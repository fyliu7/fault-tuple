
module b15s_1 ( G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, 
        G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, 
        G29, G30, G31, G32, G33, G34, G35, G36, G21356, G21357, G21358, G21359, 
        G21360, G21361, G21362, G21363, G21364, G21365, G21366, G21367, G21368, 
        G21369, G21370, G21371, G21372, G21373, G21374, G21375, G21376, G21377, 
        G21378, G21379, G21380, G21381, G21382, G21383, G21384, G21385, G21386, 
        G21387, G21388, G21389, G21390, G21391, G21392, G21393, G21394, G21395, 
        G21396, G21397, G21398, G21399, G21400, G21401, G21402, G21403, G21404, 
        G21405, G21406, G21407, G21408, G21409, G21410, G21411, G21412, G21413, 
        G21414, G21415, G21416, G21417, G21418, G21419, G21420, G21421, G21422, 
        G21423, G21424, G21425, G21426, G21427, G21428, G21429, G21430, G21431, 
        G21432, G21433, G21434, G21435, G21436, G21437, G21438, G21439, G21440, 
        G21441, G21442, G21443, G21444, G21445, G21446, G21447, G21448, G21449, 
        G21450, G21451, G21452, G21453, G21454, G21455, G21456, G21457, G21458, 
        G21459, G21460, G21461, G21462, G21463, G21464, G21465, G21466, G21467, 
        G21468, G21469, G21470, G21471, G21472, G21473, G21474, G21475, G21476, 
        G21477, G21478, G21479, G21480, G21481, G21482, G21483, G21484, G21485, 
        G21486, G21487, G21488, G21489, G21490, G21491, G21492, G21493, G21494, 
        G21495, G21496, G21497, G21498, G21499, G21500, G21501, G21502, G21503, 
        G21504, G21505, G21506, G21507, G21508, G21509, G21510, G21511, G21512, 
        G21513, G21514, G21515, G21516, G21517, G21518, G21519, G21520, G21521, 
        G21522, G21523, G21524, G21525, G21526, G21527, G21528, G21529, G21530, 
        G21531, G21532, G21533, G21534, G21535, G21536, G21537, G21538, G21539, 
        G21540, G21541, G21542, G21543, G21544, G21545, G21546, G21547, G21548, 
        G21549, G21550, G21551, G21552, G21553, G21554, G21555, G21556, G21557, 
        G21558, G21559, G21560, G21561, G21562, G21563, G21564, G21565, G21566, 
        G21567, G21568, G21569, G21570, G21571, G21572, G21573, G21574, G21575, 
        G21576, G21577, G21578, G21579, G21580, G21581, G21582, G21583, G21584, 
        G21585, G21586, G21587, G21588, G21589, G21590, G21591, G21592, G21593, 
        G21594, G21595, G21596, G21597, G21598, G21599, G21600, G21601, G21602, 
        G21603, G21604, G21605, G21606, G21607, G21608, G21609, G21610, G21611, 
        G21612, G21613, G21614, G21615, G21616, G21617, G21618, G21619, G21620, 
        G21621, G21622, G21623, G21624, G21625, G21626, G21627, G21628, G21629, 
        G21630, G21631, G21632, G21633, G21634, G21635, G21636, G21637, G21638, 
        G21639, G21640, G21641, G21642, G21643, G21644, G21645, G21646, G21647, 
        G21648, G21649, G21650, G21651, G21652, G21653, G21654, G21655, G21656, 
        G21657, G21658, G21659, G21660, G21661, G21662, G21663, G21664, G21665, 
        G21666, G21667, G21668, G21669, G21670, G21671, G21672, G21673, G21674, 
        G21675, G21676, G21677, G21678, G21679, G21680, G21681, G21682, G21683, 
        G21684, G21685, G21686, G21687, G21688, G21689, G21690, G21691, G21692, 
        G21693, G21694, G21695, G21696, G21697, G21698, G21699, G21700, G21701, 
        G21702, G21703, G21704, G21705, G21706, G21707, G21708, G21709, G21710, 
        G21711, G21712, G21713, G21714, G21715, G21716, G21717, G21718, G21719, 
        G21720, G21721, G21722, G21723, G21724, G21725, G21726, G21727, G21728, 
        G21729, G21730, G21731, G21732, G21733, G21734, G21735, G21736, G21737, 
        G21738, G21739, G21740, G21741, G21742, G21743, G21744, G21745, G21746, 
        G21747, G21748, G21749, G21750, G21751, G21752, G21753, G21754, G21755, 
        G21756, G21757, G21758, G21759, G21760, G21761, G21762, G21763, G21764, 
        G21765, G21766, G21767, G21768, G21769, G21770, G21771, G21772, G21773, 
        G21774, G21775, G21776, G21777, G21778, G21779, G21780, G21781, G21782, 
        G21783, G21784, G21785, G21786, G21787, G21788, G21789, G21790, G21791, 
        G21792, G21793, G21794, G21795, G21796, G21797, G21798, G21799, G21800, 
        G21801, G21802, G21803, G21804, G1732, G1733, G1734, G1735, G757, G758, 
        G759, G760, G761, G762, G763, G764, G765, G766, G767, G768, G769, G770, 
        G771, G772, G773, G774, G775, G776, G777, G778, G779, G780, G781, G782, 
        G783, G784, G785, G786, G787, G789, G790, G1737, G1738, G791, G792, 
        G793, G794, G795, G796, G797, G798, G799, G800, G801, G802, G803, G804, 
        G805, G806, G807, G808, G809, G810, G811, G812, G813, G814, G815, G816, 
        G817, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, 
        G829, G830, G831, G832, G833, G834, G835, G836, G837, G838, G839, G840, 
        G841, G842, G843, G844, G845, G846, G847, G848, G849, G850, G851, G852, 
        G853, G854, G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, 
        G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, 
        G877, G878, G879, G880, G881, G882, G883, G884, G885, G886, G887, G888, 
        G889, G890, G891, G892, G893, G894, G895, G896, G897, G898, G899, G900, 
        G901, G902, G903, G904, G905, G906, G907, G908, G909, G910, G911, G912, 
        G913, G914, G915, G916, G917, G918, G919, G920, G921, G922, G923, G924, 
        G925, G926, G927, G928, G929, G930, G931, G932, G933, G934, G935, G936, 
        G937, G938, G939, G940, G941, G942, G943, G944, G945, G946, G947, G948, 
        G949, G950, G951, G952, G1740, G1742, G1743, G1744, G1745, G953, G954, 
        G955, G956, G1746, G957, G958, G959, G960, G961, G962, G963, G964, 
        G965, G966, G967, G968, G969, G970, G971, G972, G973, G974, G975, G976, 
        G977, G978, G979, G980, G981, G982, G983, G984, G985, G986, G987, G988, 
        G989, G990, G991, G992, G993, G994, G995, G996, G997, G998, G999, 
        G1000, G1001, G1002, G1003, G1004, G1005, G1006, G1007, G1008, G1009, 
        G1010, G1011, G1012, G1013, G1014, G1015, G1016, G1017, G1018, G1019, 
        G1020, G1021, G1022, G1023, G1024, G1025, G1026, G1027, G1028, G1029, 
        G1030, G1031, G1032, G1033, G1034, G1035, G1036, G1037, G1038, G1039, 
        G1040, G1041, G1042, G1043, G1044, G1045, G1046, G1047, G1048, G1049, 
        G1050, G1051, G1052, G1053, G1054, G1055, G1056, G1057, G1058, G1059, 
        G1060, G1061, G1062, G1063, G1064, G1065, G1066, G1067, G1068, G1069, 
        G1070, G1071, G1072, G1073, G1074, G1075, G1076, G1077, G1078, G1079, 
        G1080, G1081, G1082, G1083, G1084, G1085, G1086, G1087, G1088, G1089, 
        G1090, G1091, G1092, G1093, G1094, G1095, G1096, G1097, G1098, G1099, 
        G1100, G1101, G1102, G1103, G1104, G1105, G1106, G1107, G1108, G1109, 
        G1110, G1111, G1112, G1113, G1114, G1115, G1116, G1117, G1118, G1119, 
        G1120, G1121, G1122, G1123, G1124, G1125, G1126, G1127, G1128, G1129, 
        G1130, G1131, G1132, G1133, G1134, G1135, G1136, G1137, G1138, G1139, 
        G1140, G1141, G1142, G1143, G1144, G1145, G1146, G1147, G1148, G1149, 
        G1150, G1151, G1152, G1153, G1154, G1155, G1156, G1157, G1158, G1159, 
        G1160, G1161, G1162, G1163, G1164, G1165, G1166, G1167, G1168, G1169, 
        G1170, G1171, G1172, G1173, G1174, G1175, G1176, G1177, G1178, G1179, 
        G1180, G1181, G1182, G1183, G1747, G1184, G1185, G1186, G1748, G1187, 
        G1749, G1188, G1189, G1750, G1751 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
         G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
         G31, G32, G33, G34, G35, G36, G21390, G21391, G21392, G21393, G21394,
         G21395, G21396, G21397, G21398, G21399, G21400, G21401, G21402,
         G21403, G21404, G21405, G21406, G21407, G21408, G21409, G21410,
         G21411, G21412, G21413, G21414, G21415, G21416, G21417, G21418,
         G21419, G21420, G21421, G21422, G21423, G21424, G21425, G21426,
         G21427, G21428, G21429, G21430, G21431, G21432, G21433, G21434,
         G21435, G21436, G21437, G21438, G21439, G21440, G21441, G21442,
         G21443, G21444, G21445, G21446, G21447, G21448, G21449, G21450,
         G21451, G21452, G21453, G21454, G21455, G21456, G21457, G21458,
         G21459, G21460, G21461, G21462, G21463, G21464, G21465, G21466,
         G21467, G21468, G21469, G21470, G21471, G21472, G21473, G21474,
         G21475, G21476, G21477, G21478, G21479, G21480, G21481, G21482,
         G21483, G21484, G21485, G21486, G21487, G21488, G21489, G21490,
         G21491, G21492, G21493, G21494, G21495, G21496, G21497, G21498,
         G21499, G21500, G21501, G21502, G21503, G21504, G21505, G21506,
         G21507, G21508, G21509, G21510, G21511, G21512, G21513, G21514,
         G21515, G21516, G21517, G21518, G21519, G21520, G21521, G21522,
         G21523, G21524, G21525, G21526, G21527, G21528, G21529, G21530,
         G21531, G21532, G21533, G21534, G21535, G21536, G21537, G21538,
         G21539, G21540, G21541, G21542, G21543, G21544, G21545, G21546,
         G21547, G21548, G21549, G21550, G21551, G21552, G21553, G21554,
         G21555, G21556, G21557, G21558, G21559, G21560, G21561, G21562,
         G21563, G21564, G21565, G21566, G21567, G21568, G21569, G21570,
         G21571, G21572, G21573, G21574, G21575, G21576, G21577, G21578,
         G21579, G21580, G21581, G21582, G21583, G21584, G21585, G21586,
         G21587, G21588, G21589, G21590, G21591, G21592, G21593, G21594,
         G21595, G21596, G21597, G21598, G21599, G21600, G21601, G21602,
         G21603, G21604, G21605, G21606, G21607, G21608, G21609, G21610,
         G21611, G21612, G21613, G21614, G21615, G21616, G21617, G21618,
         G21619, G21620, G21621, G21622, G21623, G21624, G21625, G21626,
         G21627, G21628, G21629, G21630, G21631, G21632, G21633, G21634,
         G21635, G21636, G21637, G21638, G21639, G21640, G21641, G21642,
         G21643, G21644, G21645, G21646, G21647, G21648, G21649, G21650,
         G21651, G21652, G21653, G21654, G21655, G21656, G21657, G21658,
         G21659, G21660, G21661, G21694, G21695, G21696, G21697, G21698,
         G21699, G21700, G21701, G21702, G21703, G21704, G21705, G21706,
         G21707, G21708, G21709, G21710, G21711, G21712, G21713, G21714,
         G21715, G21716, G21717, G21718, G21719, G21720, G21721, G21722,
         G21723, G21724, G21725, G21726, G21727, G21728, G21729, G21730,
         G21731, G21732, G21733, G21734, G21735, G21736, G21737, G21738,
         G21739, G21740, G21741, G21742, G21743, G21744, G21745, G21746,
         G21747, G21748, G21749, G21750, G21751, G21752, G21753, G21754,
         G21755, G21756, G21757, G21758, G21759, G21760, G21761, G21762,
         G21763, G21764, G21765, G21766, G21767, G21768, G21769, G21770,
         G21771, G21772, G21773, G21774, G21775, G21776, G21777, G21778,
         G21779, G21780, G21781, G21782, G21783, G21784, G21785, G21786,
         G21787, G21788, G21789, G21790, G21791, G21792, G21793, G21795,
         G21796, G21797, G21798, G21801, G21803, G21804,
		 
  G21356,  G21357,  G21358,  G21359,  G21360,  G21361,  G21362,  G21363, 
     G21364,  G21365,  G21366,  G21367,  G21368,  G21369,  G21370,  G21371, 
     G21372,  G21373,  G21374,  G21375,  G21376,  G21377,  G21378,  G21379, 
     G21380,  G21381,  G21382,  G21383,  G21384,  G21385,  G21386,  G21387, 
     G21388,  G21389,  G21662,  G21663,  G21664,  G21665,  G21666,  G21667, 
     G21668,  G21669,  G21670,  G21671,  G21672,  G21673,  G21674,  G21675, 
     G21676,  G21677,  G21678,  G21679,  G21680,  G21681,  G21682,  G21683, 
     G21684,  G21685,  G21686,  G21687,  G21688,  G21689,  G21690,  G21691, 
     G21692,  G21693,  G21794,  G21799,  G21800,  G21802;
	 
  output G1732, G1733, G1734, G1735, G757, G758, G759, G760, G761, G762, G763,
         G764, G765, G766, G767, G768, G769, G770, G771, G772, G773, G774,
         G775, G776, G777, G778, G779, G780, G781, G782, G783, G784, G785,
         G786, G787, G789, G790, G1737, G1738, G791, G792, G793, G794, G795,
         G796, G797, G798, G799, G800, G801, G802, G803, G804, G805, G806,
         G807, G808, G809, G810, G811, G812, G813, G814, G815, G816, G817,
         G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828,
         G829, G830, G831, G832, G833, G834, G835, G836, G837, G838, G839,
         G840, G841, G842, G843, G844, G845, G846, G847, G848, G849, G850,
         G851, G852, G853, G854, G855, G856, G857, G858, G859, G860, G861,
         G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872,
         G873, G874, G875, G876, G877, G878, G879, G880, G881, G882, G883,
         G884, G885, G886, G887, G888, G889, G890, G891, G892, G893, G894,
         G895, G896, G897, G898, G899, G900, G901, G902, G903, G904, G905,
         G906, G907, G908, G909, G910, G911, G912, G913, G914, G915, G916,
         G917, G918, G919, G920, G921, G922, G923, G924, G925, G926, G927,
         G928, G929, G930, G931, G932, G933, G934, G935, G936, G937, G938,
         G939, G940, G941, G942, G943, G944, G945, G946, G947, G948, G949,
         G950, G951, G952, G1740, G1742, G1743, G1744, G1745, G953, G954, G955,
         G956, G1746, G957, G958, G959, G960, G961, G962, G963, G964, G965,
         G966, G967, G968, G969, G970, G971, G972, G973, G974, G975, G976,
         G977, G978, G979, G980, G981, G982, G983, G984, G985, G986, G987,
         G988, G989, G990, G991, G992, G993, G994, G995, G996, G997, G998,
         G999, G1000, G1001, G1002, G1003, G1004, G1005, G1006, G1007, G1008,
         G1009, G1010, G1011, G1012, G1013, G1014, G1015, G1016, G1017, G1018,
         G1019, G1020, G1021, G1022, G1023, G1024, G1025, G1026, G1027, G1028,
         G1029, G1030, G1031, G1032, G1033, G1034, G1035, G1036, G1037, G1038,
         G1039, G1040, G1041, G1042, G1043, G1044, G1045, G1046, G1047, G1048,
         G1049, G1050, G1051, G1052, G1053, G1054, G1055, G1056, G1057, G1058,
         G1059, G1060, G1061, G1062, G1063, G1064, G1065, G1066, G1067, G1068,
         G1069, G1070, G1071, G1072, G1073, G1074, G1075, G1076, G1077, G1078,
         G1079, G1080, G1081, G1082, G1083, G1084, G1085, G1086, G1087, G1088,
         G1089, G1090, G1091, G1092, G1093, G1094, G1095, G1096, G1097, G1098,
         G1099, G1100, G1101, G1102, G1103, G1104, G1105, G1106, G1107, G1108,
         G1109, G1110, G1111, G1112, G1113, G1114, G1115, G1116, G1117, G1118,
         G1119, G1120, G1121, G1122, G1123, G1124, G1125, G1126, G1127, G1128,
         G1129, G1130, G1131, G1132, G1133, G1134, G1135, G1136, G1137, G1138,
         G1139, G1140, G1141, G1142, G1143, G1144, G1145, G1146, G1147, G1148,
         G1149, G1150, G1151, G1152, G1153, G1154, G1155, G1156, G1157, G1158,
         G1159, G1160, G1161, G1162, G1163, G1164, G1165, G1166, G1167, G1168,
         G1169, G1170, G1171, G1172, G1173, G1174, G1175, G1176, G1177, G1178,
         G1179, G1180, G1181, G1182, G1183, G1747, G1184, G1185, G1186, G1748,
         G1187, G1749, G1188, G1189, G1750, G1751;
  wire   n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592;
  nand U7357(n10305,n9290,n9110);
  nor U7358(n10047,n10042,G21428);
  not U7359(n6931,n6919);
  and U7360(n6912,n7590,n6921);
  nor U7361(n9681,n9677,n9779);
  nor U7362(n9676,n9677,n8769);
  nor U7363(n7595,n8830,n8810);
  not U7364(n9110,n7590);
  nor U7365(n7590,n9118,G21797);
  not U7366(n9936,n9953);
  nor U7367(n9953,n12764,n12765);
  nand U7368(n6921,n9293,n12973);
  nand U7369(n9346,n9651,n9652);
  nand U7370(n9344,n9649,n7456,G21428);
  and U7371(n10042,n10139,n10140);
  nand U7372(n9677,n8844,n9780);
  nor U7373(n8971,n8958,G21390);
  nor U7374(n9783,n7454,n8843);
  nor U7375(n9799,n9787,n9216);
  nor U7376(n10148,n7470,n10147);
  nor U7377(n8954,n8958,n8980);
  nor U7378(n11361,n6943,n7225);
  not U7379(n6933,n6917);
  nand U7380(n6917,n6921,n11083);
  nand U7381(n10247,n12964,n12871,n12965,n12832);
  nand U7382(n9350,n9663,n9664);
  not U7383(n7050,n7326);
  not U7384(n9101,n8737);
  nand U7385(n8737,n13571,n13572,n13573,n13574);
  and U7386(n10147,n10225,n9669);
  nand U7387(n7041,n7437,n7446);
  nand U7388(n9787,n8844,n10035);
  nand U7389(n10035,n10036,n10037,n10038,n10039);
  not U7390(n9349,n9649);
  nor U7391(n9582,n9466,n9583,n9584,n9585);
  nor U7392(n9573,n9466,n9574,n9575,n9576);
  nor U7393(n9565,n9466,n9566,n9567,n9568);
  not U7394(n9216,n10290);
  nand U7395(n11445,n11375,n10290);
  nand U7396(n11528,n11533,n10290);
  nand U7397(n11611,n11616,n10290);
  nand U7398(n11744,n11749,n10290);
  nand U7399(n12739,n12744,n10290);
  nand U7400(n12749,n12754,n10290);
  nand U7401(n12759,n12766,n10290);
  nand U7402(n10280,n10288,n10289,n10290);
  nand U7403(n10392,n10398,n10399,n10290);
  nand U7404(n12730,n12735,n12736,n10290);
  nand U7405(n10570,n10290,n10568);
  not U7406(n8958,n8972);
  not U7407(n10248,n9284);
  nor U7408(n9284,n7455,n8843);
  nand U7409(G999,n6908,n6909,n6910,n6911);
  nand U7410(n6911,n6912,n6913);
  nor U7411(n6910,n6914,n6915);
  nor U7412(n6915,n6916,n6917);
  nor U7413(n6914,n6918,n6919);
  nand U7414(n6909,n6920,G21768);
  or U7415(n6908,n6921,n6922);
  nand U7416(G998,n6923,n6924,n6925,n6926);
  nor U7417(n6926,n6927,n6928);
  nor U7418(n6928,n6929,n6921);
  and U7419(n6927,G21767,n6920);
  nand U7420(n6925,n6912,n6930);
  nand U7421(n6924,n6931,n6932);
  nand U7422(n6923,n6933,n6934);
  nand U7423(G997,n6935,n6936,n6937,n6938);
  nor U7424(n6938,n6939,n6940);
  nor U7425(n6940,n6941,n6921);
  nor U7426(n6939,n6942,n6943);
  nand U7427(n6937,n6912,n6944);
  nand U7428(n6936,n6931,n6945);
  nand U7429(n6935,n6933,n6946);
  nand U7430(G996,n6947,n6948,n6949,n6950);
  nor U7431(n6950,n6951,n6952);
  nor U7432(n6952,n6953,n6921);
  nor U7433(n6951,n6954,n6943);
  nand U7434(n6949,n6912,n6955);
  nand U7435(n6948,n6956,n6931);
  nand U7436(n6947,n6933,n6957);
  nand U7437(G995,n6958,n6959,n6960,n6961);
  nor U7438(n6961,n6962,n6963);
  nor U7439(n6963,n6964,n6921);
  nor U7440(n6962,n6965,n6943);
  nand U7441(n6960,n6912,n6966);
  nand U7442(n6959,n6967,n6931);
  nand U7443(n6958,n6933,n6968);
  nand U7444(G994,n6969,n6970,n6971,n6972);
  nor U7445(n6972,n6973,n6974);
  nor U7446(n6974,n6975,n6921);
  nor U7447(n6973,n6976,n6943);
  nand U7448(n6971,n6912,n6977);
  nand U7449(n6970,n6978,n6931);
  nand U7450(n6969,n6933,n6979);
  nand U7451(G993,n6980,n6981,n6982,n6983);
  nor U7452(n6983,n6984,n6985);
  nor U7453(n6985,n6986,n6921);
  nor U7454(n6984,n6987,n6943);
  nand U7455(n6982,n6912,n6988);
  nand U7456(n6981,n6989,n6931);
  nand U7457(n6980,n6933,n6990);
  nand U7458(G992,n6991,n6992,n6993,n6994);
  nor U7459(n6994,n6995,n6996);
  nor U7460(n6996,n6997,n6921);
  nor U7461(n6995,n6998,n6943);
  nand U7462(n6993,n6912,n6999);
  nand U7463(n6992,n7000,n6931);
  nand U7464(n6991,n6933,n7001);
  nand U7465(G991,n7002,n7003,n7004,n7005);
  nor U7466(n7005,n7006,n7007);
  nor U7467(n7007,n7008,n6921);
  and U7468(n7006,G21760,n6920);
  nand U7469(n7004,n6912,n7009);
  nand U7470(n7003,n7010,n6931);
  nand U7471(n7002,n6933,n7011);
  nand U7472(G990,n7012,n7013,n7014,n7015);
  nor U7473(n7015,n7016,n7017);
  nor U7474(n7017,n7018,n6921);
  nor U7475(n7016,n7019,n6943);
  nand U7476(n7014,n6912,n7020);
  nand U7477(n7013,n7021,n6931);
  nand U7478(n7012,n6933,n7022);
  nand U7479(G989,n7023,n7024,n7025,n7026);
  nor U7480(n7026,n7027,n7028);
  nor U7481(n7028,n7029,n6921);
  nor U7482(n7027,n7030,n6943);
  nand U7483(n7025,n6912,n7031);
  nand U7484(n7024,n6931,n7032);
  nand U7485(n7023,n6933,n7033);
  nand U7486(G988,n7034,n7035,n7036,n7037);
  nor U7487(n7037,n7038,n7039,n7040);
  nor U7488(n7040,G21598,n7041,n7042);
  nor U7489(n7039,n7043,n7044);
  nor U7490(n7043,n7045,n7046);
  and U7491(n7045,n7042,n7047);
  nor U7492(n7038,n7048,n7049);
  nand U7493(n7036,n7050,n7051);
  nand U7494(n7035,n7052,n7053);
  nand U7495(n7034,n7054,n7055);
  nand U7496(G987,n7056,n7057,n7058,n7059);
  nor U7497(n7059,n7060,n7061,n7062);
  nor U7498(n7062,n7063,n7064);
  and U7499(n7061,n7047,n7042,n7065);
  nor U7500(n7060,n7066,n7067);
  nand U7501(n7058,n7046,G21597);
  nand U7502(n7057,n7050,n7068);
  nand U7503(n7056,n7069,G21788);
  nand U7504(G986,n7070,n7071,n7072,n7073);
  nor U7505(n7073,n7074,n7075,n7076);
  nor U7506(n7076,n7063,n7077);
  nor U7507(n7075,n7041,n7078,n7079);
  nor U7508(n7074,n7080,n7067);
  nand U7509(n7072,n7046,G21596);
  nand U7510(n7071,n7050,n7081);
  nand U7511(n7070,n7069,G21787);
  nand U7512(G985,n7082,n7083,n7084,n7085);
  nor U7513(n7085,n7086,n7087,n7088);
  nor U7514(n7088,n7063,n7089);
  and U7515(n7087,n7047,n7090,n7091);
  nor U7516(n7086,n7092,n7067);
  nand U7517(n7084,n7046,G21595);
  nand U7518(n7083,n7050,n7093);
  nand U7519(n7082,n7069,G21786);
  nand U7520(G984,n7094,n7095,n7096,n7097);
  nor U7521(n7097,n7098,n7099,n7100);
  nor U7522(n7100,n7063,n7101);
  nor U7523(n7099,n7041,n7102,n7103);
  nor U7524(n7098,n7104,n7067);
  nand U7525(n7096,n7046,G21594);
  nand U7526(n7095,n7050,n7105);
  nand U7527(n7094,n7069,G21785);
  nand U7528(G983,n7106,n7107,n7108,n7109);
  nor U7529(n7109,n7110,n7111,n7112);
  nor U7530(n7112,n7063,n7113);
  nor U7531(n7111,n7041,n7114,n7115);
  nor U7532(n7110,n7116,n7067);
  nand U7533(n7108,n7046,G21593);
  nand U7534(n7107,n7050,n7117);
  nand U7535(n7106,n7069,G21784);
  nand U7536(G982,n7118,n7119,n7120,n7121);
  nor U7537(n7121,n7122,n7123,n7124);
  nor U7538(n7124,n7125,n7049);
  nor U7539(n7123,n7126,n7041);
  nor U7540(n7122,n7127,n7128);
  nand U7541(n7120,n7050,n7129);
  nand U7542(n7119,n7130,n7052);
  nand U7543(n7118,n7054,n7131);
  nand U7544(G981,n7132,n7133,n7134,n7135);
  nor U7545(n7135,n7136,n7137,n7138);
  nor U7546(n7138,n7063,n7139);
  nor U7547(n7137,n7140,n7041);
  nor U7548(n7136,n7141,n7067);
  nand U7549(n7134,n7046,G21591);
  nand U7550(n7133,n7050,n7142);
  nand U7551(n7132,n7069,G21782);
  nand U7552(G980,n7143,n7144,n7145,n7146);
  nor U7553(n7146,n7147,n7148,n7149);
  nor U7554(n7149,n7150,n7049);
  nor U7555(n7148,n7151,n7041);
  and U7556(n7147,G21590,n7046);
  nand U7557(n7145,n7050,n7152);
  nand U7558(n7144,n7153,n7052);
  nand U7559(n7143,n7054,n7154);
  nand U7560(G979,n7155,n7156,n7157,n7158);
  nor U7561(n7158,n7159,n7160,n7161);
  nor U7562(n7161,n7162,n7049);
  nor U7563(n7160,n7163,n7041);
  nor U7564(n7159,n7164,n7128);
  nand U7565(n7157,n7050,n7165);
  nand U7566(n7156,n7166,n7052);
  nand U7567(n7155,n7054,n7167);
  nand U7568(G978,n7168,n7169,n7170,n7171);
  nor U7569(n7171,n7172,n7173,n7174);
  nor U7570(n7174,n7175,n7049);
  nor U7571(n7173,n7176,n7041);
  nor U7572(n7172,n7177,n7128);
  nand U7573(n7170,n7050,n7178);
  nand U7574(n7169,n7179,n7052);
  nand U7575(n7168,n7054,n7180);
  nand U7576(G977,n7181,n7182,n7183,n7184);
  nor U7577(n7184,n7185,n7186,n7187);
  nor U7578(n7187,n7188,n7049);
  nor U7579(n7186,n7189,n7041);
  and U7580(n7185,G21587,n7046);
  nand U7581(n7183,n7050,n7190);
  nand U7582(n7182,n7191,n7052);
  nand U7583(n7181,n7054,n7192);
  nand U7584(G976,n7193,n7194,n7195,n7196);
  nor U7585(n7196,n7197,n7198,n7199);
  nor U7586(n7199,n7200,n7049);
  nor U7587(n7198,n7201,n7041);
  nor U7588(n7197,n7202,n7128);
  nand U7589(n7195,n7050,n7203);
  nand U7590(n7194,n7204,n7052);
  nand U7591(n7193,n7054,n7205);
  nand U7592(G975,n7206,n7207,n7208,n7209);
  nor U7593(n7209,n7210,n7211,n7212);
  nor U7594(n7212,n7213,n7049);
  nor U7595(n7211,n7214,n7041);
  and U7596(n7210,G21585,n7046);
  nand U7597(n7208,n7050,n7215);
  nand U7598(n7207,n7216,n7052);
  nand U7599(n7206,n7054,n7217);
  nand U7600(G974,n7218,n7219,n7220,n7221);
  nor U7601(n7221,n7222,n7223,n7224);
  nor U7602(n7224,n7225,n7049);
  nor U7603(n7223,n7226,n7041);
  nor U7604(n7222,n7227,n7128);
  nand U7605(n7220,n7050,n7228);
  nand U7606(n7219,n7229,n7052);
  nand U7607(n7218,n7054,n7230);
  nand U7608(G973,n7231,n7232,n7233,n7234);
  nor U7609(n7234,n7235,n7236,n7237);
  nor U7610(n7237,n7238,n7049);
  nor U7611(n7236,n7239,n7041);
  nor U7612(n7235,n7240,n7128);
  nand U7613(n7233,n7050,n7241);
  nand U7614(n7232,n7052,n7242);
  nand U7615(n7231,n7054,n7243);
  nand U7616(G972,n7244,n7245,n7246,n7247);
  nor U7617(n7247,n7248,n7249,n7250);
  nor U7618(n7250,G21582,n7041,n7251,n7252);
  nor U7619(n7249,n7253,n7254);
  nor U7620(n7253,n7255,n7256);
  nor U7621(n7255,G21581,n7041);
  nor U7622(n7248,n7257,n7049);
  nand U7623(n7246,n7050,n7258);
  nand U7624(n7245,n7259,n7052);
  nand U7625(n7244,n7054,n7260);
  nand U7626(G971,n7261,n7262,n7263,n7264);
  nor U7627(n7264,n7265,n7266,n7267);
  nor U7628(n7267,G21581,n7252,n7041);
  and U7629(n7266,n7256,G21581);
  nand U7630(n7256,n7128,n7268);
  nand U7631(n7268,n7047,n7252);
  nor U7632(n7265,n7269,n7049);
  nand U7633(n7263,n7050,n7270);
  nand U7634(n7262,n7271,n7052);
  nand U7635(n7261,n7054,n7272);
  nand U7636(G970,n7273,n7274,n7275,n7276);
  nor U7637(n7276,n7277,n7278,n7279);
  nor U7638(n7279,G21580,n7041,n7280,n7281);
  nor U7639(n7278,n7282,n7283);
  nor U7640(n7282,n7284,n7285);
  nor U7641(n7284,G21579,n7041);
  nor U7642(n7277,n7286,n7049);
  nand U7643(n7275,n7050,n7287);
  nand U7644(n7274,n7288,n7052);
  nand U7645(n7273,n7054,n7289);
  nand U7646(G969,n7290,n7291,n7292,n7293);
  nor U7647(n7293,n7294,n7295,n7296);
  nor U7648(n7296,G21579,n7281,n7041);
  and U7649(n7295,n7285,G21579);
  nand U7650(n7285,n7128,n7297);
  nand U7651(n7297,n7047,n7281);
  nor U7652(n7294,n7298,n7049);
  nand U7653(n7292,n7050,n7299);
  nand U7654(n7291,n7300,n7052);
  nand U7655(n7290,n7054,n7301);
  nand U7656(G968,n7302,n7303,n7304,n7305);
  nor U7657(n7305,n7306,n7307,n7308);
  nor U7658(n7308,G21578,n7041,n7309,n7310);
  nor U7659(n7307,n7311,n7312);
  not U7660(n7312,G21578);
  nor U7661(n7311,n7313,n7314);
  nor U7662(n7313,G21577,n7041);
  and U7663(n7306,G21769,n7069);
  nand U7664(n7304,n7315,n7050);
  nand U7665(n7303,n7316,n7052);
  nand U7666(n7302,n7054,n7317);
  nand U7667(G967,n7318,n7319,n7320,n7321);
  nor U7668(n7321,n7322,n7323,n7324);
  nor U7669(n7324,n7325,n7067);
  nor U7670(n7323,n6916,n7063);
  nor U7671(n7322,n6918,n7326);
  nand U7672(n7320,n7069,G21768);
  nand U7673(n7319,G21577,n7314);
  nand U7674(n7314,n7128,n7327);
  nand U7675(n7327,n7047,n7310);
  not U7676(n7310,n7328);
  nand U7677(n7318,n7047,n7328,n7309);
  not U7678(n7309,G21577);
  nand U7679(G966,n7329,n7330,n7331,n7332);
  nor U7680(n7332,n7333,n7334,n7335);
  nor U7681(n7335,n7336,n7063);
  nor U7682(n7334,n7337,n7041);
  or U7683(n7337,n7338,n7339);
  nor U7684(n7333,n7340,n7067);
  nand U7685(n7331,n7046,G21576);
  nand U7686(n7330,n7050,n6932);
  nand U7687(n7329,n7069,G21767);
  nand U7688(G965,n7341,n7342,n7343,n7344);
  nor U7689(n7344,n7345,n7346,n7347);
  and U7690(n7347,n7348,n7349,n7047);
  nor U7691(n7346,n7350,n7348);
  not U7692(n7348,G21575);
  nor U7693(n7350,n7351,n7046);
  nor U7694(n7351,n7349,n7041);
  nor U7695(n7345,n6942,n7049);
  not U7696(n6942,G21766);
  nand U7697(n7343,n7050,n6945);
  nand U7698(n7342,n7052,n6946);
  nand U7699(n7341,n7054,n6944);
  nand U7700(G964,n7352,n7353,n7354,n7355);
  nor U7701(n7355,n7356,n7357,n7358);
  nor U7702(n7358,G21574,n7041,n7359,n7360);
  nor U7703(n7357,n7361,n7362);
  nor U7704(n7361,n7363,n7364);
  nor U7705(n7363,G21573,n7041);
  nor U7706(n7356,n6954,n7049);
  not U7707(n6954,G21765);
  nand U7708(n7354,n7050,n6956);
  nand U7709(n7353,n7052,n6957);
  nand U7710(n7352,n7054,n6955);
  nand U7711(G963,n7365,n7366,n7367,n7368);
  nor U7712(n7368,n7369,n7370,n7371);
  nor U7713(n7371,G21573,n7360,n7041);
  and U7714(n7370,n7364,G21573);
  nand U7715(n7364,n7128,n7372);
  nand U7716(n7372,n7047,n7360);
  nor U7717(n7369,n6965,n7049);
  not U7718(n6965,G21764);
  nand U7719(n7367,n7050,n6967);
  nand U7720(n7366,n7052,n6968);
  nand U7721(n7365,n7054,n6966);
  nand U7722(G962,n7373,n7374,n7375,n7376);
  nor U7723(n7376,n7377,n7378,n7379);
  nor U7724(n7379,G21572,n7041,n7380,n7381);
  nor U7725(n7378,n7382,n7383);
  not U7726(n7383,G21572);
  nor U7727(n7382,n7384,n7385);
  nor U7728(n7384,G21571,n7041);
  nor U7729(n7377,n6976,n7049);
  not U7730(n6976,G21763);
  nand U7731(n7375,n7050,n6978);
  nand U7732(n7374,n7052,n6979);
  nand U7733(n7373,n7054,n6977);
  nand U7734(G961,n7386,n7387,n7388,n7389);
  nor U7735(n7389,n7390,n7391,n7392);
  nor U7736(n7392,G21571,n7381,n7041);
  nor U7737(n7391,n7393,n7380);
  not U7738(n7380,G21571);
  nor U7739(n7390,n6987,n7049);
  nand U7740(n7388,n7050,n6989);
  nand U7741(n7387,n7052,n6990);
  nand U7742(n7386,n7054,n6988);
  nand U7743(G960,n7394,n7395,n7396,n7397);
  nor U7744(n7397,n7398,n7399,n7400);
  nor U7745(n7400,n7393,n7401);
  not U7746(n7393,n7385);
  nand U7747(n7385,n7128,n7402);
  nand U7748(n7402,n7047,n7381);
  not U7749(n7381,n7403);
  nor U7750(n7399,n7041,n7403,n7404);
  nor U7751(n7398,n7405,n7063);
  nand U7752(n7396,n7069,G21761);
  nand U7753(n7395,n7054,n6999);
  nand U7754(n7394,n7050,n7000);
  nand U7755(G959,n7406,n7407,n7408,n7409);
  nor U7756(n7409,n7410,n7411,n7412);
  nor U7757(n7412,n7413,n7063);
  nor U7758(n7411,n7414,n7041);
  nor U7759(n7414,n7415,n7404);
  nor U7760(n7415,n7416,n7417);
  nor U7761(n7410,n7418,n7067);
  nand U7762(n7408,n7046,G21569);
  nand U7763(n7407,n7050,n7010);
  nand U7764(n7406,n7069,G21760);
  nand U7765(G958,n7419,n7420,n7421,n7422);
  nor U7766(n7422,n7423,n7424,n7425);
  and U7767(n7425,n7426,n7427,n7047);
  not U7768(n7047,n7041);
  nor U7769(n7424,n7428,n7426);
  nor U7770(n7428,n7429,n7046);
  nor U7771(n7423,n7019,n7049);
  not U7772(n7049,n7069);
  nand U7773(n7421,n7050,n7021);
  nand U7774(n7420,n7052,n7022);
  not U7775(n7052,n7063);
  nand U7776(n7419,n7054,n7020);
  not U7777(n7054,n7067);
  nand U7778(G957,n7430,n7431,n7432,n7433);
  nor U7779(n7433,n7434,n7429,n7435);
  nor U7780(n7435,n7436,n7063);
  nand U7781(n7063,n7437,n7438);
  nand U7782(n7438,n7439,n7440,n7441,n7442);
  not U7783(n7442,n7443);
  nor U7784(n7441,n7444,n7445);
  nor U7785(n7429,n7427,n7041);
  nor U7786(n7434,n7447,n7067);
  nand U7787(n7067,n7437,n7448);
  nand U7788(n7448,n7449,n7450);
  nand U7789(n7432,n7046,G21567);
  nand U7790(n7431,n7050,n7032);
  nand U7791(n7326,n7437,n7451);
  nand U7792(n7451,n7452,n7453,n7454,n7455);
  nor U7793(n7437,n7456,n7046);
  nand U7794(n7430,n7069,G21758);
  nor U7795(n7069,n7046,G21426);
  not U7796(n7046,n7128);
  nand U7797(n7128,n7457,n7458);
  nand U7798(n7458,n7459,n7460);
  nand U7799(n7460,n7461,n7462,n7463,n7464);
  nand U7800(n7464,n7465,n7466,n7467);
  nand U7801(n7466,n7468,n7469);
  nand U7802(n7469,n7470,n7471,n7472);
  nand U7803(n7463,n7473,n7474);
  nand U7804(n7474,n7475,n7476);
  nand U7805(n7476,n7477,n7478);
  nand U7806(n7478,n7465,n7479);
  nand U7807(n7479,n7480,n7481);
  nand U7808(n7475,n7480,n7482);
  nand U7809(n7462,n7483,n7484);
  nand U7810(G956,n7485,n7486,n7487);
  nand U7811(n7487,n7488,G21565);
  nand U7812(n7486,n7489,n7490);
  nand U7813(n7485,n7491,n7020);
  nand U7814(G955,n7492,n7493,n7494);
  nand U7815(n7494,n7488,G21564);
  nand U7816(n7493,n7495,n7489);
  nand U7817(n7492,n7491,n7009);
  nand U7818(G954,n7496,n7497,n7498);
  nand U7819(n7498,n7488,G21563);
  nand U7820(n7497,n7499,n7489);
  nand U7821(n7496,n7491,n6999);
  nor U7822(G953,n7500,n7501);
  nand U7823(G952,n7502,n7503,n7504,n7505);
  nor U7824(n7505,n7506,n7507,n7508);
  nor U7825(n7508,n7509,n7510);
  nor U7826(n7507,n7511,n7512);
  nor U7827(n7506,n7513,n7514);
  nand U7828(n7504,G32,n7515);
  nand U7829(n7503,G21556,n7516);
  nand U7830(n7502,G16,n7517);
  nand U7831(G951,n7518,n7519,n7520,n7521);
  nor U7832(n7521,n7522,n7523,n7524);
  nor U7833(n7524,n7525,n7510);
  nor U7834(n7523,n7511,n7526);
  nor U7835(n7522,n7513,n7527);
  nand U7836(n7520,G31,n7515);
  nand U7837(n7519,G21555,n7516);
  nand U7838(n7518,G15,n7517);
  nand U7839(G950,n7528,n7529,n7530,n7531);
  nor U7840(n7531,n7532,n7533,n7534);
  nor U7841(n7534,n7535,n7510);
  nor U7842(n7533,n7511,n7536);
  nor U7843(n7532,n7513,n7537);
  nand U7844(n7530,G30,n7515);
  nand U7845(n7529,G21554,n7516);
  nand U7846(n7528,G14,n7517);
  nand U7847(G949,n7538,n7539,n7540,n7541);
  nor U7848(n7541,n7542,n7543,n7544);
  nor U7849(n7544,n7545,n7510);
  nor U7850(n7543,n7511,n7546);
  nor U7851(n7542,n7513,n7547);
  nand U7852(n7540,G29,n7515);
  nand U7853(n7539,G21553,n7516);
  nand U7854(n7538,G13,n7517);
  nand U7855(G948,n7548,n7549,n7550,n7551);
  nor U7856(n7551,n7552,n7553,n7554);
  nor U7857(n7554,n7555,n7510);
  nor U7858(n7553,n7511,n7556);
  nor U7859(n7552,n7513,n7557);
  nand U7860(n7550,G28,n7515);
  nand U7861(n7549,G21552,n7516);
  nand U7862(n7548,G12,n7517);
  nand U7863(G947,n7558,n7559,n7560,n7561);
  nor U7864(n7561,n7562,n7563,n7564);
  nor U7865(n7564,n7565,n7510);
  nor U7866(n7563,n7511,n7566);
  nor U7867(n7562,n7513,n7567);
  nand U7868(n7560,G27,n7515);
  nand U7869(n7559,G21551,n7516);
  nand U7870(n7558,G11,n7517);
  nand U7871(G946,n7568,n7569,n7570,n7571);
  nor U7872(n7571,n7572,n7573,n7574);
  nor U7873(n7574,n7575,n7510);
  nor U7874(n7573,n7511,n7576);
  nor U7875(n7572,n7513,n7577);
  nand U7876(n7570,G26,n7515);
  nand U7877(n7569,G21550,n7516);
  nand U7878(n7568,G10,n7517);
  nand U7879(G945,n7578,n7579,n7580,n7581);
  nor U7880(n7581,n7582,n7583,n7584);
  nor U7881(n7584,n7585,n7510);
  nor U7882(n7583,n7511,n7586);
  and U7883(n7511,n7587,n7588);
  nand U7884(n7588,n7589,n7590);
  nand U7885(n7587,n7591,G21426);
  nor U7886(n7582,n7513,n7592);
  nand U7887(n7580,G25,n7515);
  nand U7888(n7515,n7593,n7594);
  nand U7889(n7594,n7589,n7595,n7513,n7596);
  not U7890(n7589,n7597);
  nand U7891(n7593,n7598,n7599);
  nand U7892(n7579,G21549,n7516);
  nand U7893(n7516,n7600,n7601);
  nand U7894(n7601,n7602,n7603,n7604);
  nand U7895(n7604,n7605,n7591);
  nand U7896(n7602,n7599,n7606);
  not U7897(n7599,n7510);
  nand U7898(n7600,n7598,n7510);
  nand U7899(n7510,n7607,n7608);
  and U7900(n7598,n7609,n7597);
  nand U7901(n7597,n7610,n7611);
  nand U7902(n7609,n7612,n7613);
  nand U7903(n7613,n7513,n7596,n7595);
  nand U7904(n7578,G9,n7517);
  and U7905(n7517,n7591,n7513,n7595);
  not U7906(n7591,n7596);
  nand U7907(G944,n7614,n7615,n7616,n7617);
  nor U7908(n7617,n7618,n7619,n7620);
  nor U7909(n7620,n7509,n7621);
  nor U7910(n7619,n7622,n7512);
  nor U7911(n7618,n7623,n7514);
  nand U7912(n7616,G32,n7624);
  nand U7913(n7615,G21548,n7625);
  nand U7914(n7614,n7626,G16);
  nand U7915(G943,n7627,n7628,n7629,n7630);
  nor U7916(n7630,n7631,n7632,n7633);
  nor U7917(n7633,n7525,n7621);
  nor U7918(n7632,n7622,n7526);
  nor U7919(n7631,n7623,n7527);
  nand U7920(n7629,G31,n7624);
  nand U7921(n7628,G21547,n7625);
  nand U7922(n7627,n7626,G15);
  nand U7923(G942,n7634,n7635,n7636,n7637);
  nor U7924(n7637,n7638,n7639,n7640);
  nor U7925(n7640,n7535,n7621);
  nor U7926(n7639,n7622,n7536);
  nor U7927(n7638,n7623,n7537);
  nand U7928(n7636,G30,n7624);
  nand U7929(n7635,G21546,n7625);
  nand U7930(n7634,n7626,G14);
  nand U7931(G941,n7641,n7642,n7643,n7644);
  nor U7932(n7644,n7645,n7646,n7647);
  nor U7933(n7647,n7545,n7621);
  nor U7934(n7646,n7622,n7546);
  nor U7935(n7645,n7623,n7547);
  nand U7936(n7643,G29,n7624);
  nand U7937(n7642,G21545,n7625);
  nand U7938(n7641,n7626,G13);
  nand U7939(G940,n7648,n7649,n7650,n7651);
  nor U7940(n7651,n7652,n7653,n7654);
  nor U7941(n7654,n7555,n7621);
  nor U7942(n7653,n7622,n7556);
  nor U7943(n7652,n7623,n7557);
  nand U7944(n7650,G28,n7624);
  nand U7945(n7649,G21544,n7625);
  nand U7946(n7648,n7626,G12);
  nand U7947(G939,n7655,n7656,n7657,n7658);
  nor U7948(n7658,n7659,n7660,n7661);
  nor U7949(n7661,n7565,n7621);
  nor U7950(n7660,n7622,n7566);
  nor U7951(n7659,n7623,n7567);
  nand U7952(n7657,G27,n7624);
  nand U7953(n7656,G21543,n7625);
  nand U7954(n7655,n7626,G11);
  nand U7955(G938,n7662,n7663,n7664,n7665);
  nor U7956(n7665,n7666,n7667,n7668);
  nor U7957(n7668,n7575,n7621);
  nor U7958(n7667,n7622,n7576);
  nor U7959(n7666,n7623,n7577);
  nand U7960(n7664,G26,n7624);
  nand U7961(n7663,G21542,n7625);
  nand U7962(n7662,n7626,G10);
  nand U7963(G937,n7669,n7670,n7671,n7672);
  nor U7964(n7672,n7673,n7674,n7675);
  nor U7965(n7675,n7585,n7621);
  nor U7966(n7674,n7622,n7586);
  and U7967(n7622,n7676,n7677);
  nand U7968(n7677,n7678,n7590);
  nand U7969(n7676,n7679,G21426);
  nor U7970(n7673,n7623,n7592);
  nand U7971(n7671,G25,n7624);
  nand U7972(n7624,n7680,n7681);
  nand U7973(n7681,n7678,n7595,n7623,n7682);
  not U7974(n7678,n7683);
  nand U7975(n7680,n7684,n7685);
  nand U7976(n7670,G21541,n7625);
  nand U7977(n7625,n7686,n7687);
  nand U7978(n7687,n7688,n7603,n7689);
  nand U7979(n7689,n7605,n7679);
  nand U7980(n7688,n7685,n7606);
  not U7981(n7685,n7621);
  nand U7982(n7686,n7684,n7621);
  nand U7983(n7621,n7690,n7608);
  and U7984(n7684,n7691,n7683);
  nand U7985(n7683,n7692,n7611);
  nand U7986(n7691,n7612,n7693);
  nand U7987(n7693,n7623,n7682,n7595);
  nand U7988(n7669,n7626,G9);
  and U7989(n7626,n7679,n7623,n7595);
  not U7990(n7679,n7682);
  nand U7991(G936,n7694,n7695,n7696,n7697);
  nor U7992(n7697,n7698,n7699,n7700);
  nor U7993(n7700,n7509,n7701);
  nor U7994(n7699,n7702,n7512);
  nor U7995(n7698,n7703,n7514);
  nand U7996(n7696,G32,n7704);
  nand U7997(n7695,G21540,n7705);
  nand U7998(n7694,n7706,G16);
  nand U7999(G935,n7707,n7708,n7709,n7710);
  nor U8000(n7710,n7711,n7712,n7713);
  nor U8001(n7713,n7525,n7701);
  nor U8002(n7712,n7702,n7526);
  nor U8003(n7711,n7703,n7527);
  nand U8004(n7709,G31,n7704);
  nand U8005(n7708,G21539,n7705);
  nand U8006(n7707,n7706,G15);
  nand U8007(G934,n7714,n7715,n7716,n7717);
  nor U8008(n7717,n7718,n7719,n7720);
  nor U8009(n7720,n7535,n7701);
  nor U8010(n7719,n7702,n7536);
  nor U8011(n7718,n7703,n7537);
  nand U8012(n7716,G30,n7704);
  nand U8013(n7715,G21538,n7705);
  nand U8014(n7714,n7706,G14);
  nand U8015(G933,n7721,n7722,n7723,n7724);
  nor U8016(n7724,n7725,n7726,n7727);
  nor U8017(n7727,n7545,n7701);
  nor U8018(n7726,n7702,n7546);
  nor U8019(n7725,n7703,n7547);
  nand U8020(n7723,G29,n7704);
  nand U8021(n7722,G21537,n7705);
  nand U8022(n7721,n7706,G13);
  nand U8023(G932,n7728,n7729,n7730,n7731);
  nor U8024(n7731,n7732,n7733,n7734);
  nor U8025(n7734,n7555,n7701);
  nor U8026(n7733,n7702,n7556);
  nor U8027(n7732,n7703,n7557);
  nand U8028(n7730,G28,n7704);
  nand U8029(n7729,G21536,n7705);
  nand U8030(n7728,n7706,G12);
  nand U8031(G931,n7735,n7736,n7737,n7738);
  nor U8032(n7738,n7739,n7740,n7741);
  nor U8033(n7741,n7565,n7701);
  nor U8034(n7740,n7702,n7566);
  nor U8035(n7739,n7703,n7567);
  nand U8036(n7737,G27,n7704);
  nand U8037(n7736,G21535,n7705);
  nand U8038(n7735,n7706,G11);
  nand U8039(G930,n7742,n7743,n7744,n7745);
  nor U8040(n7745,n7746,n7747,n7748);
  nor U8041(n7748,n7575,n7701);
  nor U8042(n7747,n7702,n7576);
  nor U8043(n7746,n7703,n7577);
  nand U8044(n7744,G26,n7704);
  nand U8045(n7743,G21534,n7705);
  nand U8046(n7742,n7706,G10);
  nand U8047(G929,n7749,n7750,n7751,n7752);
  nor U8048(n7752,n7753,n7754,n7755);
  nor U8049(n7755,n7585,n7701);
  nor U8050(n7754,n7702,n7586);
  and U8051(n7702,n7756,n7757);
  nand U8052(n7757,n7758,n7590);
  nand U8053(n7756,n7759,G21426);
  nor U8054(n7753,n7703,n7592);
  nand U8055(n7751,G25,n7704);
  nand U8056(n7704,n7760,n7761);
  nand U8057(n7761,n7758,n7595,n7703,n7762);
  not U8058(n7758,n7763);
  nand U8059(n7760,n7764,n7765);
  nand U8060(n7750,G21533,n7705);
  nand U8061(n7705,n7766,n7767);
  nand U8062(n7767,n7768,n7603,n7769);
  nand U8063(n7769,n7605,n7759);
  nand U8064(n7768,n7765,n7606);
  not U8065(n7765,n7701);
  nand U8066(n7766,n7764,n7701);
  nand U8067(n7701,n7770,n7608);
  and U8068(n7764,n7771,n7763);
  nand U8069(n7763,n7772,n7611);
  nand U8070(n7771,n7612,n7773);
  nand U8071(n7773,n7703,n7762,n7595);
  nand U8072(n7749,n7706,G9);
  and U8073(n7706,n7759,n7703,n7595);
  not U8074(n7759,n7762);
  nand U8075(G928,n7774,n7775,n7776,n7777);
  nor U8076(n7777,n7778,n7779,n7780);
  nor U8077(n7780,n7509,n7781);
  nor U8078(n7779,n7782,n7512);
  nor U8079(n7778,n7783,n7514);
  nand U8080(n7776,G32,n7784);
  nand U8081(n7775,G21532,n7785);
  nand U8082(n7774,n7786,G16);
  nand U8083(G927,n7787,n7788,n7789,n7790);
  nor U8084(n7790,n7791,n7792,n7793);
  nor U8085(n7793,n7525,n7781);
  nor U8086(n7792,n7782,n7526);
  nor U8087(n7791,n7783,n7527);
  nand U8088(n7789,G31,n7784);
  nand U8089(n7788,G21531,n7785);
  nand U8090(n7787,n7786,G15);
  nand U8091(G926,n7794,n7795,n7796,n7797);
  nor U8092(n7797,n7798,n7799,n7800);
  nor U8093(n7800,n7535,n7781);
  nor U8094(n7799,n7782,n7536);
  nor U8095(n7798,n7783,n7537);
  nand U8096(n7796,G30,n7784);
  nand U8097(n7795,G21530,n7785);
  nand U8098(n7794,n7786,G14);
  nand U8099(G925,n7801,n7802,n7803,n7804);
  nor U8100(n7804,n7805,n7806,n7807);
  nor U8101(n7807,n7545,n7781);
  nor U8102(n7806,n7782,n7546);
  nor U8103(n7805,n7783,n7547);
  nand U8104(n7803,G29,n7784);
  nand U8105(n7802,G21529,n7785);
  nand U8106(n7801,n7786,G13);
  nand U8107(G924,n7808,n7809,n7810,n7811);
  nor U8108(n7811,n7812,n7813,n7814);
  nor U8109(n7814,n7555,n7781);
  nor U8110(n7813,n7782,n7556);
  nor U8111(n7812,n7783,n7557);
  nand U8112(n7810,G28,n7784);
  nand U8113(n7809,G21528,n7785);
  nand U8114(n7808,n7786,G12);
  nand U8115(G923,n7815,n7816,n7817,n7818);
  nor U8116(n7818,n7819,n7820,n7821);
  nor U8117(n7821,n7565,n7781);
  nor U8118(n7820,n7782,n7566);
  nor U8119(n7819,n7783,n7567);
  nand U8120(n7817,G27,n7784);
  nand U8121(n7816,G21527,n7785);
  nand U8122(n7815,n7786,G11);
  nand U8123(G922,n7822,n7823,n7824,n7825);
  nor U8124(n7825,n7826,n7827,n7828);
  nor U8125(n7828,n7575,n7781);
  nor U8126(n7827,n7782,n7576);
  nor U8127(n7826,n7783,n7577);
  nand U8128(n7824,G26,n7784);
  nand U8129(n7823,G21526,n7785);
  nand U8130(n7822,n7786,G10);
  nand U8131(G921,n7829,n7830,n7831,n7832);
  nor U8132(n7832,n7833,n7834,n7835);
  nor U8133(n7835,n7585,n7781);
  nor U8134(n7834,n7782,n7586);
  and U8135(n7782,n7836,n7837);
  nand U8136(n7837,n7838,n7590);
  nand U8137(n7836,n7839,G21426);
  nor U8138(n7833,n7783,n7592);
  nand U8139(n7831,G25,n7784);
  nand U8140(n7784,n7840,n7841);
  nand U8141(n7841,n7838,n7595,n7783,n7842);
  not U8142(n7838,n7843);
  nand U8143(n7840,n7844,n7845);
  nand U8144(n7830,G21525,n7785);
  nand U8145(n7785,n7846,n7847);
  nand U8146(n7847,n7848,n7603,n7849);
  nand U8147(n7849,n7605,n7839);
  nand U8148(n7848,n7845,n7606);
  not U8149(n7845,n7781);
  nand U8150(n7846,n7844,n7781);
  nand U8151(n7781,n7608,n7850);
  nor U8152(n7608,G21564,G21563);
  and U8153(n7844,n7851,n7843);
  nand U8154(n7843,n7852,n7611);
  nor U8155(n7611,n7853,n7854);
  nand U8156(n7851,n7612,n7855);
  nand U8157(n7855,n7783,n7842,n7595);
  nand U8158(n7829,n7786,G9);
  and U8159(n7786,n7839,n7783,n7595);
  not U8160(n7839,n7842);
  nand U8161(G920,n7856,n7857,n7858,n7859);
  nor U8162(n7859,n7860,n7861,n7862);
  nor U8163(n7862,n7509,n7863);
  nor U8164(n7861,n7864,n7512);
  nor U8165(n7860,n7865,n7514);
  nand U8166(n7858,G32,n7866);
  nand U8167(n7857,G21524,n7867);
  nand U8168(n7856,n7868,G16);
  nand U8169(G919,n7869,n7870,n7871,n7872);
  nor U8170(n7872,n7873,n7874,n7875);
  nor U8171(n7875,n7525,n7863);
  nor U8172(n7874,n7864,n7526);
  nor U8173(n7873,n7865,n7527);
  nand U8174(n7871,G31,n7866);
  nand U8175(n7870,G21523,n7867);
  nand U8176(n7869,n7868,G15);
  nand U8177(G918,n7876,n7877,n7878,n7879);
  nor U8178(n7879,n7880,n7881,n7882);
  nor U8179(n7882,n7535,n7863);
  nor U8180(n7881,n7864,n7536);
  nor U8181(n7880,n7865,n7537);
  nand U8182(n7878,G30,n7866);
  nand U8183(n7877,G21522,n7867);
  nand U8184(n7876,n7868,G14);
  nand U8185(G917,n7883,n7884,n7885,n7886);
  nor U8186(n7886,n7887,n7888,n7889);
  nor U8187(n7889,n7545,n7863);
  nor U8188(n7888,n7864,n7546);
  nor U8189(n7887,n7865,n7547);
  nand U8190(n7885,G29,n7866);
  nand U8191(n7884,G21521,n7867);
  nand U8192(n7883,n7868,G13);
  nand U8193(G916,n7890,n7891,n7892,n7893);
  nor U8194(n7893,n7894,n7895,n7896);
  nor U8195(n7896,n7555,n7863);
  nor U8196(n7895,n7864,n7556);
  nor U8197(n7894,n7865,n7557);
  nand U8198(n7892,G28,n7866);
  nand U8199(n7891,G21520,n7867);
  nand U8200(n7890,n7868,G12);
  nand U8201(G915,n7897,n7898,n7899,n7900);
  nor U8202(n7900,n7901,n7902,n7903);
  nor U8203(n7903,n7565,n7863);
  nor U8204(n7902,n7864,n7566);
  nor U8205(n7901,n7865,n7567);
  nand U8206(n7899,G27,n7866);
  nand U8207(n7898,G21519,n7867);
  nand U8208(n7897,n7868,G11);
  nand U8209(G914,n7904,n7905,n7906,n7907);
  nor U8210(n7907,n7908,n7909,n7910);
  nor U8211(n7910,n7575,n7863);
  nor U8212(n7909,n7864,n7576);
  nor U8213(n7908,n7865,n7577);
  nand U8214(n7906,G26,n7866);
  nand U8215(n7905,G21518,n7867);
  nand U8216(n7904,n7868,G10);
  nand U8217(G913,n7911,n7912,n7913,n7914);
  nor U8218(n7914,n7915,n7916,n7917);
  nor U8219(n7917,n7585,n7863);
  nor U8220(n7916,n7864,n7586);
  and U8221(n7864,n7918,n7919);
  nand U8222(n7919,n7920,n7590);
  nand U8223(n7918,n7921,G21426);
  nor U8224(n7915,n7865,n7592);
  nand U8225(n7913,G25,n7866);
  nand U8226(n7866,n7922,n7923);
  nand U8227(n7923,n7920,n7595,n7865,n7924);
  not U8228(n7920,n7925);
  nand U8229(n7922,n7926,n7927);
  nand U8230(n7912,G21517,n7867);
  nand U8231(n7867,n7928,n7929);
  nand U8232(n7929,n7930,n7603,n7931);
  nand U8233(n7931,n7605,n7921);
  nand U8234(n7930,n7927,n7606);
  not U8235(n7927,n7863);
  nand U8236(n7928,n7926,n7863);
  nand U8237(n7863,n7607,n7932);
  and U8238(n7926,n7933,n7925);
  nand U8239(n7925,n7934,n7610);
  nand U8240(n7933,n7612,n7935);
  nand U8241(n7935,n7865,n7924,n7595);
  nand U8242(n7911,n7868,G9);
  and U8243(n7868,n7921,n7865,n7595);
  not U8244(n7921,n7924);
  nand U8245(G912,n7936,n7937,n7938,n7939);
  nor U8246(n7939,n7940,n7941,n7942);
  nor U8247(n7942,n7509,n7943);
  nor U8248(n7941,n7944,n7512);
  nor U8249(n7940,n7945,n7514);
  nand U8250(n7938,G32,n7946);
  nand U8251(n7937,G21516,n7947);
  nand U8252(n7936,n7948,G16);
  nand U8253(G911,n7949,n7950,n7951,n7952);
  nor U8254(n7952,n7953,n7954,n7955);
  nor U8255(n7955,n7525,n7943);
  nor U8256(n7954,n7944,n7526);
  nor U8257(n7953,n7945,n7527);
  nand U8258(n7951,G31,n7946);
  nand U8259(n7950,G21515,n7947);
  nand U8260(n7949,n7948,G15);
  nand U8261(G910,n7956,n7957,n7958,n7959);
  nor U8262(n7959,n7960,n7961,n7962);
  nor U8263(n7962,n7535,n7943);
  nor U8264(n7961,n7944,n7536);
  nor U8265(n7960,n7945,n7537);
  nand U8266(n7958,G30,n7946);
  nand U8267(n7957,G21514,n7947);
  nand U8268(n7956,n7948,G14);
  nand U8269(G909,n7963,n7964,n7965,n7966);
  nor U8270(n7966,n7967,n7968,n7969);
  nor U8271(n7969,n7545,n7943);
  nor U8272(n7968,n7944,n7546);
  nor U8273(n7967,n7945,n7547);
  nand U8274(n7965,G29,n7946);
  nand U8275(n7964,G21513,n7947);
  nand U8276(n7963,n7948,G13);
  nand U8277(G908,n7970,n7971,n7972,n7973);
  nor U8278(n7973,n7974,n7975,n7976);
  nor U8279(n7976,n7555,n7943);
  nor U8280(n7975,n7944,n7556);
  nor U8281(n7974,n7945,n7557);
  nand U8282(n7972,G28,n7946);
  nand U8283(n7971,G21512,n7947);
  nand U8284(n7970,n7948,G12);
  nand U8285(G907,n7977,n7978,n7979,n7980);
  nor U8286(n7980,n7981,n7982,n7983);
  nor U8287(n7983,n7565,n7943);
  nor U8288(n7982,n7944,n7566);
  nor U8289(n7981,n7945,n7567);
  nand U8290(n7979,G27,n7946);
  nand U8291(n7978,G21511,n7947);
  nand U8292(n7977,n7948,G11);
  nand U8293(G906,n7984,n7985,n7986,n7987);
  nor U8294(n7987,n7988,n7989,n7990);
  nor U8295(n7990,n7575,n7943);
  nor U8296(n7989,n7944,n7576);
  nor U8297(n7988,n7945,n7577);
  nand U8298(n7986,G26,n7946);
  nand U8299(n7985,G21510,n7947);
  nand U8300(n7984,n7948,G10);
  nand U8301(G905,n7991,n7992,n7993,n7994);
  nor U8302(n7994,n7995,n7996,n7997);
  nor U8303(n7997,n7585,n7943);
  nor U8304(n7996,n7944,n7586);
  and U8305(n7944,n7998,n7999);
  nand U8306(n7999,n8000,n7590);
  nand U8307(n7998,n8001,G21426);
  nor U8308(n7995,n7945,n7592);
  nand U8309(n7993,G25,n7946);
  nand U8310(n7946,n8002,n8003);
  nand U8311(n8003,n8000,n7595,n7945,n8004);
  not U8312(n8000,n8005);
  nand U8313(n8002,n8006,n8007);
  nand U8314(n7992,G21509,n7947);
  nand U8315(n7947,n8008,n8009);
  nand U8316(n8009,n8010,n7603,n8011);
  nand U8317(n8011,n7605,n8001);
  nand U8318(n8010,n8007,n7606);
  not U8319(n8007,n7943);
  nand U8320(n8008,n8006,n7943);
  nand U8321(n7943,n7690,n7932);
  and U8322(n8006,n8012,n8005);
  nand U8323(n8005,n7934,n7692);
  nand U8324(n8012,n7612,n8013);
  nand U8325(n8013,n7945,n8004,n7595);
  nand U8326(n7991,n7948,G9);
  and U8327(n7948,n8001,n7945,n7595);
  not U8328(n8001,n8004);
  nand U8329(G904,n8014,n8015,n8016,n8017);
  nor U8330(n8017,n8018,n8019,n8020);
  nor U8331(n8020,n7509,n8021);
  nor U8332(n8019,n8022,n7512);
  nor U8333(n8018,n8023,n7514);
  nand U8334(n8016,G32,n8024);
  nand U8335(n8015,G21508,n8025);
  nand U8336(n8014,n8026,G16);
  nand U8337(G903,n8027,n8028,n8029,n8030);
  nor U8338(n8030,n8031,n8032,n8033);
  nor U8339(n8033,n7525,n8021);
  nor U8340(n8032,n8022,n7526);
  nor U8341(n8031,n8023,n7527);
  nand U8342(n8029,G31,n8024);
  nand U8343(n8028,G21507,n8025);
  nand U8344(n8027,n8026,G15);
  nand U8345(G902,n8034,n8035,n8036,n8037);
  nor U8346(n8037,n8038,n8039,n8040);
  nor U8347(n8040,n7535,n8021);
  nor U8348(n8039,n8022,n7536);
  nor U8349(n8038,n8023,n7537);
  nand U8350(n8036,G30,n8024);
  nand U8351(n8035,G21506,n8025);
  nand U8352(n8034,n8026,G14);
  nand U8353(G901,n8041,n8042,n8043,n8044);
  nor U8354(n8044,n8045,n8046,n8047);
  nor U8355(n8047,n7545,n8021);
  nor U8356(n8046,n8022,n7546);
  nor U8357(n8045,n8023,n7547);
  nand U8358(n8043,G29,n8024);
  nand U8359(n8042,G21505,n8025);
  nand U8360(n8041,n8026,G13);
  nand U8361(G900,n8048,n8049,n8050,n8051);
  nor U8362(n8051,n8052,n8053,n8054);
  nor U8363(n8054,n7555,n8021);
  nor U8364(n8053,n8022,n7556);
  nor U8365(n8052,n8023,n7557);
  nand U8366(n8050,G28,n8024);
  nand U8367(n8049,G21504,n8025);
  nand U8368(n8048,n8026,G12);
  nand U8369(G899,n8055,n8056,n8057,n8058);
  nor U8370(n8058,n8059,n8060,n8061);
  nor U8371(n8061,n7565,n8021);
  nor U8372(n8060,n8022,n7566);
  nor U8373(n8059,n8023,n7567);
  nand U8374(n8057,G27,n8024);
  nand U8375(n8056,G21503,n8025);
  nand U8376(n8055,n8026,G11);
  nand U8377(G898,n8062,n8063,n8064,n8065);
  nor U8378(n8065,n8066,n8067,n8068);
  nor U8379(n8068,n7575,n8021);
  nor U8380(n8067,n8022,n7576);
  nor U8381(n8066,n8023,n7577);
  nand U8382(n8064,G26,n8024);
  nand U8383(n8063,G21502,n8025);
  nand U8384(n8062,n8026,G10);
  nand U8385(G897,n8069,n8070,n8071,n8072);
  nor U8386(n8072,n8073,n8074,n8075);
  nor U8387(n8075,n7585,n8021);
  nor U8388(n8074,n8022,n7586);
  and U8389(n8022,n8076,n8077);
  nand U8390(n8077,n8078,n7590);
  nand U8391(n8076,n8079,G21426);
  nor U8392(n8073,n8023,n7592);
  nand U8393(n8071,G25,n8024);
  nand U8394(n8024,n8080,n8081);
  nand U8395(n8081,n8078,n7595,n8023,n8082);
  not U8396(n8078,n8083);
  nand U8397(n8080,n8084,n8085);
  nand U8398(n8070,G21501,n8025);
  nand U8399(n8025,n8086,n8087);
  nand U8400(n8087,n8088,n7603,n8089);
  nand U8401(n8089,n7605,n8079);
  nand U8402(n8088,n8085,n7606);
  not U8403(n8085,n8021);
  nand U8404(n8086,n8084,n8021);
  nand U8405(n8021,n7770,n7932);
  and U8406(n8084,n8090,n8083);
  nand U8407(n8083,n7934,n7772);
  nand U8408(n8090,n7612,n8091);
  nand U8409(n8091,n8023,n8082,n7595);
  nand U8410(n8069,n8026,G9);
  and U8411(n8026,n8079,n8023,n7595);
  not U8412(n8079,n8082);
  nand U8413(G896,n8092,n8093,n8094,n8095);
  nor U8414(n8095,n8096,n8097,n8098);
  nor U8415(n8098,n7509,n8099);
  nor U8416(n8097,n8100,n7512);
  nor U8417(n8096,n8101,n7514);
  nand U8418(n8094,G32,n8102);
  nand U8419(n8093,G21500,n8103);
  nand U8420(n8092,n8104,G16);
  nand U8421(G895,n8105,n8106,n8107,n8108);
  nor U8422(n8108,n8109,n8110,n8111);
  nor U8423(n8111,n7525,n8099);
  nor U8424(n8110,n8100,n7526);
  nor U8425(n8109,n8101,n7527);
  nand U8426(n8107,G31,n8102);
  nand U8427(n8106,G21499,n8103);
  nand U8428(n8105,n8104,G15);
  nand U8429(G894,n8112,n8113,n8114,n8115);
  nor U8430(n8115,n8116,n8117,n8118);
  nor U8431(n8118,n7535,n8099);
  nor U8432(n8117,n8100,n7536);
  nor U8433(n8116,n8101,n7537);
  nand U8434(n8114,G30,n8102);
  nand U8435(n8113,G21498,n8103);
  nand U8436(n8112,n8104,G14);
  nand U8437(G893,n8119,n8120,n8121,n8122);
  nor U8438(n8122,n8123,n8124,n8125);
  nor U8439(n8125,n7545,n8099);
  nor U8440(n8124,n8100,n7546);
  nor U8441(n8123,n8101,n7547);
  nand U8442(n8121,G29,n8102);
  nand U8443(n8120,G21497,n8103);
  nand U8444(n8119,n8104,G13);
  nand U8445(G892,n8126,n8127,n8128,n8129);
  nor U8446(n8129,n8130,n8131,n8132);
  nor U8447(n8132,n7555,n8099);
  nor U8448(n8131,n8100,n7556);
  nor U8449(n8130,n8101,n7557);
  nand U8450(n8128,G28,n8102);
  nand U8451(n8127,G21496,n8103);
  nand U8452(n8126,n8104,G12);
  nand U8453(G891,n8133,n8134,n8135,n8136);
  nor U8454(n8136,n8137,n8138,n8139);
  nor U8455(n8139,n7565,n8099);
  nor U8456(n8138,n8100,n7566);
  nor U8457(n8137,n8101,n7567);
  nand U8458(n8135,G27,n8102);
  nand U8459(n8134,G21495,n8103);
  nand U8460(n8133,n8104,G11);
  nand U8461(G890,n8140,n8141,n8142,n8143);
  nor U8462(n8143,n8144,n8145,n8146);
  nor U8463(n8146,n7575,n8099);
  nor U8464(n8145,n8100,n7576);
  nor U8465(n8144,n8101,n7577);
  nand U8466(n8142,G26,n8102);
  nand U8467(n8141,G21494,n8103);
  nand U8468(n8140,n8104,G10);
  nand U8469(G889,n8147,n8148,n8149,n8150);
  nor U8470(n8150,n8151,n8152,n8153);
  nor U8471(n8153,n7585,n8099);
  nor U8472(n8152,n8100,n7586);
  and U8473(n8100,n8154,n8155);
  nand U8474(n8155,n8156,n7590);
  nand U8475(n8154,n8157,G21426);
  nor U8476(n8151,n8101,n7592);
  nand U8477(n8149,G25,n8102);
  nand U8478(n8102,n8158,n8159);
  nand U8479(n8159,n8156,n7595,n8101,n8160);
  not U8480(n8156,n8161);
  nand U8481(n8158,n8162,n8163);
  nand U8482(n8148,G21493,n8103);
  nand U8483(n8103,n8164,n8165);
  nand U8484(n8165,n8166,n7603,n8167);
  nand U8485(n8167,n8163,n7606);
  nand U8486(n8166,n7605,n8157);
  nand U8487(n8164,n8162,n8099);
  and U8488(n8162,n8168,n8161);
  nand U8489(n8161,n7934,n7852);
  nor U8490(n7934,n7853,n8169);
  not U8491(n7853,n8170);
  nand U8492(n8168,n7612,n8171);
  nand U8493(n8171,n8101,n8160,n7595);
  nand U8494(n8147,n8104,G9);
  and U8495(n8104,n8157,n8101,n7595);
  not U8496(n8157,n8160);
  nand U8497(G888,n8172,n8173,n8174,n8175);
  nor U8498(n8175,n8176,n8177,n8178);
  nor U8499(n8178,n7509,n8179);
  nor U8500(n8177,n8180,n7512);
  nor U8501(n8176,n8181,n7514);
  nand U8502(n8174,G32,n8182);
  nand U8503(n8173,G21492,n8183);
  nand U8504(n8172,n8184,G16);
  nand U8505(G887,n8185,n8186,n8187,n8188);
  nor U8506(n8188,n8189,n8190,n8191);
  nor U8507(n8191,n7525,n8179);
  nor U8508(n8190,n8180,n7526);
  nor U8509(n8189,n8181,n7527);
  nand U8510(n8187,G31,n8182);
  nand U8511(n8186,G21491,n8183);
  nand U8512(n8185,n8184,G15);
  nand U8513(G886,n8192,n8193,n8194,n8195);
  nor U8514(n8195,n8196,n8197,n8198);
  nor U8515(n8198,n7535,n8179);
  nor U8516(n8197,n8180,n7536);
  nor U8517(n8196,n8181,n7537);
  nand U8518(n8194,G30,n8182);
  nand U8519(n8193,G21490,n8183);
  nand U8520(n8192,n8184,G14);
  nand U8521(G885,n8199,n8200,n8201,n8202);
  nor U8522(n8202,n8203,n8204,n8205);
  nor U8523(n8205,n7545,n8179);
  nor U8524(n8204,n8180,n7546);
  nor U8525(n8203,n8181,n7547);
  nand U8526(n8201,G29,n8182);
  nand U8527(n8200,G21489,n8183);
  nand U8528(n8199,n8184,G13);
  nand U8529(G884,n8206,n8207,n8208,n8209);
  nor U8530(n8209,n8210,n8211,n8212);
  nor U8531(n8212,n7555,n8179);
  nor U8532(n8211,n8180,n7556);
  nor U8533(n8210,n8181,n7557);
  nand U8534(n8208,G28,n8182);
  nand U8535(n8207,G21488,n8183);
  nand U8536(n8206,n8184,G12);
  nand U8537(G883,n8213,n8214,n8215,n8216);
  nor U8538(n8216,n8217,n8218,n8219);
  nor U8539(n8219,n7565,n8179);
  nor U8540(n8218,n8180,n7566);
  nor U8541(n8217,n8181,n7567);
  nand U8542(n8215,G27,n8182);
  nand U8543(n8214,G21487,n8183);
  nand U8544(n8213,n8184,G11);
  nand U8545(G882,n8220,n8221,n8222,n8223);
  nor U8546(n8223,n8224,n8225,n8226);
  nor U8547(n8226,n7575,n8179);
  nor U8548(n8225,n8180,n7576);
  nor U8549(n8224,n8181,n7577);
  nand U8550(n8222,G26,n8182);
  nand U8551(n8221,G21486,n8183);
  nand U8552(n8220,n8184,G10);
  nand U8553(G881,n8227,n8228,n8229,n8230);
  nor U8554(n8230,n8231,n8232,n8233);
  nor U8555(n8233,n7585,n8179);
  nor U8556(n8232,n8180,n7586);
  and U8557(n8180,n8234,n8235);
  nand U8558(n8235,n8236,n7590);
  nand U8559(n8234,n8237,G21426);
  nor U8560(n8231,n8181,n7592);
  nand U8561(n8229,G25,n8182);
  nand U8562(n8182,n8238,n8239);
  nand U8563(n8239,n8236,n7595,n8181,n8240);
  not U8564(n8236,n8241);
  nand U8565(n8238,n8242,n8243);
  nand U8566(n8228,G21485,n8183);
  nand U8567(n8183,n8244,n8245);
  nand U8568(n8245,n8246,n7603,n8247);
  nand U8569(n8247,n7605,n8237);
  nand U8570(n8246,n8243,n7606);
  not U8571(n8243,n8179);
  nand U8572(n8244,n8242,n8179);
  nand U8573(n8179,n8248,n7607);
  and U8574(n8242,n8249,n8241);
  nand U8575(n8241,n8250,n7610);
  nand U8576(n8249,n7612,n8251);
  nand U8577(n8251,n8181,n8240,n7595);
  nand U8578(n8227,n8184,G9);
  and U8579(n8184,n8237,n8181,n7595);
  not U8580(n8237,n8240);
  nand U8581(G880,n8252,n8253,n8254,n8255);
  nor U8582(n8255,n8256,n8257,n8258);
  nor U8583(n8258,n7509,n8259);
  nor U8584(n8257,n8260,n7512);
  nor U8585(n8256,n8261,n7514);
  nand U8586(n8254,G32,n8262);
  nand U8587(n8253,G21484,n8263);
  nand U8588(n8252,n8264,G16);
  nand U8589(G879,n8265,n8266,n8267,n8268);
  nor U8590(n8268,n8269,n8270,n8271);
  nor U8591(n8271,n7525,n8259);
  nor U8592(n8270,n8260,n7526);
  nor U8593(n8269,n8261,n7527);
  nand U8594(n8267,G31,n8262);
  nand U8595(n8266,G21483,n8263);
  nand U8596(n8265,n8264,G15);
  nand U8597(G878,n8272,n8273,n8274,n8275);
  nor U8598(n8275,n8276,n8277,n8278);
  nor U8599(n8278,n7535,n8259);
  nor U8600(n8277,n8260,n7536);
  nor U8601(n8276,n8261,n7537);
  nand U8602(n8274,G30,n8262);
  nand U8603(n8273,G21482,n8263);
  nand U8604(n8272,n8264,G14);
  nand U8605(G877,n8279,n8280,n8281,n8282);
  nor U8606(n8282,n8283,n8284,n8285);
  nor U8607(n8285,n7545,n8259);
  nor U8608(n8284,n8260,n7546);
  nor U8609(n8283,n8261,n7547);
  nand U8610(n8281,G29,n8262);
  nand U8611(n8280,G21481,n8263);
  nand U8612(n8279,n8264,G13);
  nand U8613(G876,n8286,n8287,n8288,n8289);
  nor U8614(n8289,n8290,n8291,n8292);
  nor U8615(n8292,n7555,n8259);
  nor U8616(n8291,n8260,n7556);
  nor U8617(n8290,n8261,n7557);
  nand U8618(n8288,G28,n8262);
  nand U8619(n8287,G21480,n8263);
  nand U8620(n8286,n8264,G12);
  nand U8621(G875,n8293,n8294,n8295,n8296);
  nor U8622(n8296,n8297,n8298,n8299);
  nor U8623(n8299,n7565,n8259);
  nor U8624(n8298,n8260,n7566);
  nor U8625(n8297,n8261,n7567);
  nand U8626(n8295,G27,n8262);
  nand U8627(n8294,G21479,n8263);
  nand U8628(n8293,n8264,G11);
  nand U8629(G874,n8300,n8301,n8302,n8303);
  nor U8630(n8303,n8304,n8305,n8306);
  nor U8631(n8306,n7575,n8259);
  nor U8632(n8305,n8260,n7576);
  nor U8633(n8304,n8261,n7577);
  nand U8634(n8302,G26,n8262);
  nand U8635(n8301,G21478,n8263);
  nand U8636(n8300,n8264,G10);
  nand U8637(G873,n8307,n8308,n8309,n8310);
  nor U8638(n8310,n8311,n8312,n8313);
  nor U8639(n8313,n7585,n8259);
  nor U8640(n8312,n8260,n7586);
  and U8641(n8260,n8314,n8315);
  nand U8642(n8315,n8316,n7590);
  nand U8643(n8314,n8317,G21426);
  nor U8644(n8311,n8261,n7592);
  nand U8645(n8309,G25,n8262);
  nand U8646(n8262,n8318,n8319);
  nand U8647(n8319,n8316,n7595,n8261,n8320);
  not U8648(n8316,n8321);
  nand U8649(n8318,n8322,n8323);
  nand U8650(n8308,G21477,n8263);
  nand U8651(n8263,n8324,n8325);
  nand U8652(n8325,n8326,n7603,n8327);
  nand U8653(n8327,n7605,n8317);
  nand U8654(n8326,n8323,n7606);
  not U8655(n8323,n8259);
  nand U8656(n8324,n8322,n8259);
  nand U8657(n8259,n8248,n7690);
  and U8658(n8322,n8328,n8321);
  nand U8659(n8321,n8250,n7692);
  nand U8660(n8328,n7612,n8329);
  nand U8661(n8329,n8261,n8320,n7595);
  nand U8662(n8307,n8264,G9);
  and U8663(n8264,n8317,n8261,n7595);
  not U8664(n8317,n8320);
  nand U8665(G872,n8330,n8331,n8332,n8333);
  nor U8666(n8333,n8334,n8335,n8336);
  nor U8667(n8336,n7509,n8337);
  nor U8668(n8335,n8338,n7512);
  nor U8669(n8334,n8339,n7514);
  nand U8670(n8332,G32,n8340);
  nand U8671(n8331,G21476,n8341);
  nand U8672(n8330,n8342,G16);
  nand U8673(G871,n8343,n8344,n8345,n8346);
  nor U8674(n8346,n8347,n8348,n8349);
  nor U8675(n8349,n7525,n8337);
  nor U8676(n8348,n8338,n7526);
  nor U8677(n8347,n8339,n7527);
  nand U8678(n8345,G31,n8340);
  nand U8679(n8344,G21475,n8341);
  nand U8680(n8343,n8342,G15);
  nand U8681(G870,n8350,n8351,n8352,n8353);
  nor U8682(n8353,n8354,n8355,n8356);
  nor U8683(n8356,n7535,n8337);
  nor U8684(n8355,n8338,n7536);
  nor U8685(n8354,n8339,n7537);
  nand U8686(n8352,G30,n8340);
  nand U8687(n8351,G21474,n8341);
  nand U8688(n8350,n8342,G14);
  nand U8689(G869,n8357,n8358,n8359,n8360);
  nor U8690(n8360,n8361,n8362,n8363);
  nor U8691(n8363,n7545,n8337);
  nor U8692(n8362,n8338,n7546);
  nor U8693(n8361,n8339,n7547);
  nand U8694(n8359,G29,n8340);
  nand U8695(n8358,G21473,n8341);
  nand U8696(n8357,n8342,G13);
  nand U8697(G868,n8364,n8365,n8366,n8367);
  nor U8698(n8367,n8368,n8369,n8370);
  nor U8699(n8370,n7555,n8337);
  nor U8700(n8369,n8338,n7556);
  nor U8701(n8368,n8339,n7557);
  nand U8702(n8366,G28,n8340);
  nand U8703(n8365,G21472,n8341);
  nand U8704(n8364,n8342,G12);
  nand U8705(G867,n8371,n8372,n8373,n8374);
  nor U8706(n8374,n8375,n8376,n8377);
  nor U8707(n8377,n7565,n8337);
  nor U8708(n8376,n8338,n7566);
  nor U8709(n8375,n8339,n7567);
  nand U8710(n8373,G27,n8340);
  nand U8711(n8372,G21471,n8341);
  nand U8712(n8371,n8342,G11);
  nand U8713(G866,n8378,n8379,n8380,n8381);
  nor U8714(n8381,n8382,n8383,n8384);
  nor U8715(n8384,n7575,n8337);
  nor U8716(n8383,n8338,n7576);
  nor U8717(n8382,n8339,n7577);
  nand U8718(n8380,G26,n8340);
  nand U8719(n8379,G21470,n8341);
  nand U8720(n8378,n8342,G10);
  nand U8721(G865,n8385,n8386,n8387,n8388);
  nor U8722(n8388,n8389,n8390,n8391);
  nor U8723(n8391,n7585,n8337);
  nor U8724(n8390,n8338,n7586);
  and U8725(n8338,n8392,n8393);
  nand U8726(n8393,n8394,n7590);
  nand U8727(n8392,n8395,G21426);
  nor U8728(n8389,n8339,n7592);
  nand U8729(n8387,G25,n8340);
  nand U8730(n8340,n8396,n8397);
  nand U8731(n8397,n8394,n7595,n8339,n8398);
  not U8732(n8394,n8399);
  nand U8733(n8396,n8400,n8401);
  nand U8734(n8386,G21469,n8341);
  nand U8735(n8341,n8402,n8403);
  nand U8736(n8403,n8404,n7603,n8405);
  nand U8737(n8405,n7605,n8395);
  nand U8738(n8404,n8401,n7606);
  not U8739(n8401,n8337);
  nand U8740(n8402,n8400,n8337);
  nand U8741(n8337,n8248,n7770);
  and U8742(n8400,n8406,n8399);
  nand U8743(n8399,n8250,n7772);
  nand U8744(n8406,n7612,n8407);
  nand U8745(n8407,n8339,n8398,n7595);
  nand U8746(n8385,n8342,G9);
  and U8747(n8342,n8395,n8339,n7595);
  not U8748(n8395,n8398);
  nand U8749(G864,n8408,n8409,n8410,n8411);
  nor U8750(n8411,n8412,n8413,n8414);
  nor U8751(n8414,n7509,n8415);
  nor U8752(n8413,n8416,n7512);
  nor U8753(n8412,n8417,n7514);
  nand U8754(n8410,G32,n8418);
  nand U8755(n8409,G21468,n8419);
  nand U8756(n8408,n8420,G16);
  nand U8757(G863,n8421,n8422,n8423,n8424);
  nor U8758(n8424,n8425,n8426,n8427);
  nor U8759(n8427,n7525,n8415);
  nor U8760(n8426,n8416,n7526);
  nor U8761(n8425,n8417,n7527);
  nand U8762(n8423,G31,n8418);
  nand U8763(n8422,G21467,n8419);
  nand U8764(n8421,n8420,G15);
  nand U8765(G862,n8428,n8429,n8430,n8431);
  nor U8766(n8431,n8432,n8433,n8434);
  nor U8767(n8434,n7535,n8415);
  nor U8768(n8433,n8416,n7536);
  nor U8769(n8432,n8417,n7537);
  nand U8770(n8430,G30,n8418);
  nand U8771(n8429,G21466,n8419);
  nand U8772(n8428,n8420,G14);
  nand U8773(G861,n8435,n8436,n8437,n8438);
  nor U8774(n8438,n8439,n8440,n8441);
  nor U8775(n8441,n7545,n8415);
  nor U8776(n8440,n8416,n7546);
  nor U8777(n8439,n8417,n7547);
  nand U8778(n8437,G29,n8418);
  nand U8779(n8436,G21465,n8419);
  nand U8780(n8435,n8420,G13);
  nand U8781(G860,n8442,n8443,n8444,n8445);
  nor U8782(n8445,n8446,n8447,n8448);
  nor U8783(n8448,n7555,n8415);
  nor U8784(n8447,n8416,n7556);
  nor U8785(n8446,n8417,n7557);
  nand U8786(n8444,G28,n8418);
  nand U8787(n8443,G21464,n8419);
  nand U8788(n8442,n8420,G12);
  nand U8789(G859,n8449,n8450,n8451,n8452);
  nor U8790(n8452,n8453,n8454,n8455);
  nor U8791(n8455,n7565,n8415);
  nor U8792(n8454,n8416,n7566);
  nor U8793(n8453,n8417,n7567);
  nand U8794(n8451,G27,n8418);
  nand U8795(n8450,G21463,n8419);
  nand U8796(n8449,n8420,G11);
  nand U8797(G858,n8456,n8457,n8458,n8459);
  nor U8798(n8459,n8460,n8461,n8462);
  nor U8799(n8462,n7575,n8415);
  nor U8800(n8461,n8416,n7576);
  nor U8801(n8460,n8417,n7577);
  nand U8802(n8458,G26,n8418);
  nand U8803(n8457,G21462,n8419);
  nand U8804(n8456,n8420,G10);
  nand U8805(G857,n8463,n8464,n8465,n8466);
  nor U8806(n8466,n8467,n8468,n8469);
  nor U8807(n8469,n7585,n8415);
  nor U8808(n8468,n8416,n7586);
  and U8809(n8416,n8470,n8471);
  nand U8810(n8471,n8472,n7590);
  nand U8811(n8470,n8473,G21426);
  nor U8812(n8467,n8417,n7592);
  nand U8813(n8465,G25,n8418);
  nand U8814(n8418,n8474,n8475);
  nand U8815(n8475,n8472,n7595,n8417,n8476);
  not U8816(n8472,n8477);
  nand U8817(n8474,n8478,n8479);
  nand U8818(n8464,G21461,n8419);
  nand U8819(n8419,n8480,n8481);
  nand U8820(n8481,n8482,n7603,n8483);
  nand U8821(n8483,n7605,n8473);
  nand U8822(n8482,n8479,n7606);
  not U8823(n8479,n8415);
  nand U8824(n8480,n8478,n8415);
  nand U8825(n8415,n8248,n7850);
  and U8826(n8478,n8484,n8477);
  nand U8827(n8477,n8250,n7852);
  nor U8828(n8250,n7854,n8170);
  nand U8829(n8484,n7612,n8485);
  nand U8830(n8485,n8417,n8476,n7595);
  nand U8831(n8463,n8420,G9);
  and U8832(n8420,n8473,n8417,n7595);
  not U8833(n8473,n8476);
  nand U8834(G856,n8486,n8487,n8488,n8489);
  nor U8835(n8489,n8490,n8491,n8492);
  nor U8836(n8492,n7509,n8493);
  nor U8837(n8491,n8494,n7512);
  nor U8838(n8490,n8495,n7514);
  nand U8839(n8488,G32,n8496);
  nand U8840(n8487,G21460,n8497);
  nand U8841(n8486,n8498,G16);
  nand U8842(G855,n8499,n8500,n8501,n8502);
  nor U8843(n8502,n8503,n8504,n8505);
  nor U8844(n8505,n7525,n8493);
  nor U8845(n8504,n8494,n7526);
  nor U8846(n8503,n8495,n7527);
  nand U8847(n8501,G31,n8496);
  nand U8848(n8500,G21459,n8497);
  nand U8849(n8499,n8498,G15);
  nand U8850(G854,n8506,n8507,n8508,n8509);
  nor U8851(n8509,n8510,n8511,n8512);
  nor U8852(n8512,n7535,n8493);
  nor U8853(n8511,n8494,n7536);
  nor U8854(n8510,n8495,n7537);
  nand U8855(n8508,G30,n8496);
  nand U8856(n8507,G21458,n8497);
  nand U8857(n8506,n8498,G14);
  nand U8858(G853,n8513,n8514,n8515,n8516);
  nor U8859(n8516,n8517,n8518,n8519);
  nor U8860(n8519,n7545,n8493);
  nor U8861(n8518,n8494,n7546);
  nor U8862(n8517,n8495,n7547);
  nand U8863(n8515,G29,n8496);
  nand U8864(n8514,G21457,n8497);
  nand U8865(n8513,n8498,G13);
  nand U8866(G852,n8520,n8521,n8522,n8523);
  nor U8867(n8523,n8524,n8525,n8526);
  nor U8868(n8526,n7555,n8493);
  nor U8869(n8525,n8494,n7556);
  nor U8870(n8524,n8495,n7557);
  nand U8871(n8522,G28,n8496);
  nand U8872(n8521,G21456,n8497);
  nand U8873(n8520,n8498,G12);
  nand U8874(G851,n8527,n8528,n8529,n8530);
  nor U8875(n8530,n8531,n8532,n8533);
  nor U8876(n8533,n7565,n8493);
  nor U8877(n8532,n8494,n7566);
  nor U8878(n8531,n8495,n7567);
  nand U8879(n8529,G27,n8496);
  nand U8880(n8528,G21455,n8497);
  nand U8881(n8527,n8498,G11);
  nand U8882(G850,n8534,n8535,n8536,n8537);
  nor U8883(n8537,n8538,n8539,n8540);
  nor U8884(n8540,n7575,n8493);
  nor U8885(n8539,n8494,n7576);
  nor U8886(n8538,n8495,n7577);
  nand U8887(n8536,G26,n8496);
  nand U8888(n8535,G21454,n8497);
  nand U8889(n8534,n8498,G10);
  nand U8890(G849,n8541,n8542,n8543,n8544);
  nor U8891(n8544,n8545,n8546,n8547);
  nor U8892(n8547,n7585,n8493);
  nor U8893(n8546,n8494,n7586);
  and U8894(n8494,n8548,n8549);
  nand U8895(n8549,n8550,n7590);
  nand U8896(n8548,n8551,G21426);
  nor U8897(n8545,n8495,n7592);
  nand U8898(n8543,G25,n8496);
  nand U8899(n8496,n8552,n8553);
  nand U8900(n8553,n8550,n7595,n8495,n8554);
  not U8901(n8550,n8555);
  nand U8902(n8552,n8556,n8557);
  nand U8903(n8542,G21453,n8497);
  nand U8904(n8497,n8558,n8559);
  nand U8905(n8559,n8560,n7603,n8561);
  nand U8906(n8561,n7605,n8551);
  nand U8907(n8560,n8557,n7606);
  not U8908(n8557,n8493);
  nand U8909(n8558,n8556,n8493);
  nand U8910(n8493,n8562,n7607);
  nor U8911(n7607,G21566,G21565);
  and U8912(n8556,n8563,n8555);
  nand U8913(n8555,n8564,n7610);
  nor U8914(n7610,n8565,n8566);
  nand U8915(n8563,n7612,n8567);
  nand U8916(n8567,n8495,n8554,n7595);
  nand U8917(n8541,n8498,G9);
  and U8918(n8498,n8551,n8495,n7595);
  not U8919(n8551,n8554);
  nand U8920(G848,n8568,n8569,n8570,n8571);
  nor U8921(n8571,n8572,n8573,n8574);
  nor U8922(n8574,n7509,n8575);
  nor U8923(n8573,n8576,n7512);
  nor U8924(n8572,n8577,n7514);
  nand U8925(n8570,G32,n8578);
  nand U8926(n8569,G21452,n8579);
  nand U8927(n8568,n8580,G16);
  nand U8928(G847,n8581,n8582,n8583,n8584);
  nor U8929(n8584,n8585,n8586,n8587);
  nor U8930(n8587,n7525,n8575);
  nor U8931(n8586,n8576,n7526);
  nor U8932(n8585,n8577,n7527);
  nand U8933(n8583,G31,n8578);
  nand U8934(n8582,G21451,n8579);
  nand U8935(n8581,n8580,G15);
  nand U8936(G846,n8588,n8589,n8590,n8591);
  nor U8937(n8591,n8592,n8593,n8594);
  nor U8938(n8594,n7535,n8575);
  nor U8939(n8593,n8576,n7536);
  nor U8940(n8592,n8577,n7537);
  nand U8941(n8590,G30,n8578);
  nand U8942(n8589,G21450,n8579);
  nand U8943(n8588,n8580,G14);
  nand U8944(G845,n8595,n8596,n8597,n8598);
  nor U8945(n8598,n8599,n8600,n8601);
  nor U8946(n8601,n7545,n8575);
  nor U8947(n8600,n8576,n7546);
  nor U8948(n8599,n8577,n7547);
  nand U8949(n8597,G29,n8578);
  nand U8950(n8596,G21449,n8579);
  nand U8951(n8595,n8580,G13);
  nand U8952(G844,n8602,n8603,n8604,n8605);
  nor U8953(n8605,n8606,n8607,n8608);
  nor U8954(n8608,n7555,n8575);
  nor U8955(n8607,n8576,n7556);
  nor U8956(n8606,n8577,n7557);
  nand U8957(n8604,G28,n8578);
  nand U8958(n8603,G21448,n8579);
  nand U8959(n8602,n8580,G12);
  nand U8960(G843,n8609,n8610,n8611,n8612);
  nor U8961(n8612,n8613,n8614,n8615);
  nor U8962(n8615,n7565,n8575);
  nor U8963(n8614,n8576,n7566);
  nor U8964(n8613,n8577,n7567);
  nand U8965(n8611,G27,n8578);
  nand U8966(n8610,G21447,n8579);
  nand U8967(n8609,n8580,G11);
  nand U8968(G842,n8616,n8617,n8618,n8619);
  nor U8969(n8619,n8620,n8621,n8622);
  nor U8970(n8622,n7575,n8575);
  nor U8971(n8621,n8576,n7576);
  nor U8972(n8620,n8577,n7577);
  nand U8973(n8618,G26,n8578);
  nand U8974(n8617,G21446,n8579);
  nand U8975(n8616,n8580,G10);
  nand U8976(G841,n8623,n8624,n8625,n8626);
  nor U8977(n8626,n8627,n8628,n8629);
  nor U8978(n8629,n7585,n8575);
  nor U8979(n8628,n8576,n7586);
  and U8980(n8576,n8630,n8631);
  nand U8981(n8631,n8632,n7590);
  nand U8982(n8630,n8633,G21426);
  nor U8983(n8627,n8577,n7592);
  nand U8984(n8625,G25,n8578);
  nand U8985(n8578,n8634,n8635);
  nand U8986(n8635,n8632,n7595,n8577,n8636);
  not U8987(n8632,n8637);
  nand U8988(n8634,n8638,n8639);
  nand U8989(n8624,G21445,n8579);
  nand U8990(n8579,n8640,n8641);
  nand U8991(n8641,n8642,n7603,n8643);
  nand U8992(n8643,n7605,n8633);
  nand U8993(n8642,n8639,n7606);
  not U8994(n8639,n8575);
  nand U8995(n8640,n8638,n8575);
  nand U8996(n8575,n8562,n7690);
  and U8997(n8638,n8644,n8637);
  nand U8998(n8637,n8564,n7692);
  nor U8999(n7692,n8565,G21566);
  nand U9000(n8644,n7612,n8645);
  nand U9001(n8645,n8577,n8636,n7595);
  nand U9002(n8623,n8580,G9);
  and U9003(n8580,n8633,n8577,n7595);
  not U9004(n8633,n8636);
  nand U9005(G840,n8646,n8647,n8648,n8649);
  nor U9006(n8649,n8650,n8651,n8652);
  nor U9007(n8652,n7509,n8653);
  nor U9008(n8651,n8654,n7512);
  nor U9009(n8650,n8655,n7514);
  nand U9010(n8648,G32,n8656);
  nand U9011(n8647,G21444,n8657);
  nand U9012(n8646,n8658,G16);
  nand U9013(G839,n8659,n8660,n8661,n8662);
  nor U9014(n8662,n8663,n8664,n8665);
  nor U9015(n8665,n7525,n8653);
  nor U9016(n8664,n8654,n7526);
  nor U9017(n8663,n8655,n7527);
  nand U9018(n8661,G31,n8656);
  nand U9019(n8660,G21443,n8657);
  nand U9020(n8659,n8658,G15);
  nand U9021(G838,n8666,n8667,n8668,n8669);
  nor U9022(n8669,n8670,n8671,n8672);
  nor U9023(n8672,n7535,n8653);
  nor U9024(n8671,n8654,n7536);
  nor U9025(n8670,n8655,n7537);
  nand U9026(n8668,G30,n8656);
  nand U9027(n8667,G21442,n8657);
  nand U9028(n8666,n8658,G14);
  nand U9029(G837,n8673,n8674,n8675,n8676);
  nor U9030(n8676,n8677,n8678,n8679);
  nor U9031(n8679,n7545,n8653);
  nor U9032(n8678,n8654,n7546);
  nor U9033(n8677,n8655,n7547);
  nand U9034(n8675,G29,n8656);
  nand U9035(n8674,G21441,n8657);
  nand U9036(n8673,n8658,G13);
  nand U9037(G836,n8680,n8681,n8682,n8683);
  nor U9038(n8683,n8684,n8685,n8686);
  nor U9039(n8686,n7555,n8653);
  nor U9040(n8685,n8654,n7556);
  nor U9041(n8684,n8655,n7557);
  nand U9042(n8682,G28,n8656);
  nand U9043(n8681,G21440,n8657);
  nand U9044(n8680,n8658,G12);
  nand U9045(G835,n8687,n8688,n8689,n8690);
  nor U9046(n8690,n8691,n8692,n8693);
  nor U9047(n8693,n7565,n8653);
  nor U9048(n8692,n8654,n7566);
  nor U9049(n8691,n8655,n7567);
  nand U9050(n8689,G27,n8656);
  nand U9051(n8688,G21439,n8657);
  nand U9052(n8687,n8658,G11);
  nand U9053(G834,n8694,n8695,n8696,n8697);
  nor U9054(n8697,n8698,n8699,n8700);
  nor U9055(n8700,n7575,n8653);
  nor U9056(n8699,n8654,n7576);
  nor U9057(n8698,n8655,n7577);
  nand U9058(n8696,G26,n8656);
  nand U9059(n8695,G21438,n8657);
  nand U9060(n8694,n8658,G10);
  nand U9061(G833,n8701,n8702,n8703,n8704);
  nor U9062(n8704,n8705,n8706,n8707);
  nor U9063(n8707,n7585,n8653);
  nor U9064(n8706,n8654,n7586);
  and U9065(n8654,n8708,n8709);
  nand U9066(n8709,n8710,n7590);
  nand U9067(n8708,n8711,G21426);
  nor U9068(n8705,n8655,n7592);
  nand U9069(n8703,G25,n8656);
  nand U9070(n8656,n8712,n8713);
  nand U9071(n8713,n8710,n7595,n8655,n8714);
  not U9072(n8710,n8715);
  nand U9073(n8712,n8716,n8717);
  nand U9074(n8702,G21437,n8657);
  nand U9075(n8657,n8718,n8719);
  nand U9076(n8719,n8720,n7603,n8721);
  nand U9077(n8721,n7605,n8711);
  nand U9078(n8720,n8717,n7606);
  not U9079(n8717,n8653);
  nand U9080(n8718,n8716,n8653);
  nand U9081(n8653,n8562,n7770);
  and U9082(n8716,n8722,n8715);
  nand U9083(n8715,n8564,n7772);
  nor U9084(n7772,n8566,n8723);
  nand U9085(n8722,n7612,n8724);
  nand U9086(n8724,n8655,n8714,n7595);
  nand U9087(n8701,n8658,G9);
  and U9088(n8658,n8711,n8655,n7595);
  not U9089(n8711,n8714);
  nand U9090(G832,n8725,n8726,n8727,n8728);
  nor U9091(n8728,n8729,n8730,n8731);
  nor U9092(n8731,n8732,n7514);
  nand U9093(n7514,G8,n7595);
  nor U9094(n8730,n7509,n8733);
  and U9095(n7509,n8734,n8735);
  or U9096(n8735,n7512,n7456);
  nand U9097(n8734,n8736,n8737);
  nor U9098(n8729,n8738,n7512);
  nand U9099(n7512,G32,n7606);
  nand U9100(n8727,G32,n8739);
  nand U9101(n8726,G21436,n8740);
  nand U9102(n8725,n8741,G16);
  nand U9103(G831,n8742,n8743,n8744,n8745);
  nor U9104(n8745,n8746,n8747,n8748);
  nor U9105(n8748,n8732,n7527);
  nand U9106(n7527,G7,n7595);
  nor U9107(n8747,n7525,n8733);
  and U9108(n7525,n8749,n8750);
  or U9109(n8750,n7526,n7456);
  nand U9110(n8749,n8736,n7470);
  nor U9111(n8746,n8738,n7526);
  nand U9112(n7526,G31,n7606);
  nand U9113(n8744,G31,n8739);
  nand U9114(n8743,G21435,n8740);
  nand U9115(n8742,n8741,G15);
  nand U9116(G830,n8751,n8752,n8753,n8754);
  nor U9117(n8754,n8755,n8756,n8757);
  nor U9118(n8757,n8732,n7537);
  nand U9119(n7537,G6,n7595);
  nor U9120(n8756,n7535,n8733);
  and U9121(n7535,n8758,n8759);
  or U9122(n8759,n7536,n7456);
  nand U9123(n8758,n8736,n7482);
  nor U9124(n8755,n8738,n7536);
  nand U9125(n7536,G30,n7606);
  nand U9126(n8753,G30,n8739);
  nand U9127(n8752,G21434,n8740);
  nand U9128(n8751,n8741,G14);
  nand U9129(G829,n8760,n8761,n8762,n8763);
  nor U9130(n8763,n8764,n8765,n8766);
  nor U9131(n8766,n8732,n7547);
  nand U9132(n7547,G5,n7595);
  nor U9133(n8765,n7545,n8733);
  and U9134(n7545,n8767,n8768);
  or U9135(n8768,n7546,n7456);
  nand U9136(n8767,n8736,n8769);
  nor U9137(n8764,n8738,n7546);
  nand U9138(n7546,G29,n7606);
  nand U9139(n8762,G29,n8739);
  nand U9140(n8761,G21433,n8740);
  nand U9141(n8760,n8741,G13);
  nand U9142(G828,n8770,n8771,n8772,n8773);
  nor U9143(n8773,n8774,n8775,n8776);
  nor U9144(n8776,n8732,n7557);
  nand U9145(n7557,G4,n7595);
  nor U9146(n8775,n7555,n8733);
  and U9147(n7555,n8777,n8778);
  or U9148(n8778,n7556,n7456);
  nand U9149(n8777,n8736,n7484);
  nor U9150(n8774,n8738,n7556);
  nand U9151(n7556,G28,n7606);
  nand U9152(n8772,G28,n8739);
  nand U9153(n8771,G21432,n8740);
  nand U9154(n8770,n8741,G12);
  nand U9155(G827,n8779,n8780,n8781,n8782);
  nor U9156(n8782,n8783,n8784,n8785);
  nor U9157(n8785,n8732,n7567);
  nand U9158(n7567,G3,n7595);
  nor U9159(n8784,n7565,n8733);
  and U9160(n7565,n8786,n8787);
  or U9161(n8787,n7566,n7456);
  nand U9162(n8786,n8736,n8788);
  nor U9163(n8783,n8738,n7566);
  nand U9164(n7566,G27,n7606);
  nand U9165(n8781,G27,n8739);
  nand U9166(n8780,G21431,n8740);
  nand U9167(n8779,n8741,G11);
  nand U9168(G826,n8789,n8790,n8791,n8792);
  nor U9169(n8792,n8793,n8794,n8795);
  nor U9170(n8795,n8732,n7577);
  nand U9171(n7577,G2,n7595);
  nor U9172(n8794,n7575,n8733);
  and U9173(n7575,n8796,n8797);
  or U9174(n8797,n7576,n7456);
  nand U9175(n8796,n8736,n8798);
  nor U9176(n8793,n8738,n7576);
  nand U9177(n7576,G26,n7606);
  nand U9178(n8791,G26,n8739);
  nand U9179(n8790,G21430,n8740);
  nand U9180(n8789,n8741,G10);
  nand U9181(G825,n8799,n8800,n8801,n8802);
  nor U9182(n8802,n8803,n8804,n8805);
  nor U9183(n8805,n8732,n7592);
  nand U9184(n7592,G1,n7595);
  nor U9185(n8804,n7585,n8733);
  and U9186(n7585,n8806,n8807);
  nand U9187(n8807,n8736,n8808);
  nor U9188(n8736,n8809,n8810);
  or U9189(n8806,n7586,n7456);
  nor U9190(n8803,n8738,n7586);
  nand U9191(n7586,G25,n7606);
  and U9192(n8738,n8811,n8812);
  nand U9193(n8812,n8813,n7590);
  nand U9194(n8811,n8814,G21426);
  nand U9195(n8801,G25,n8739);
  nand U9196(n8739,n8815,n8816);
  nand U9197(n8816,n7595,n8732,n8813);
  not U9198(n8813,n8817);
  nand U9199(n8815,n8818,n8819);
  nand U9200(n8800,G21429,n8740);
  nand U9201(n8740,n8820,n8821);
  nand U9202(n8821,n8822,n7603,n8823);
  nand U9203(n8823,n8819,n7606);
  not U9204(n8819,n8733);
  nand U9205(n7603,n7605,n7456);
  nand U9206(n8822,n7605,n8814);
  nor U9207(n7605,n8810,n8824);
  nand U9208(n8820,n8818,n8733);
  nand U9209(n8733,n8562,n7850);
  nor U9210(n8562,n8825,n8826);
  and U9211(n8818,n8827,n8817);
  nand U9212(n8817,n8564,n7852);
  nor U9213(n7852,G21566,n8723);
  nor U9214(n8564,n8169,n8170);
  nand U9215(n8827,n7612,n8828);
  nand U9216(n8828,n8732,n8829,n7595);
  nand U9217(n7612,n7590,n7606);
  nand U9218(n8799,n8741,G9);
  and U9219(n8741,n7595,n8814);
  not U9220(n8814,n8829);
  nand U9221(G824,n8831,n8832,n8833,n8834);
  nand U9222(n8834,n8835,G21428);
  nand U9223(n8833,n8836,n8837);
  nand U9224(n8836,n8838,n8839,n8840);
  nand U9225(n8840,n8841,n7483);
  nand U9226(n8839,n8842,n8843);
  nand U9227(n8842,G21425,n7483,n8824);
  nand U9228(n8838,n8844,n8845);
  nand U9229(G823,n8846,n8847,n8848);
  nand U9230(n8848,G21427,n8849);
  nand U9231(n8849,n8837,n8832);
  nand U9232(n8832,G21428,n7456,G35);
  nand U9233(n8846,n8850,n8837);
  nand U9234(n8850,n8851,n8852);
  nand U9235(n8852,G21428,n7471,n8853);
  not U9236(n8851,n7459);
  nand U9237(G822,n8854,n8855,n8856,n8857);
  or U9238(n8857,n8830,G21428);
  nand U9239(n8856,n7456,n7471,G21427,G21428);
  nand U9240(G821,n8858,n8859,n8860);
  nand U9241(n8860,n8835,G21425);
  not U9242(n8835,n8837);
  nand U9243(n8837,n8861,n8862,n8863,n8864);
  nand U9244(n8864,n8843,n7471);
  nand U9245(n8863,G21428,n8865);
  or U9246(n8865,n8845,G21427);
  nand U9247(n8845,n8866,n7453,n8867,n8868);
  nor U9248(n8868,n8869,n8870,n8871,n8872);
  nor U9249(n8872,n7450,n8873);
  nor U9250(n8871,n8874,n8875);
  nor U9251(n8870,n7467,n7455);
  nor U9252(n8869,n8876,n8877);
  nor U9253(n8867,n8878,n8879);
  nor U9254(n8879,n8880,n7483);
  nor U9255(n8880,n8881,n8882,n8883);
  nor U9256(n8883,n8737,n8884);
  nor U9257(n8878,n8885,n8886);
  nor U9258(n8885,G21795,G21796);
  not U9259(n7453,n8887);
  nand U9260(n8866,n8888,n7500,n8889);
  nand U9261(n8889,G21563,n8877);
  nand U9262(n8888,n8890,n8891,n8892);
  or U9263(n8892,n8877,G21563);
  nand U9264(n8877,n8893,n8894);
  nand U9265(n8894,n8895,n8896);
  or U9266(n8893,n8897,n8895);
  nand U9267(n8891,n8898,n8899,n8900);
  nand U9268(n8900,G21564,n8876);
  nand U9269(n8899,n8901,n8875);
  nand U9270(n8901,n8902,n8903);
  nand U9271(n8903,n8904,n8905);
  nand U9272(n8905,n8906,n8907);
  nand U9273(n8907,n8908,G21566);
  not U9274(n8904,n8909);
  nand U9275(n8902,n8908,n7850);
  not U9276(n8908,n8910);
  nand U9277(n8898,n8895,n8911);
  nand U9278(n8911,n8912,n8913,n8914);
  nand U9279(n8914,G21566,n8915);
  nand U9280(n8912,n7850,n8916);
  or U9281(n8890,n8876,G21564);
  nand U9282(n8876,n8917,n8918);
  nand U9283(n8918,n8895,n8919);
  or U9284(n8917,n8920,n8895);
  not U9285(n8895,n8875);
  nand U9286(n8862,n8921,n8882);
  nand U9287(n8861,n8922,n8923);
  not U9288(n8859,n8924);
  nor U9289(G820,n8925,n8926);
  nor U9290(G819,n8925,n8927);
  nor U9291(G818,n8925,n8928);
  nor U9292(G817,n8925,n8929);
  nor U9293(G816,n8925,n8930);
  nor U9294(G815,n8925,n8931);
  nor U9295(G814,n8925,n8932);
  nor U9296(G813,n8925,n8933);
  nor U9297(G812,n8925,n8934);
  nor U9298(G811,n8925,n8935);
  nor U9299(G810,n8925,n8936);
  nor U9300(G809,n8925,n8937);
  nor U9301(G808,n8925,n8938);
  nor U9302(G807,n8925,n8939);
  nor U9303(G806,n8925,n8940);
  nor U9304(G805,n8925,n8941);
  and U9305(G804,n8942,G21408);
  and U9306(G803,n8942,G21407);
  and U9307(G802,n8942,G21406);
  and U9308(G801,n8942,G21405);
  and U9309(G800,n8942,G21404);
  and U9310(G799,n8942,G21403);
  and U9311(G798,n8942,G21402);
  and U9312(G797,n8942,G21401);
  nor U9313(G796,n8925,n8943);
  nor U9314(G795,n8925,n8944);
  nor U9315(G794,n8925,n8945);
  nor U9316(G793,n8925,n8946);
  and U9317(G792,n8942,G21396);
  and U9318(G791,n8942,G21395);
  nand U9319(G790,n8947,n8948,n8949);
  nor U9320(n8949,n8950,n8951,n8952);
  nor U9321(n8952,n8953,G21392,G21391);
  nor U9322(n8950,G21798,n8954);
  or U9323(n8948,n8955,n8956);
  nand U9324(n8947,n8957,n8958);
  nand U9325(G789,n8959,n8960,n8961,n8962);
  nand U9326(n8962,n8963,n8964);
  nand U9327(n8963,n8965,n8966);
  nand U9328(n8966,G21392,n8967,G21798);
  nand U9329(n8961,n8968,n8965,n8969,G21391);
  nand U9330(n8969,n8956,n8970);
  nand U9331(n8968,n8957,n7471);
  not U9332(n8957,n8967);
  nand U9333(n8967,G36,G21390);
  not U9334(n8960,n8971);
  nand U9335(n8959,n8972,G35);
  nand U9336(G787,n8973,n8974,n8975,n8976);
  not U9337(n8976,n8954);
  nand U9338(n8975,G21392,n8977,G36);
  nand U9339(n8977,n8978,n8979,n8980);
  nand U9340(n8979,n8964,n8970);
  nand U9341(n8978,G35,n8953,G21391);
  or U9342(n8974,n8980,n8956,n8964);
  nor U9343(n8956,G36,G35);
  nand U9344(n8973,n8981,n8953);
  not U9345(n8953,G33);
  nand U9346(n8981,n8965,n8982);
  nand U9347(n8982,G21798,G35,n8983);
  nand U9348(n8965,G21390,n8984);
  nand U9349(G786,n8985,n8986,n8987);
  nand U9350(n8987,G21389,n8958);
  nand U9351(n8986,n8954,G21759);
  nand U9352(n8985,n8971,G21760);
  nand U9353(G785,n8988,n8989,n8990);
  nand U9354(n8990,G21388,n8958);
  nand U9355(n8989,n8954,G21760);
  nand U9356(n8988,n8971,G21761);
  nand U9357(G784,n8991,n8992,n8993);
  nand U9358(n8993,G21387,n8958);
  nand U9359(n8992,n8954,G21761);
  nand U9360(n8991,n8971,G21762);
  nand U9361(G783,n8994,n8995,n8996);
  nand U9362(n8996,G21386,n8958);
  nand U9363(n8995,n8954,G21762);
  nand U9364(n8994,n8971,G21763);
  nand U9365(G782,n8997,n8998,n8999);
  nand U9366(n8999,G21385,n8958);
  nand U9367(n8998,n8954,G21763);
  nand U9368(n8997,n8971,G21764);
  nand U9369(G781,n9000,n9001,n9002);
  nand U9370(n9002,G21384,n8958);
  nand U9371(n9001,n8954,G21764);
  nand U9372(n9000,n8971,G21765);
  nand U9373(G780,n9003,n9004,n9005);
  nand U9374(n9005,G21383,n8958);
  nand U9375(n9004,n8954,G21765);
  nand U9376(n9003,n8971,G21766);
  nand U9377(G779,n9006,n9007,n9008);
  nand U9378(n9008,G21382,n8958);
  nand U9379(n9007,n8954,G21766);
  nand U9380(n9006,n8971,G21767);
  nand U9381(G778,n9009,n9010,n9011);
  nand U9382(n9011,G21381,n8958);
  nand U9383(n9010,n8954,G21767);
  nand U9384(n9009,n8971,G21768);
  nand U9385(G777,n9012,n9013,n9014);
  nand U9386(n9014,G21380,n8958);
  nand U9387(n9013,n8954,G21768);
  nand U9388(n9012,n8971,G21769);
  nand U9389(G776,n9015,n9016,n9017);
  nand U9390(n9017,G21379,n8958);
  nand U9391(n9016,n8954,G21769);
  nand U9392(n9015,n8971,G21770);
  nand U9393(G775,n9018,n9019,n9020);
  nand U9394(n9020,G21378,n8958);
  nand U9395(n9019,n8954,G21770);
  nand U9396(n9018,n8971,G21771);
  nand U9397(G774,n9021,n9022,n9023);
  nand U9398(n9023,G21377,n8958);
  nand U9399(n9022,n8954,G21771);
  nand U9400(n9021,n8971,G21772);
  nand U9401(G773,n9024,n9025,n9026);
  nand U9402(n9026,G21376,n8958);
  nand U9403(n9025,n8954,G21772);
  nand U9404(n9024,n8971,G21773);
  nand U9405(G772,n9027,n9028,n9029);
  nand U9406(n9029,G21375,n8958);
  nand U9407(n9028,n8954,G21773);
  nand U9408(n9027,n8971,G21774);
  nand U9409(G771,n9030,n9031,n9032);
  nand U9410(n9032,G21374,n8958);
  nand U9411(n9031,n8954,G21774);
  nand U9412(n9030,n8971,G21775);
  nand U9413(G770,n9033,n9034,n9035);
  nand U9414(n9035,G21373,n8958);
  nand U9415(n9034,n8954,G21775);
  nand U9416(n9033,n8971,G21776);
  nand U9417(G769,n9036,n9037,n9038);
  nand U9418(n9038,G21372,n8958);
  nand U9419(n9037,n8954,G21776);
  nand U9420(n9036,n8971,G21777);
  nand U9421(G768,n9039,n9040,n9041);
  nand U9422(n9041,G21371,n8958);
  nand U9423(n9040,n8954,G21777);
  nand U9424(n9039,n8971,G21778);
  nand U9425(G767,n9042,n9043,n9044);
  nand U9426(n9044,G21370,n8958);
  nand U9427(n9043,n8954,G21778);
  nand U9428(n9042,n8971,G21779);
  nand U9429(G766,n9045,n9046,n9047);
  nand U9430(n9047,G21369,n8958);
  nand U9431(n9046,n8954,G21779);
  nand U9432(n9045,n8971,G21780);
  nand U9433(G765,n9048,n9049,n9050);
  nand U9434(n9050,G21368,n8958);
  nand U9435(n9049,n8954,G21780);
  nand U9436(n9048,n8971,G21781);
  nand U9437(G764,n9051,n9052,n9053);
  nand U9438(n9053,G21367,n8958);
  nand U9439(n9052,n8954,G21781);
  nand U9440(n9051,n8971,G21782);
  nand U9441(G763,n9054,n9055,n9056);
  nand U9442(n9056,G21366,n8958);
  nand U9443(n9055,n8954,G21782);
  nand U9444(n9054,n8971,G21783);
  nand U9445(G762,n9057,n9058,n9059);
  nand U9446(n9059,G21365,n8958);
  nand U9447(n9058,n8954,G21783);
  nand U9448(n9057,n8971,G21784);
  nand U9449(G761,n9060,n9061,n9062);
  nand U9450(n9062,G21364,n8958);
  nand U9451(n9061,n8954,G21784);
  nand U9452(n9060,n8971,G21785);
  nand U9453(G760,n9063,n9064,n9065);
  nand U9454(n9065,G21363,n8958);
  nand U9455(n9064,n8954,G21785);
  nand U9456(n9063,n8971,G21786);
  nand U9457(G759,n9066,n9067,n9068);
  nand U9458(n9068,G21362,n8958);
  nand U9459(n9067,n8954,G21786);
  nand U9460(n9066,n8971,G21787);
  nand U9461(G758,n9069,n9070,n9071);
  nand U9462(n9071,G21361,n8958);
  nand U9463(n9070,n8954,G21787);
  nand U9464(n9069,n8971,G21788);
  nand U9465(G757,n9072,n9073,n9074);
  nand U9466(n9074,G21360,n8958);
  nand U9467(n9073,n8954,G21788);
  nand U9468(n9072,n8971,G21789);
  nand U9469(G1751,n9075,n9076);
  nand U9470(n9076,G21804,n9077);
  nand U9471(n9075,n9078,n9079);
  nand U9472(G1750,n9080,n9081);
  nand U9473(n9081,n9077,G21803);
  or U9474(n9080,n9082,n9077);
  not U9475(n9077,n9079);
  nand U9476(n9079,n9083,n9084);
  nand U9477(n9084,n8824,n9085);
  nor U9478(n9082,n9086,n9087,n7456);
  nand U9479(G1749,n9088,n9089);
  nand U9480(n9089,G21800,n8958);
  nand U9481(n9088,G21804,n8972);
  nand U9482(G1748,n9090,n9091);
  or U9483(n9091,n9092,n8970);
  not U9484(n8970,G21798);
  nand U9485(n9090,n9093,n9092);
  nand U9486(n9092,n9094,n9095,n9083);
  nand U9487(n9095,n8923,n9085,n8922);
  nand U9488(n8922,G21428,G21426);
  nand U9489(n9094,G21427,n7471,n9096);
  nand U9490(n9093,n8809,n9097);
  nand U9491(n9097,G21428,n9098);
  nand U9492(n9098,G21426,n9099,n9100,n7471);
  or U9493(n9100,n9101,G21797,n7470);
  or U9494(n9099,n7480,n9102);
  nand U9495(G1747,n9103,n9104);
  or U9496(n9104,n8958,G21803);
  nand U9497(n9103,G21794,n8958);
  nand U9498(G1746,n9105,n9106,n9107,n9108);
  nand U9499(n9108,G21428,n7483,n7501);
  nand U9500(n9107,n7488,G21566);
  nand U9501(n9106,n9109,n7456,n7489);
  nor U9502(n7489,n9110,n7488);
  not U9503(n7488,n7501);
  nand U9504(n9105,n7491,n7031);
  and U9505(n7491,n9111,n7501);
  nand U9506(n7501,n9112,n9113,n8810);
  not U9507(n8810,n7606);
  nand U9508(n7606,n9114,n9115,n9116);
  or U9509(n9116,n8858,n9117);
  nand U9510(n9115,n9096,n9118);
  nand U9511(n9114,n7456,n8843,G21427);
  nand U9512(n9112,n8924,n9117);
  nand U9513(n9111,n8855,n9119);
  nand U9514(n9119,n9110,n7456);
  nand U9515(G1745,n9120,n9121);
  nand U9516(n9121,n9122,G21561);
  nand U9517(n9120,n9123,n9124);
  nand U9518(n9123,n9125,n9126,n9127);
  nand U9519(n9127,n8844,n8910);
  nand U9520(n8910,n9128,n9129,n9130);
  nor U9521(n9130,n9131,n9132,n9133);
  nor U9522(n9133,n9134,n9135);
  and U9523(n9132,n8916,n8881);
  nor U9524(n9131,n9136,n9137);
  nand U9525(n9129,n7031,n9138);
  nand U9526(n9128,n7033,n9139);
  nand U9527(n9126,G21427,n9140);
  nand U9528(n9140,G21567,n9137);
  nand U9529(n9125,n9141,n7033);
  nand U9530(G1744,n9142,n9143);
  nand U9531(n9143,n9122,G21560);
  nand U9532(n9142,n9144,n9124);
  nand U9533(n9144,n9145,n9146,n9147);
  nand U9534(n9147,n9148,n9149);
  nand U9535(n9146,n9141,n7022);
  nand U9536(n9145,n8844,n8909);
  nand U9537(n8909,n9150,n9151,n9152,n9153);
  nor U9538(n9153,n9154,n9155,n9156);
  nor U9539(n9156,n9134,n9157);
  nor U9540(n9155,n9158,n9159);
  nor U9541(n9158,n9160,n9161);
  nor U9542(n9154,n9136,n9162);
  nand U9543(n9152,n9163,n9164);
  nand U9544(n9151,n7020,n9138);
  nand U9545(n9150,n7022,n9139);
  nand U9546(G1743,n9165,n9166);
  nand U9547(n9166,n9122,G21559);
  nand U9548(n9165,n9167,n9124);
  nand U9549(n9167,n9168,n9169,n9170);
  nand U9550(n9170,n9148,n9171);
  nand U9551(n9169,n9141,n7011);
  nand U9552(n9168,n8844,n8920);
  nand U9553(n8920,n9172,n9173,n9174,n9175);
  nor U9554(n9175,n9176,n9177,n9178);
  nor U9555(n9178,n9136,n9179);
  nor U9556(n9177,n9134,n9180);
  nor U9557(n9176,n9181,n7418);
  nand U9558(n9174,n9163,n9182);
  nand U9559(n9173,n9139,n7011);
  nand U9560(n9172,n9183,n7446);
  nand U9561(G1742,n9184,n9185);
  nand U9562(n9185,n9122,G21558);
  nand U9563(n9184,n9186,n9124);
  nand U9564(n9186,n9187,n9188);
  nand U9565(n9188,n9141,n7001);
  nor U9566(n9141,n9117,G21426);
  nand U9567(n9187,n8844,n8897);
  nand U9568(n8897,n9189,n9190,n9191,n9192);
  nor U9569(n9192,n9193,n9194,n9195);
  nor U9570(n9195,n9136,n9196);
  and U9571(n9136,n9197,n7455);
  nor U9572(n9194,n9134,n9198);
  nor U9573(n9134,n9199,n9200);
  nor U9574(n9193,n9181,n9201);
  not U9575(n9181,n9138);
  nand U9576(n9138,n7439,n7440,n9202);
  nor U9577(n9202,n9203,n7444,n7445);
  nor U9578(n7445,n8808,n7482,n7470,n9101);
  nor U9579(n9203,n7477,n9204);
  and U9580(n7440,n9205,n9206,n9207,n9208);
  nand U9581(n9208,n9209,n8808);
  nand U9582(n9207,n9210,n7484);
  nand U9583(n9206,n7470,n8737,n7482);
  and U9584(n7439,n9211,n9212,n9213);
  nand U9585(n9213,n7472,n9214);
  nand U9586(n9214,n9215,n9216);
  nand U9587(n9215,n9217,n9218);
  nand U9588(n9212,n9101,n9219);
  nand U9589(n9191,n9220,n9163);
  nand U9590(n9190,n7001,n9139);
  nand U9591(n9139,n9221,n9222,n7452,n7450);
  nand U9592(n9222,n9223,n7484);
  nand U9593(n9223,n9224,n9225);
  nand U9594(n9225,n9226,n9227);
  nand U9595(n9189,n7446,n9228);
  not U9596(n7446,n9159);
  nand U9597(G1740,n9229,n9230);
  nand U9598(n9230,n6990,n9231,n8844,n9124);
  nand U9599(n9229,n9122,G21557);
  not U9600(n9122,n9124);
  nand U9601(n9124,n8858,n9113,n9232);
  nand U9602(n9232,n7459,n8875);
  nand U9603(n8875,n7461,n9233,n9234,n9235);
  nand U9604(n9235,n7467,n7471,n9236);
  nand U9605(n9234,n7473,n9237);
  nand U9606(n9237,n7450,n9238);
  nand U9607(n9238,n7480,n9239);
  nand U9608(n9239,n9211,n9240);
  nand U9609(n9233,n7483,n8881);
  nand U9610(n8881,n7454,n9159);
  and U9611(n7461,n9241,n9242,n9243,n9244);
  nor U9612(n9244,n9245,n9246);
  or U9613(n9246,n9247,n7481);
  nand U9614(n9241,n9248,n7472);
  nand U9615(n9113,n8924,G21795);
  nor U9616(n8924,n8923,n8843);
  nand U9617(n8858,G21425,n8843);
  nand U9618(G1738,n9249,n9250);
  nand U9619(n9250,G21394,n8942);
  nand U9620(n9249,n9251,n8925);
  nand U9621(n9251,n9252,n9253);
  nand U9622(G1737,n9254,n9255);
  nand U9623(n9255,n9253,n9252,n8925);
  not U9624(n9252,G34);
  not U9625(n9253,n8951);
  nand U9626(n9254,G21393,n8942);
  nand U9627(G1735,n9256,n9257);
  nand U9628(n9257,G21359,n8958);
  nand U9629(n9256,G21793,n8972);
  nand U9630(G1734,n9258,n9259);
  nand U9631(n9259,G21358,n8958);
  nand U9632(n9258,G21792,n8972);
  nand U9633(G1733,n9260,n9261);
  nand U9634(n9261,G21357,n8958);
  nand U9635(n9260,G21791,n8972);
  nand U9636(G1732,n9262,n9263);
  nand U9637(n9263,G21356,n8958);
  nand U9638(n9262,G21790,n8972);
  nand U9639(G1189,n8942,n9264);
  nand U9640(n9264,G21802,G21392);
  nand U9641(G1188,n9265,n9266);
  nand U9642(n9266,G21428,n9085,n8824);
  nand U9643(n9265,G21801,n9267);
  nand U9644(n9267,n9268,n7459);
  nand U9645(G1187,n9269,n9270,n9271);
  or U9646(n9270,n8958,G21801);
  nand U9647(n9269,G21799,n8958);
  nor U9648(n8972,n8964,G21392);
  nand U9649(G1186,n9272,n9273,n9271);
  nand U9650(n9271,n8951,n8964);
  nor U9651(n8951,G21392,G21390);
  nand U9652(n9273,G34,n8925);
  not U9653(n8925,n8942);
  nand U9654(n9272,n8942,G21797);
  nor U9655(n8942,n9274,n8983);
  nor U9656(n8983,n8984,n8955);
  nor U9657(n9274,G21392,G21391);
  nand U9658(G1185,n9275,n9276);
  nand U9659(n9276,n9277,n8886);
  nand U9660(n9277,n9278,n9279);
  nand U9661(n9279,n9280,n9281);
  nand U9662(n9280,n9282,n9283);
  nand U9663(n9283,n8844,n9284);
  nand U9664(n9278,n9117,n9285);
  nand U9665(n9285,n9286,n9287,n9288);
  nand U9666(n9288,n7459,n8882);
  nand U9667(n9286,n8844,n9289);
  nand U9668(n9289,n9290,n9291);
  nand U9669(n9275,G21796,n9292);
  nand U9670(G1184,n9293,n9294);
  nand U9671(n9294,G21795,n9292);
  nand U9672(n9292,n7459,n8886);
  nand U9673(n8886,n9268,n9295);
  nand U9674(n9295,n9296,n7471);
  nand U9675(n9296,n9297,n9298);
  or U9676(n9297,n7477,n7465);
  and U9677(n9268,n9299,n9300,n9301,n9302);
  nand U9678(n9301,n7465,n9303);
  nand U9679(n9303,n7481,n9304,n9305);
  nand U9680(n9304,n7470,n9281);
  nand U9681(n9300,n9117,n9306);
  nand U9682(n9306,n7465,n7470);
  not U9683(n9299,n9245);
  nand U9684(n9245,n8808,n9307,n9308);
  nand U9685(n9308,n7482,n9309);
  nand U9686(n9309,n9310,n9101);
  nand U9687(G1183,n9311,n9312,n9313);
  nand U9688(n9312,G21793,n9314);
  or U9689(n9311,n9314,n7030);
  nand U9690(G1182,n9313,n9315,n9316);
  nand U9691(n9316,G21792,n9314);
  not U9692(n9313,n9317);
  nand U9693(G1181,n9318,n9319,n9320);
  nand U9694(n9320,G21791,n9314);
  nand U9695(n9319,n9321,n7019,n9322);
  nand U9696(n9321,G21393,G21758);
  nand U9697(n9318,n9317,G21758);
  nor U9698(n9317,n9314,n7019);
  nand U9699(G1180,n9323,n9315,n9324);
  nand U9700(n9324,G21790,n9314);
  nand U9701(n9315,n9325,n7030,n9322);
  not U9702(n9325,G21393);
  nand U9703(n9323,n9322,n7019);
  nor U9704(n9322,n9314,G21394);
  nand U9705(n9314,n9326,n9327,n9328,n9329);
  nor U9706(n9329,n9330,n9331,n9332,n9333);
  nand U9707(n9333,n8941,n8940,n8939,n8938);
  not U9708(n8938,G21412);
  not U9709(n8939,G21411);
  not U9710(n8940,G21410);
  not U9711(n8941,G21409);
  nand U9712(n9332,n8937,n8936,n8935,n8934);
  not U9713(n8934,G21416);
  not U9714(n8935,G21415);
  not U9715(n8936,G21414);
  not U9716(n8937,G21413);
  nand U9717(n9331,n8933,n8932,n8931,n8930);
  not U9718(n8930,G21420);
  not U9719(n8931,G21419);
  not U9720(n8932,G21418);
  not U9721(n8933,G21417);
  nand U9722(n9330,n8929,n8928,n8927,n8926);
  not U9723(n8926,G21424);
  not U9724(n8927,G21423);
  not U9725(n8928,G21422);
  not U9726(n8929,G21421);
  nor U9727(n9328,n9334,n9335,G21396,G21395);
  and U9728(n9335,G21394,G21393);
  nand U9729(n9334,n8946,n8945,n8944,n8943);
  not U9730(n8943,G21400);
  not U9731(n8944,G21399);
  not U9732(n8945,G21398);
  not U9733(n8946,G21397);
  nor U9734(n9327,G21408,G21407,G21406,G21405);
  nor U9735(n9326,G21404,G21403,G21402,G21401);
  nand U9736(G1179,n9336,n9337,n9338,n9339);
  nor U9737(n9339,n9340,n9341,n9342);
  nor U9738(n9342,n9343,n9344);
  nor U9739(n9341,n9345,n9346);
  nor U9740(n9340,n9347,n9348);
  not U9741(n9348,n7053);
  nand U9742(n9338,n9349,G21789);
  nand U9743(n9337,n7055,n9350);
  nand U9744(n9336,n9351,n7051);
  nand U9745(G1178,n9352,n9353,n9354,n9355);
  nor U9746(n9355,n9356,n9357,n9358);
  nor U9747(n9358,n9359,n9344);
  nor U9748(n9357,n9360,n9346);
  not U9749(n9360,G21756);
  nor U9750(n9356,n9347,n7064);
  nand U9751(n9354,n9349,G21788);
  nand U9752(n9353,n9361,n9350);
  nand U9753(n9352,n9351,n7068);
  nand U9754(G1177,n9362,n9363,n9364,n9365);
  nor U9755(n9365,n9366,n9367,n9368);
  nor U9756(n9368,n9369,n9344);
  nor U9757(n9367,n9370,n9346);
  not U9758(n9370,G21755);
  nor U9759(n9366,n9347,n7077);
  nand U9760(n9364,n9349,G21787);
  nand U9761(n9363,n9371,n9350);
  nand U9762(n9362,n9351,n7081);
  nand U9763(G1176,n9372,n9373,n9374,n9375);
  nor U9764(n9375,n9376,n9377,n9378);
  nor U9765(n9378,n9379,n9344);
  nor U9766(n9377,n9380,n9346);
  not U9767(n9380,G21754);
  nor U9768(n9376,n9347,n7089);
  nand U9769(n9374,n9349,G21786);
  nand U9770(n9373,n9381,n9350);
  nand U9771(n9372,n9351,n7093);
  nand U9772(G1175,n9382,n9383,n9384,n9385);
  nor U9773(n9385,n9386,n9387,n9388);
  nor U9774(n9388,n9389,n9344);
  nor U9775(n9387,n9390,n9346);
  nor U9776(n9386,n9347,n7101);
  nand U9777(n9384,n9349,G21785);
  nand U9778(n9383,n9391,n9350);
  nand U9779(n9382,n9351,n7105);
  nand U9780(G1174,n9392,n9393,n9394,n9395);
  nor U9781(n9395,n9396,n9397,n9398);
  nor U9782(n9398,n9399,n9344);
  nor U9783(n9397,n9400,n9346);
  not U9784(n9400,G21752);
  nor U9785(n9396,n9347,n7113);
  nand U9786(n9394,n9349,G21784);
  nand U9787(n9393,n9401,n9350);
  nand U9788(n9392,n9351,n7117);
  nand U9789(G1173,n9402,n9403,n9404,n9405);
  nor U9790(n9405,n9406,n9407,n9408);
  nor U9791(n9408,n9409,n9344);
  nor U9792(n9407,n9410,n9346);
  not U9793(n9410,G21751);
  nor U9794(n9406,n9347,n9411);
  nand U9795(n9404,n9349,G21783);
  nand U9796(n9403,n7131,n9350);
  nand U9797(n9402,n9351,n7129);
  nand U9798(G1172,n9412,n9413,n9414,n9415);
  nor U9799(n9415,n9416,n9417,n9418);
  nor U9800(n9418,n9419,n9344);
  nor U9801(n9417,n9420,n9346);
  nor U9802(n9416,n9347,n7139);
  nand U9803(n9414,n9349,G21782);
  nand U9804(n9413,n9421,n9350);
  nand U9805(n9412,n9351,n7142);
  nand U9806(G1171,n9422,n9423,n9424,n9425);
  nor U9807(n9425,n9426,n9427,n9428);
  nor U9808(n9428,n9429,n9344);
  nor U9809(n9427,n9430,n9346);
  nor U9810(n9426,n9347,n9431);
  nand U9811(n9424,n9349,G21781);
  nand U9812(n9423,n7154,n9350);
  nand U9813(n9422,n9351,n7152);
  nand U9814(G1170,n9432,n9433,n9434,n9435);
  nor U9815(n9435,n9436,n9437,n9438);
  nor U9816(n9438,n9439,n9344);
  nor U9817(n9437,n9440,n9346);
  nor U9818(n9436,n9347,n9441);
  nand U9819(n9434,n9349,G21780);
  nand U9820(n9433,n7167,n9350);
  nand U9821(n9432,n9351,n7165);
  nand U9822(G1169,n9442,n9443,n9444,n9445);
  nor U9823(n9445,n9446,n9447,n9448);
  nor U9824(n9448,n9449,n9344);
  nor U9825(n9447,n9450,n9346);
  nor U9826(n9446,n9347,n9451);
  nand U9827(n9444,n9349,G21779);
  nand U9828(n9443,n7180,n9350);
  nand U9829(n9442,n9351,n7178);
  nand U9830(G1168,n9452,n9453,n9454,n9455);
  nor U9831(n9455,n9456,n9457,n9458);
  nor U9832(n9458,n9459,n9344);
  nor U9833(n9457,n9460,n9346);
  nor U9834(n9456,n9347,n9461);
  nand U9835(n9454,n9349,G21778);
  nand U9836(n9453,n7192,n9350);
  nand U9837(n9452,n9351,n7190);
  nand U9838(G1167,n9462,n9463,n9464,n9465);
  nor U9839(n9465,n9466,n9467,n9468,n9469);
  nor U9840(n9469,n9347,n9470);
  nor U9841(n9468,n9471,n9344);
  nor U9842(n9467,n9472,n9346);
  nand U9843(n9464,n9349,G21777);
  nand U9844(n9463,n7205,n9350);
  nand U9845(n9462,n9351,n7203);
  nand U9846(G1166,n9473,n9474,n9475,n9476);
  nor U9847(n9476,n9466,n9477,n9478,n9479);
  nor U9848(n9479,n9347,n9480);
  nor U9849(n9478,n9481,n9344);
  nor U9850(n9477,n9482,n9346);
  nand U9851(n9475,n9349,G21776);
  nand U9852(n9474,n7217,n9350);
  nand U9853(n9473,n9351,n7215);
  nand U9854(G1165,n9483,n9484,n9485,n9486);
  nor U9855(n9486,n9466,n9487,n9488,n9489);
  nor U9856(n9489,n9347,n9490);
  nor U9857(n9488,n9491,n9344);
  nor U9858(n9487,n9492,n9346);
  nand U9859(n9485,n9349,G21775);
  nand U9860(n9484,n7230,n9350);
  nand U9861(n9483,n9351,n7228);
  nand U9862(G1164,n9493,n9494,n9495,n9496);
  nor U9863(n9496,n9466,n9497,n9498,n9499);
  nor U9864(n9499,n9347,n9500);
  nor U9865(n9498,n9501,n9344);
  nor U9866(n9497,n9502,n9346);
  nand U9867(n9495,n9349,G21774);
  nand U9868(n9494,n7243,n9350);
  nand U9869(n9493,n9351,n7241);
  nand U9870(G1163,n9503,n9504,n9505,n9506);
  nor U9871(n9506,n9466,n9507,n9508,n9509);
  nor U9872(n9509,n9347,n9510);
  nor U9873(n9508,n9511,n9344);
  nor U9874(n9507,n9512,n9346);
  not U9875(n9512,G21741);
  nand U9876(n9505,n9349,G21773);
  nand U9877(n9504,n7260,n9350);
  nand U9878(n9503,n9351,n7258);
  nand U9879(G1162,n9513,n9514,n9515,n9516);
  nor U9880(n9516,n9466,n9517,n9518,n9519);
  nor U9881(n9519,n9347,n9520);
  nor U9882(n9518,n9521,n9344);
  nor U9883(n9517,n9522,n9346);
  not U9884(n9522,G21740);
  nand U9885(n9515,n9349,G21772);
  nand U9886(n9514,n7272,n9350);
  nand U9887(n9513,n9351,n7270);
  nand U9888(G1161,n9523,n9524,n9525,n9526);
  nor U9889(n9526,n9466,n9527,n9528,n9529);
  nor U9890(n9529,n9347,n9530);
  nor U9891(n9528,n9531,n9344);
  nor U9892(n9527,n9532,n9346);
  not U9893(n9532,G21739);
  nand U9894(n9525,n9349,G21771);
  nand U9895(n9524,n7289,n9350);
  nand U9896(n9523,n9351,n7287);
  nand U9897(G1160,n9533,n9534,n9535,n9536);
  nor U9898(n9536,n9466,n9537,n9538,n9539);
  nor U9899(n9539,n9347,n9540);
  nor U9900(n9538,n9541,n9344);
  nor U9901(n9537,n9542,n9346);
  not U9902(n9542,G21738);
  nand U9903(n9535,n9349,G21770);
  nand U9904(n9534,n7301,n9350);
  nand U9905(n9533,n9351,n7299);
  nand U9906(G1159,n9543,n9544,n9545,n9546);
  nor U9907(n9546,n9466,n9547,n9548,n9549);
  nor U9908(n9549,n9347,n9550);
  nor U9909(n9548,n9551,n9344);
  nor U9910(n9547,n9552,n9346);
  not U9911(n9552,G21737);
  nand U9912(n9545,n9349,G21769);
  nand U9913(n9544,n7317,n9350);
  nand U9914(n9543,n9351,n7315);
  nand U9915(G1158,n9553,n9554,n9555,n9556);
  nor U9916(n9556,n9466,n9557,n9558,n9559);
  nor U9917(n9559,n9347,n6916);
  nor U9918(n9558,n6922,n9344);
  not U9919(n6922,G21609);
  nor U9920(n9557,n9560,n9346);
  not U9921(n9560,G21736);
  nand U9922(n9555,n9349,G21768);
  nand U9923(n9554,n9350,n6913);
  nand U9924(n9553,n9351,n9561);
  nand U9925(G1157,n9562,n9563,n9564,n9565);
  nor U9926(n9568,n9347,n7336);
  nor U9927(n9567,n6929,n9344);
  not U9928(n6929,G21608);
  nor U9929(n9566,n9569,n9346);
  not U9930(n9569,G21735);
  nand U9931(n9564,n9349,G21767);
  nand U9932(n9563,n6930,n9350);
  nand U9933(n9562,n9351,n6932);
  nand U9934(G1156,n9570,n9571,n9572,n9573);
  nor U9935(n9576,n9347,n9577);
  nor U9936(n9575,n6941,n9344);
  not U9937(n6941,G21607);
  nor U9938(n9574,n9578,n9346);
  not U9939(n9578,G21734);
  nand U9940(n9572,n9349,G21766);
  nand U9941(n9571,n6944,n9350);
  nand U9942(n9570,n9351,n6945);
  nand U9943(G1155,n9579,n9580,n9581,n9582);
  nor U9944(n9585,n9347,n9586);
  nor U9945(n9584,n6953,n9344);
  not U9946(n6953,G21606);
  nor U9947(n9583,n9587,n9346);
  not U9948(n9587,G21733);
  nand U9949(n9581,n9349,G21765);
  nand U9950(n9580,n6955,n9350);
  nand U9951(n9579,n9351,n6956);
  nand U9952(G1154,n9588,n9589,n9590,n9591);
  nor U9953(n9591,n9466,n9592,n9593,n9594);
  nor U9954(n9594,n9347,n9595);
  nor U9955(n9593,n6964,n9344);
  not U9956(n6964,G21605);
  nor U9957(n9592,n9596,n9346);
  not U9958(n9596,G21732);
  nand U9959(n9590,n9349,G21764);
  nand U9960(n9589,n6966,n9350);
  nand U9961(n9588,n9351,n6967);
  not U9962(n9351,n9597);
  nand U9963(G1153,n9598,n9599,n9600,n9601);
  nor U9964(n9601,n9466,n9602,n9603,n9604);
  nor U9965(n9604,n9605,n9606);
  nor U9966(n9603,n6975,n9344);
  not U9967(n6975,G21604);
  nor U9968(n9602,n9607,n9346);
  not U9969(n9607,G21731);
  nand U9970(n9600,n9349,G21763);
  nand U9971(n9599,n6977,n9350);
  nand U9972(n9598,n6978,n9608);
  nand U9973(G1152,n9609,n9610,n9611,n9612);
  nor U9974(n9612,n9466,n9613,n9614,n9615);
  nor U9975(n9615,n9605,n8873);
  nor U9976(n9614,n6986,n9344);
  nor U9977(n9613,n9616,n9346);
  not U9978(n9616,G21730);
  nor U9979(n9466,G21427,G21428,n9349);
  nand U9980(n9611,n9349,G21762);
  nand U9981(n9610,n6988,n9350);
  nand U9982(n9609,n6989,n9608);
  nand U9983(G1151,n9617,n9618,n9619,n9620);
  nor U9984(n9620,n9621,n9622,n9623);
  nor U9985(n9623,n6997,n9344);
  nor U9986(n9622,n9624,n9346);
  not U9987(n9624,G21729);
  nor U9988(n9621,n9605,n7405);
  nand U9989(n9619,n9349,G21761);
  nand U9990(n9618,n6999,n9350);
  nand U9991(n9617,n7000,n9608);
  nand U9992(G1150,n9625,n9626,n9627,n9628);
  nor U9993(n9628,n9629,n9630,n9631);
  nor U9994(n9631,n7008,n9344);
  nor U9995(n9630,n9632,n9346);
  not U9996(n9632,G21728);
  nor U9997(n9629,n7413,n9605);
  nand U9998(n9627,n9349,G21760);
  nand U9999(n9626,n7009,n9350);
  nand U10000(n9625,n7010,n9608);
  nand U10001(G1149,n9633,n9634,n9635,n9636);
  nor U10002(n9636,n9637,n9638,n9639);
  nor U10003(n9639,n7018,n9344);
  nor U10004(n9638,n9640,n9346);
  not U10005(n9640,G21727);
  nor U10006(n9637,n9605,n9641);
  nand U10007(n9635,n9349,G21759);
  nand U10008(n9634,n7020,n9350);
  nand U10009(n9633,n7021,n9608);
  nand U10010(G1148,n9642,n9643,n9644,n9645);
  nor U10011(n9645,n9646,n9647,n9648);
  nor U10012(n9648,n7029,n9344);
  nor U10013(n9647,n9650,n9346);
  nand U10014(n9652,n9653,n9654);
  nand U10015(n9654,n9655,n9656,n9657);
  or U10016(n9653,n9658,n8921);
  not U10017(n9650,G21726);
  nor U10018(n9646,n9605,n7436);
  and U10019(n9605,n9347,n9659);
  nand U10020(n9659,n8798,n7470,n9651);
  and U10021(n9347,n9660,n9661);
  nand U10022(n9661,n9662,n9657,n9651);
  nand U10023(n9660,G21427,n9649,n7055);
  nand U10024(n9644,n9349,G21758);
  nand U10025(n9643,n7031,n9350);
  nand U10026(n9664,n9651,n9657,n9665,n9656);
  not U10027(n9665,n9655);
  or U10028(n9663,n7055,n9349,n9118);
  nand U10029(n9642,n7032,n9608);
  nand U10030(n9608,n9597,n9666);
  nand U10031(n9666,n9649,n8798,n9667);
  nand U10032(n9597,n8921,n9227,n9651);
  nor U10033(n9651,n7456,n9349);
  nand U10034(n9649,n9083,n7457,n8847,n8831);
  nand U10035(n8831,G21425,G21428,n8824);
  nand U10036(n8847,n7456,n8843,n7590);
  nand U10037(n7457,n9085,n8843,n8824);
  and U10038(n9083,n9668,n9669,n9670);
  or U10039(n9668,n9287,n9117);
  nand U10040(n9287,n9671,n9672,n9673);
  nor U10041(n8921,n9656,n9298);
  not U10042(n9656,n9662);
  nor U10043(n9662,G21797,G35);
  nand U10044(G1147,n9674,n9675);
  nand U10045(n9675,n9676,n7055);
  nand U10046(n9674,G21757,n9677);
  nand U10047(G1146,n9678,n9679,n9680);
  nand U10048(n9680,G21756,n9677);
  nand U10049(n9679,n9676,n9361);
  nand U10050(n9678,n9681,n9682);
  nand U10051(G1145,n9683,n9684,n9685);
  nand U10052(n9685,G21755,n9677);
  nand U10053(n9684,n9676,n9371);
  nand U10054(n9683,n9681,n9686);
  nand U10055(G1144,n9687,n9688,n9689);
  nand U10056(n9689,G21754,n9677);
  nand U10057(n9688,n9676,n9381);
  nand U10058(n9687,n9681,n9690);
  nand U10059(G1143,n9691,n9692,n9693);
  nand U10060(n9693,G21753,n9677);
  nand U10061(n9692,n9676,n9391);
  nand U10062(n9691,n9681,n9694);
  nand U10063(G1142,n9695,n9696,n9697);
  nand U10064(n9697,G21752,n9677);
  nand U10065(n9696,n9676,n9401);
  nand U10066(n9695,n9681,n9698);
  nand U10067(G1141,n9699,n9700,n9701);
  nand U10068(n9701,G21751,n9677);
  nand U10069(n9700,n9676,n7131);
  nand U10070(n9699,n9681,n7130);
  nand U10071(G1140,n9702,n9703,n9704);
  nand U10072(n9704,G21750,n9677);
  nand U10073(n9703,n9676,n9421);
  nand U10074(n9702,n9681,n9705);
  nand U10075(G1139,n9706,n9707,n9708);
  nand U10076(n9708,G21749,n9677);
  nand U10077(n9707,n9676,n7154);
  nand U10078(n9706,n9681,n7153);
  nand U10079(G1138,n9709,n9710,n9711);
  nand U10080(n9711,G21748,n9677);
  nand U10081(n9710,n9676,n7167);
  nand U10082(n9709,n9681,n7166);
  nand U10083(G1137,n9712,n9713,n9714);
  nand U10084(n9714,G21747,n9677);
  nand U10085(n9713,n9676,n7180);
  nand U10086(n9712,n9681,n7179);
  nand U10087(G1136,n9715,n9716,n9717);
  nand U10088(n9717,G21746,n9677);
  nand U10089(n9716,n9676,n7192);
  nand U10090(n9715,n9681,n7191);
  nand U10091(G1135,n9718,n9719,n9720);
  nand U10092(n9720,G21745,n9677);
  nand U10093(n9719,n9676,n7205);
  nand U10094(n9718,n9681,n7204);
  nand U10095(G1134,n9721,n9722,n9723);
  nand U10096(n9723,G21744,n9677);
  nand U10097(n9722,n9676,n7217);
  nand U10098(n9721,n9681,n7216);
  nand U10099(G1133,n9724,n9725,n9726);
  nand U10100(n9726,G21743,n9677);
  nand U10101(n9725,n9676,n7230);
  nand U10102(n9724,n9681,n7229);
  nand U10103(G1132,n9727,n9728,n9729);
  nand U10104(n9729,G21742,n9677);
  nand U10105(n9728,n9676,n7243);
  nand U10106(n9727,n9681,n7242);
  nand U10107(G1131,n9730,n9731,n9732);
  nand U10108(n9732,G21741,n9677);
  nand U10109(n9731,n9676,n7260);
  nand U10110(n9730,n9681,n7259);
  nand U10111(G1130,n9733,n9734,n9735);
  nand U10112(n9735,G21740,n9677);
  nand U10113(n9734,n9676,n7272);
  nand U10114(n9733,n9681,n7271);
  nand U10115(G1129,n9736,n9737,n9738);
  nand U10116(n9738,G21739,n9677);
  nand U10117(n9737,n9676,n7289);
  nand U10118(n9736,n9681,n7288);
  nand U10119(G1128,n9739,n9740,n9741);
  nand U10120(n9741,G21738,n9677);
  nand U10121(n9740,n9676,n7301);
  nand U10122(n9739,n9681,n7300);
  nand U10123(G1127,n9742,n9743,n9744);
  nand U10124(n9744,G21737,n9677);
  nand U10125(n9743,n9676,n7317);
  nand U10126(n9742,n9681,n7316);
  not U10127(n7316,n9550);
  nand U10128(G1126,n9745,n9746,n9747);
  nand U10129(n9747,G21736,n9677);
  nand U10130(n9746,n9676,n6913);
  nand U10131(n9745,n9681,n9748);
  not U10132(n9748,n6916);
  nand U10133(G1125,n9749,n9750,n9751);
  nand U10134(n9751,G21735,n9677);
  nand U10135(n9750,n9676,n6930);
  nand U10136(n9749,n9681,n6934);
  nand U10137(G1124,n9752,n9753,n9754);
  nand U10138(n9754,G21734,n9677);
  nand U10139(n9753,n9676,n6944);
  nand U10140(n9752,n9681,n6946);
  nand U10141(G1123,n9755,n9756,n9757);
  nand U10142(n9757,G21733,n9677);
  nand U10143(n9756,n9676,n6955);
  nand U10144(n9755,n9681,n6957);
  nand U10145(G1122,n9758,n9759,n9760);
  nand U10146(n9760,G21732,n9677);
  nand U10147(n9759,n9676,n6966);
  nand U10148(n9758,n9681,n6968);
  nand U10149(G1121,n9761,n9762,n9763);
  nand U10150(n9763,G21731,n9677);
  nand U10151(n9762,n9676,n6977);
  nand U10152(n9761,n9681,n6979);
  nand U10153(G1120,n9764,n9765,n9766);
  nand U10154(n9766,G21730,n9677);
  nand U10155(n9765,n9676,n6988);
  nand U10156(n9764,n9681,n6990);
  nand U10157(G1119,n9767,n9768,n9769);
  nand U10158(n9769,G21729,n9677);
  nand U10159(n9768,n9676,n6999);
  nand U10160(n9767,n9681,n7001);
  nand U10161(G1118,n9770,n9771,n9772);
  nand U10162(n9772,G21728,n9677);
  nand U10163(n9771,n9676,n7009);
  nand U10164(n9770,n9681,n7011);
  nand U10165(G1117,n9773,n9774,n9775);
  nand U10166(n9775,G21727,n9677);
  nand U10167(n9774,n9676,n7020);
  nand U10168(n9773,n9681,n7022);
  nand U10169(G1116,n9776,n9777,n9778);
  nand U10170(n9778,G21726,n9677);
  nand U10171(n9777,n9676,n7031);
  nand U10172(n9776,n9681,n7033);
  nand U10173(n9780,n9781,n9782);
  nand U10174(n9782,n9783,n7483);
  nand U10175(G1115,n9784,n9785,n9786);
  nand U10176(n9786,G21725,n9787);
  nand U10177(n9785,n9788,G1);
  nand U10178(n9784,n9789,n7055);
  nand U10179(G1114,n9790,n9791,n9792);
  nor U10180(n9792,n9793,n9794,n9795);
  and U10181(n9795,G2,n9788);
  nor U10182(n9794,n9796,n9797);
  not U10183(n9797,G18);
  nor U10184(n9793,n7066,n9798);
  nand U10185(n9791,n9799,n7068);
  nand U10186(n9790,G21724,n9787);
  nand U10187(G1113,n9800,n9801,n9802);
  nor U10188(n9802,n9803,n9804,n9805);
  and U10189(n9805,G3,n9788);
  nor U10190(n9804,n9796,n9806);
  not U10191(n9806,G19);
  nor U10192(n9803,n7080,n9798);
  nand U10193(n9801,n9799,n7081);
  nand U10194(n9800,G21723,n9787);
  nand U10195(G1112,n9807,n9808,n9809);
  nor U10196(n9809,n9810,n9811,n9812);
  and U10197(n9812,G4,n9788);
  nor U10198(n9811,n9796,n9813);
  not U10199(n9813,G20);
  nor U10200(n9810,n7092,n9798);
  nand U10201(n9808,n9799,n7093);
  nand U10202(n9807,G21722,n9787);
  nand U10203(G1111,n9814,n9815,n9816);
  nor U10204(n9816,n9817,n9818,n9819);
  and U10205(n9819,G5,n9788);
  nor U10206(n9818,n9796,n9820);
  not U10207(n9820,G21);
  nor U10208(n9817,n7104,n9798);
  nand U10209(n9815,n9799,n7105);
  nand U10210(n9814,G21721,n9787);
  nand U10211(G1110,n9821,n9822,n9823);
  nor U10212(n9823,n9824,n9825,n9826);
  and U10213(n9826,G6,n9788);
  nor U10214(n9825,n9796,n9827);
  not U10215(n9827,G22);
  nor U10216(n9824,n7116,n9798);
  nand U10217(n9822,n9799,n7117);
  nand U10218(n9821,G21720,n9787);
  nand U10219(G1109,n9828,n9829,n9830);
  nor U10220(n9830,n9831,n9832,n9833);
  and U10221(n9833,G7,n9788);
  nor U10222(n9832,n9796,n9834);
  not U10223(n9834,G23);
  nor U10224(n9831,n9835,n9798);
  nand U10225(n9829,n9799,n7129);
  nand U10226(n9828,G21719,n9787);
  nand U10227(G1108,n9836,n9837,n9838);
  nor U10228(n9838,n9839,n9840,n9841);
  and U10229(n9841,G8,n9788);
  nor U10230(n9840,n9796,n9842);
  not U10231(n9842,G24);
  nor U10232(n9839,n7141,n9798);
  nand U10233(n9837,n9799,n7142);
  nand U10234(n9836,G21718,n9787);
  nand U10235(G1107,n9843,n9844,n9845);
  nor U10236(n9845,n9846,n9847,n9848);
  and U10237(n9848,G9,n9788);
  nor U10238(n9847,n9849,n9796);
  not U10239(n9849,G25);
  nor U10240(n9846,n9850,n9798);
  nand U10241(n9844,n9799,n7152);
  nand U10242(n9843,G21717,n9787);
  nand U10243(G1106,n9851,n9852,n9853);
  nor U10244(n9853,n9854,n9855,n9856);
  and U10245(n9856,G10,n9788);
  nor U10246(n9855,n9857,n9796);
  not U10247(n9857,G26);
  nor U10248(n9854,n9858,n9798);
  nand U10249(n9852,n9799,n7165);
  nand U10250(n9851,G21716,n9787);
  nand U10251(G1105,n9859,n9860,n9861);
  nor U10252(n9861,n9862,n9863,n9864);
  and U10253(n9864,G11,n9788);
  nor U10254(n9863,n9865,n9796);
  not U10255(n9865,G27);
  nor U10256(n9862,n9866,n9798);
  nand U10257(n9860,n9799,n7178);
  nand U10258(n9859,G21715,n9787);
  nand U10259(G1104,n9867,n9868,n9869);
  nor U10260(n9869,n9870,n9871,n9872);
  and U10261(n9872,G12,n9788);
  nor U10262(n9871,n9873,n9796);
  not U10263(n9873,G28);
  nor U10264(n9870,n9874,n9798);
  nand U10265(n9868,n9799,n7190);
  nand U10266(n9867,G21714,n9787);
  nand U10267(G1103,n9875,n9876,n9877);
  nor U10268(n9877,n9878,n9879,n9880);
  and U10269(n9880,G13,n9788);
  nor U10270(n9879,n9881,n9796);
  not U10271(n9881,G29);
  nor U10272(n9878,n9882,n9798);
  nand U10273(n9876,n9799,n7203);
  nand U10274(n9875,G21713,n9787);
  nand U10275(G1102,n9883,n9884,n9885);
  nor U10276(n9885,n9886,n9887,n9888);
  and U10277(n9888,G14,n9788);
  nor U10278(n9887,n9889,n9796);
  not U10279(n9889,G30);
  nor U10280(n9886,n9890,n9798);
  nand U10281(n9884,n9799,n7215);
  nand U10282(n9883,G21712,n9787);
  nand U10283(G1101,n9891,n9892,n9893);
  nor U10284(n9893,n9894,n9895,n9896);
  and U10285(n9896,G15,n9788);
  nor U10286(n9895,n9897,n9796);
  not U10287(n9897,G31);
  nor U10288(n9894,n9898,n9798);
  nand U10289(n9892,n9799,n7228);
  nand U10290(n9891,G21711,n9787);
  nand U10291(G1100,n9899,n9900,n9901);
  nor U10292(n9901,n9902,n9903,n9904);
  and U10293(n9904,G16,n9788);
  nor U10294(n9788,n9787,n7465);
  nor U10295(n9903,n9905,n9796);
  or U10296(n9796,n9787,n9101);
  not U10297(n9905,G32);
  nor U10298(n9902,n9906,n9798);
  not U10299(n9798,n9789);
  nand U10300(n9900,n9799,n7241);
  nand U10301(n9899,G21710,n9787);
  nand U10302(G1099,n9907,n9908,n9909,n9910);
  nand U10303(n9910,n9789,n7260);
  nand U10304(n9909,n9799,n7258);
  nand U10305(n9908,G17,n9911);
  nand U10306(n9907,G21709,n9787);
  nand U10307(G1098,n9912,n9913,n9914,n9915);
  nand U10308(n9915,n9789,n7272);
  nand U10309(n9914,n9799,n7270);
  nand U10310(n9913,n9911,G18);
  nand U10311(n9912,G21708,n9787);
  nand U10312(G1097,n9916,n9917,n9918,n9919);
  nand U10313(n9919,n9789,n7289);
  nand U10314(n9918,n9799,n7287);
  nand U10315(n9917,n9911,G19);
  nand U10316(n9916,G21707,n9787);
  nand U10317(G1096,n9920,n9921,n9922,n9923);
  nand U10318(n9923,n9789,n7301);
  nand U10319(n9922,n9799,n7299);
  nand U10320(n9921,n9911,G20);
  nand U10321(n9920,G21706,n9787);
  nand U10322(G1095,n9924,n9925,n9926,n9927);
  nand U10323(n9927,n9789,n7317);
  nand U10324(n9926,n9799,n7315);
  nand U10325(n9925,n9911,G21);
  nand U10326(n9924,G21705,n9787);
  nand U10327(G1094,n9928,n9929,n9930,n9931);
  nand U10328(n9931,n9799,n9561);
  not U10329(n9561,n6918);
  nand U10330(n6918,n9932,n9933,n9934);
  nand U10331(n9934,n9935,n9936);
  nand U10332(n9935,n9937,n9938);
  or U10333(n9938,n9939,n9940);
  nand U10334(n9933,n9941,n9939);
  or U10335(n9932,n9937,n9939);
  nand U10336(n9930,n9789,n6913);
  nand U10337(n9929,n9911,G22);
  nand U10338(n9928,G21704,n9787);
  nand U10339(G1093,n9942,n9943,n9944,n9945);
  nand U10340(n9945,n9799,n6932);
  nand U10341(n6932,n9946,n9947,n9948);
  not U10342(n9948,n9941);
  nor U10343(n9941,n9949,n9936,n9950);
  nand U10344(n9947,n9951,n9936);
  or U10345(n9951,n9952,n9949);
  nand U10346(n9946,n9940,n9953);
  nand U10347(n9944,n9789,n6930);
  nand U10348(n9943,n9911,G23);
  nand U10349(n9942,G21703,n9787);
  nand U10350(G1092,n9954,n9955,n9956,n9957);
  nand U10351(n9957,n9799,n6945);
  or U10352(n6945,n9958,n9959);
  or U10353(n9959,n9953,n9960);
  nand U10354(n9956,n9789,n6944);
  nand U10355(n9955,n9911,G24);
  nand U10356(n9954,G21702,n9787);
  nand U10357(G1091,n9961,n9962,n9963,n9964);
  nand U10358(n9964,n9799,n6956);
  or U10359(n6956,n9965,n9966);
  and U10360(n9966,n9967,n9968);
  nand U10361(n9963,n9789,n6955);
  nand U10362(n9962,n9911,G25);
  nand U10363(n9961,G21701,n9787);
  nand U10364(G1090,n9969,n9970,n9971,n9972);
  nand U10365(n9972,n9799,n6967);
  and U10366(n6967,n9973,n9974);
  nand U10367(n9974,n9975,n9976);
  not U10368(n9975,n9977);
  nand U10369(n9973,n9978,n9979,n9980);
  nand U10370(n9978,n9976,n9981);
  nand U10371(n9971,n9789,n6966);
  nand U10372(n9970,n9911,G26);
  nand U10373(n9969,G21700,n9787);
  nand U10374(G1089,n9982,n9983,n9984,n9985);
  nand U10375(n9985,n9799,n6978);
  or U10376(n6978,n9986,n9987);
  and U10377(n9987,n9979,n9988);
  nand U10378(n9984,n9789,n6977);
  nand U10379(n9983,n9911,G27);
  nand U10380(n9982,G21699,n9787);
  nand U10381(G1088,n9989,n9990,n9991,n9992);
  nand U10382(n9992,n9799,n6989);
  or U10383(n6989,n9993,n9994);
  and U10384(n9994,n9995,n9996);
  nand U10385(n9991,n9789,n6988);
  nand U10386(n9990,n9911,G28);
  nand U10387(n9989,G21698,n9787);
  nand U10388(G1087,n9997,n9998,n9999,n10000);
  nand U10389(n10000,n9799,n7000);
  and U10390(n7000,n10001,n10002);
  nand U10391(n10002,n10003,n10004);
  nand U10392(n10004,n10005,n10006);
  not U10393(n10003,n10007);
  nand U10394(n10001,n10005,n10006,n10007);
  nand U10395(n9999,n9789,n6999);
  nand U10396(n9998,n9911,G29);
  nand U10397(n9997,G21697,n9787);
  nand U10398(G1086,n10008,n10009,n10010,n10011);
  nand U10399(n10011,n9799,n7010);
  and U10400(n7010,n10012,n10013);
  nand U10401(n10013,n10014,n10015,n10016);
  nand U10402(n10014,n10017,n10018);
  nand U10403(n10012,n10019,n10017);
  not U10404(n10019,n10020);
  nand U10405(n10010,n9789,n7009);
  nand U10406(n10009,n9911,G30);
  nand U10407(n10008,G21696,n9787);
  nand U10408(G1085,n10021,n10022,n10023,n10024);
  nand U10409(n10024,n9799,n7021);
  or U10410(n7021,n10025,n10026);
  and U10411(n10026,n10015,n10027);
  nand U10412(n10023,n9789,n7020);
  nand U10413(n10022,n9911,G31);
  nand U10414(n10021,G21695,n9787);
  nand U10415(G1084,n10028,n10029,n10030,n10031);
  nand U10416(n10031,n9789,n7031);
  nor U10417(n9789,n9787,n9307);
  nand U10418(n10030,n9799,n7032);
  or U10419(n7032,n10032,n9953);
  nand U10420(n10032,n10033,n10034);
  nand U10421(n10029,n9911,G32);
  nor U10422(n9911,n9787,n9248);
  nand U10423(n10028,G21694,n9787);
  nand U10424(n10038,n7467,n7471,n9284);
  not U10425(n7471,G35);
  nand U10426(n10037,n10040,n7473);
  nor U10427(n7473,n9117,G35);
  nand U10428(n10036,n10041,n7483);
  and U10429(G1083,G21693,n10042);
  nand U10430(G1082,n10043,n10044,n10045);
  nand U10431(n10045,G21692,n10042);
  nand U10432(n10044,n10046,G21724);
  nand U10433(n10043,G21647,n10047);
  nand U10434(G1081,n10048,n10049,n10050);
  nand U10435(n10050,G21691,n10042);
  nand U10436(n10049,n10046,G21723);
  nand U10437(n10048,G21648,n10047);
  nand U10438(G1080,n10051,n10052,n10053);
  nand U10439(n10053,G21690,n10042);
  nand U10440(n10052,n10046,G21722);
  nand U10441(n10051,G21649,n10047);
  nand U10442(G1079,n10054,n10055,n10056);
  nand U10443(n10056,G21689,n10042);
  nand U10444(n10055,n10046,G21721);
  nand U10445(n10054,G21650,n10047);
  nand U10446(G1078,n10057,n10058,n10059);
  nand U10447(n10059,G21688,n10042);
  nand U10448(n10058,n10046,G21720);
  nand U10449(n10057,G21651,n10047);
  nand U10450(G1077,n10060,n10061,n10062);
  nand U10451(n10062,G21687,n10042);
  nand U10452(n10061,n10046,G21719);
  nand U10453(n10060,G21652,n10047);
  nand U10454(G1076,n10063,n10064,n10065);
  nand U10455(n10065,G21686,n10042);
  nand U10456(n10064,n10046,G21718);
  nand U10457(n10063,G21653,n10047);
  nand U10458(G1075,n10066,n10067,n10068);
  nand U10459(n10068,G21685,n10042);
  nand U10460(n10067,n10046,G21717);
  nand U10461(n10066,G21654,n10047);
  nand U10462(G1074,n10069,n10070,n10071);
  nand U10463(n10071,G21684,n10042);
  nand U10464(n10070,n10046,G21716);
  nand U10465(n10069,G21655,n10047);
  nand U10466(G1073,n10072,n10073,n10074);
  nand U10467(n10074,G21683,n10042);
  nand U10468(n10073,n10046,G21715);
  nand U10469(n10072,G21656,n10047);
  nand U10470(G1072,n10075,n10076,n10077);
  nand U10471(n10077,G21682,n10042);
  nand U10472(n10076,n10046,G21714);
  nand U10473(n10075,G21657,n10047);
  nand U10474(G1071,n10078,n10079,n10080);
  nand U10475(n10080,G21681,n10042);
  nand U10476(n10079,n10046,G21713);
  nand U10477(n10078,G21658,n10047);
  nand U10478(G1070,n10081,n10082,n10083);
  nand U10479(n10083,G21680,n10042);
  nand U10480(n10082,n10046,G21712);
  nand U10481(n10081,G21659,n10047);
  nand U10482(G1069,n10084,n10085,n10086);
  nand U10483(n10086,G21679,n10042);
  nand U10484(n10085,n10046,G21711);
  nand U10485(n10084,G21660,n10047);
  nand U10486(G1068,n10087,n10088,n10089);
  nand U10487(n10089,G21678,n10042);
  nand U10488(n10088,n10046,G21710);
  and U10489(n10046,n10090,n8737);
  nand U10490(n10087,G21661,n10047);
  nand U10491(G1067,n10091,n10092,n10093);
  nand U10492(n10093,G21677,n10042);
  nand U10493(n10092,n10090,G21709);
  nand U10494(n10091,G21631,n10047);
  nand U10495(G1066,n10094,n10095,n10096);
  nand U10496(n10096,G21676,n10042);
  nand U10497(n10095,n10090,G21708);
  nand U10498(n10094,G21632,n10047);
  nand U10499(G1065,n10097,n10098,n10099);
  nand U10500(n10099,G21675,n10042);
  nand U10501(n10098,n10090,G21707);
  nand U10502(n10097,G21633,n10047);
  nand U10503(G1064,n10100,n10101,n10102);
  nand U10504(n10102,G21674,n10042);
  nand U10505(n10101,n10090,G21706);
  nand U10506(n10100,G21634,n10047);
  nand U10507(G1063,n10103,n10104,n10105);
  nand U10508(n10105,G21673,n10042);
  nand U10509(n10104,n10090,G21705);
  nand U10510(n10103,G21635,n10047);
  nand U10511(G1062,n10106,n10107,n10108);
  nand U10512(n10108,G21672,n10042);
  nand U10513(n10107,n10090,G21704);
  nand U10514(n10106,G21636,n10047);
  nand U10515(G1061,n10109,n10110,n10111);
  nand U10516(n10111,G21671,n10042);
  nand U10517(n10110,n10090,G21703);
  nand U10518(n10109,G21637,n10047);
  nand U10519(G1060,n10112,n10113,n10114);
  nand U10520(n10114,G21670,n10042);
  nand U10521(n10113,n10090,G21702);
  nand U10522(n10112,G21638,n10047);
  nand U10523(G1059,n10115,n10116,n10117);
  nand U10524(n10117,G21669,n10042);
  nand U10525(n10116,n10090,G21701);
  nand U10526(n10115,G21639,n10047);
  nand U10527(G1058,n10118,n10119,n10120);
  nand U10528(n10120,G21668,n10042);
  nand U10529(n10119,n10090,G21700);
  nand U10530(n10118,G21640,n10047);
  nand U10531(G1057,n10121,n10122,n10123);
  nand U10532(n10123,G21667,n10042);
  nand U10533(n10122,n10090,G21699);
  nand U10534(n10121,G21641,n10047);
  nand U10535(G1056,n10124,n10125,n10126);
  nand U10536(n10126,G21666,n10042);
  nand U10537(n10125,n10090,G21698);
  nand U10538(n10124,G21642,n10047);
  nand U10539(G1055,n10127,n10128,n10129);
  nand U10540(n10129,G21665,n10042);
  nand U10541(n10128,n10090,G21697);
  nand U10542(n10127,G21643,n10047);
  nand U10543(G1054,n10130,n10131,n10132);
  nand U10544(n10132,G21664,n10042);
  nand U10545(n10131,n10090,G21696);
  nand U10546(n10130,G21644,n10047);
  nand U10547(G1053,n10133,n10134,n10135);
  nand U10548(n10135,G21663,n10042);
  nand U10549(n10134,n10090,G21695);
  nand U10550(n10133,G21645,n10047);
  nand U10551(G1052,n10136,n10137,n10138);
  nand U10552(n10138,G21662,n10042);
  nand U10553(n10137,n10090,G21694);
  nor U10554(n10090,n8843,n10042);
  nand U10555(n10136,G21646,n10047);
  nand U10556(n10140,n7480,n10141);
  nand U10557(n10141,n9669,n10142);
  nand U10558(n10142,n9200,n7483,n7459);
  not U10559(n7480,n9298);
  nand U10560(n9298,n8984,n10143);
  not U10561(n8984,G21392);
  nand U10562(n10139,n9096,G21427);
  nand U10563(G1051,n10144,n10145,n10146);
  nand U10564(n10146,n10147,G21661);
  nand U10565(n10144,n10148,G21710);
  nand U10566(G1050,n10149,n10150,n10151);
  nand U10567(n10151,n10147,G21660);
  nand U10568(n10149,n10148,G21711);
  nand U10569(G1049,n10152,n10153,n10154);
  nand U10570(n10154,n10147,G21659);
  nand U10571(n10152,n10148,G21712);
  nand U10572(G1048,n10155,n10156,n10157);
  nand U10573(n10157,n10147,G21658);
  nand U10574(n10155,n10148,G21713);
  nand U10575(G1047,n10158,n10159,n10160);
  nand U10576(n10160,n10147,G21657);
  nand U10577(n10158,n10148,G21714);
  nand U10578(G1046,n10161,n10162,n10163);
  nand U10579(n10163,n10147,G21656);
  nand U10580(n10161,n10148,G21715);
  nand U10581(G1045,n10164,n10165,n10166);
  nand U10582(n10166,n10147,G21655);
  nand U10583(n10164,n10148,G21716);
  nand U10584(G1044,n10167,n10168,n10169);
  nand U10585(n10169,n10147,G21654);
  nand U10586(n10167,n10148,G21717);
  nand U10587(G1043,n10170,n10171,n10172);
  nand U10588(n10172,n10147,G21653);
  nand U10589(n10170,n10148,G21718);
  nand U10590(G1042,n10173,n10174,n10175);
  nand U10591(n10175,n10147,G21652);
  nand U10592(n10173,n10148,G21719);
  nand U10593(G1041,n10176,n10177,n10178);
  nand U10594(n10178,n10147,G21651);
  nand U10595(n10176,n10148,G21720);
  nand U10596(G1040,n10179,n10180,n10181);
  nand U10597(n10181,n10147,G21650);
  nand U10598(n10179,n10148,G21721);
  nand U10599(G1039,n10182,n10183,n10184);
  nand U10600(n10184,n10147,G21649);
  nand U10601(n10182,n10148,G21722);
  nand U10602(G1038,n10185,n10186,n10187);
  nand U10603(n10187,n10147,G21648);
  nand U10604(n10185,n10148,G21723);
  nand U10605(G1037,n10188,n10189,n10190);
  nand U10606(n10190,n10147,G21647);
  nand U10607(n10188,n10148,G21724);
  nand U10608(G1036,n10191,n10145,n10192);
  nand U10609(n10192,n10147,G21646);
  nand U10610(n10145,n10193,G32);
  nand U10611(n10191,n10148,G21694);
  nand U10612(G1035,n10194,n10150,n10195);
  nand U10613(n10195,n10147,G21645);
  nand U10614(n10150,n10193,G31);
  nand U10615(n10194,n10148,G21695);
  nand U10616(G1034,n10196,n10153,n10197);
  nand U10617(n10197,n10147,G21644);
  nand U10618(n10153,n10193,G30);
  nand U10619(n10196,n10148,G21696);
  nand U10620(G1033,n10198,n10156,n10199);
  nand U10621(n10199,n10147,G21643);
  nand U10622(n10156,n10193,G29);
  nand U10623(n10198,n10148,G21697);
  nand U10624(G1032,n10200,n10159,n10201);
  nand U10625(n10201,n10147,G21642);
  nand U10626(n10159,n10193,G28);
  nand U10627(n10200,n10148,G21698);
  nand U10628(G1031,n10202,n10162,n10203);
  nand U10629(n10203,n10147,G21641);
  nand U10630(n10162,n10193,G27);
  nand U10631(n10202,n10148,G21699);
  nand U10632(G1030,n10204,n10165,n10205);
  nand U10633(n10205,n10147,G21640);
  nand U10634(n10165,n10193,G26);
  nand U10635(n10204,n10148,G21700);
  nand U10636(G1029,n10206,n10168,n10207);
  nand U10637(n10207,n10147,G21639);
  nand U10638(n10168,n10193,G25);
  nand U10639(n10206,n10148,G21701);
  nand U10640(G1028,n10208,n10171,n10209);
  nand U10641(n10209,n10147,G21638);
  nand U10642(n10171,n10193,G24);
  nand U10643(n10208,n10148,G21702);
  nand U10644(G1027,n10210,n10174,n10211);
  nand U10645(n10211,n10147,G21637);
  nand U10646(n10174,n10193,G23);
  nand U10647(n10210,n10148,G21703);
  nand U10648(G1026,n10212,n10177,n10213);
  nand U10649(n10213,n10147,G21636);
  nand U10650(n10177,n10193,G22);
  nand U10651(n10212,n10148,G21704);
  nand U10652(G1025,n10214,n10180,n10215);
  nand U10653(n10215,n10147,G21635);
  nand U10654(n10180,n10193,G21);
  nand U10655(n10214,n10148,G21705);
  nand U10656(G1024,n10216,n10183,n10217);
  nand U10657(n10217,n10147,G21634);
  nand U10658(n10183,n10193,G20);
  nand U10659(n10216,n10148,G21706);
  nand U10660(G1023,n10218,n10186,n10219);
  nand U10661(n10219,n10147,G21633);
  nand U10662(n10186,n10193,G19);
  nand U10663(n10218,n10148,G21707);
  nand U10664(G1022,n10220,n10189,n10221);
  nand U10665(n10221,n10147,G21632);
  nand U10666(n10189,n10193,G18);
  nand U10667(n10220,n10148,G21708);
  nand U10668(G1021,n10222,n10223,n10224);
  nand U10669(n10224,n10147,G21631);
  nand U10670(n10223,n10193,G17);
  nor U10671(n10193,n7477,n10147);
  nand U10672(n10222,n10148,G21709);
  nand U10673(n9669,n8882,n7483,n7459);
  nor U10674(n7459,n8854,n8843);
  not U10675(n8854,n8844);
  or U10676(n10225,n9670,G35);
  nand U10677(n9670,n9284,n7467,n8844);
  nor U10678(n8844,n7456,G21427);
  nand U10679(G1020,n10226,n10227,n10228,n10229);
  nor U10680(n10229,n10230,n10231);
  nor U10681(n10231,n6921,n9343);
  nor U10682(n10230,n6943,n7048);
  nand U10683(n10228,n6933,n7053);
  nand U10684(n10227,n7051,n6931);
  or U10685(n7051,n10232,n10233);
  or U10686(n10233,n9953,n10234);
  nand U10687(n10234,n10235,n10236,n10237,n10238);
  nand U10688(n10238,n7055,n9953);
  nand U10689(n10237,n7053,n10239);
  or U10690(n7053,n10240,n10241);
  nor U10691(n10241,n10242,n7590);
  nor U10692(n10242,n10243,n10244,n10245);
  nor U10693(n10245,n10246,n9343);
  and U10694(n10244,n10247,G21598);
  nor U10695(n10243,n10248,n7048);
  not U10696(n7048,G21789);
  nand U10697(n10236,G21789,n10249);
  nand U10698(n10235,G21598,n10250);
  nand U10699(n10232,n10251,n10252);
  nand U10700(n10252,n10253,n9936);
  nand U10701(n10253,n10254,n10255);
  or U10702(n10251,n10254,n10255);
  nand U10703(n10226,n7055,n6912);
  or U10704(n7055,n10256,n10257);
  nor U10705(n10257,n10258,n10259,n10260,n10261);
  nor U10706(n10261,n9110,n9343);
  not U10707(n9343,G21630);
  nor U10708(n10260,n10262,n7044);
  nor U10709(n10259,n10263,n9345);
  and U10710(n10258,n10264,G21725);
  or U10711(n10256,n10265,n10248);
  nand U10712(G1019,n10266,n10267,n10268,n10269);
  nor U10713(n10269,n10270,n10271);
  nor U10714(n10271,n6921,n9359);
  nor U10715(n10270,n6943,n10272);
  nand U10716(n10268,n9361,n6912);
  nand U10717(n10267,n6931,n7068);
  or U10718(n7068,n10255,n10273);
  or U10719(n10273,n9953,n10254);
  nand U10720(n10254,n10274,n10275);
  nand U10721(n10275,n9953,n10276);
  or U10722(n10276,n10277,n10278);
  nand U10723(n10274,n10278,n10277);
  nand U10724(n10255,n10279,n10280,n10281,n10282);
  nor U10725(n10282,n10283,n10284);
  nor U10726(n10284,n10285,n10286);
  nor U10727(n10283,n10287,n10272);
  nand U10728(n10281,n9361,n9953);
  nand U10729(n10289,n9682,n10291);
  nand U10730(n10288,n10292,n7064);
  nand U10731(n10292,n10293,n10291);
  nor U10732(n10291,n7089,n7077);
  nand U10733(n10279,n9682,n10294);
  nand U10734(n10266,n9682,n6933);
  not U10735(n9682,n7064);
  nand U10736(n7064,n10240,n10295);
  nand U10737(n10295,n10296,n10297);
  or U10738(n10240,n10297,n10296);
  or U10739(n10296,n10298,n9110);
  nand U10740(n10298,n10299,n10300,n10301,n10302);
  nor U10741(n10302,n10303,n10304);
  nor U10742(n10304,n10248,n10272);
  not U10743(n10272,G21788);
  nor U10744(n10303,n10246,n9359);
  nand U10745(n10301,G21597,n10247);
  nand U10746(n10300,n9361,n10305);
  not U10747(n9361,n7066);
  nand U10748(n7066,n10265,n10306);
  nand U10749(n10306,n10307,n10308);
  or U10750(n10265,n10308,n10307);
  or U10751(n10307,n10309,n10248);
  nand U10752(n10309,n10310,n10311,n10312,n10313);
  nor U10753(n10313,n10314,n10315);
  nor U10754(n10315,n9110,n9359);
  not U10755(n9359,G21629);
  nor U10756(n10314,n10262,n10286);
  nand U10757(n10312,G21756,n10316);
  nand U10758(n10311,n7065,n7042,n9783);
  nand U10759(n7042,n10317,n10318,n7078);
  nand U10760(n10318,n9101,n10286);
  not U10761(n10286,G21597);
  or U10762(n10317,n10319,n9101);
  nand U10763(n7065,n10320,n10321,n10322);
  nand U10764(n10321,G21597,n9101);
  nand U10765(n10320,n10319,n8737);
  nand U10766(n10319,n10323,n10324,n10325,n10326);
  nor U10767(n10326,n10327,n10328,n10329,n10330);
  nor U10768(n10330,n10331,n10332);
  nor U10769(n10329,n10333,n10334);
  nor U10770(n10328,n10335,n10336);
  nor U10771(n10327,n10337,n10338);
  nor U10772(n10325,n10339,n10340,n10341,n10342);
  nor U10773(n10342,n10343,n10344);
  nor U10774(n10341,n10345,n10346);
  nor U10775(n10340,n10347,n10348);
  nor U10776(n10339,n10349,n10350);
  nor U10777(n10324,n10351,n10352,n10353,n10354);
  nor U10778(n10354,n10355,n10356);
  nor U10779(n10353,n10357,n10358);
  nor U10780(n10352,n10359,n10360);
  nor U10781(n10351,n10361,n10362);
  nor U10782(n10323,n10363,n10364,n10365,n10366);
  nor U10783(n10366,n10367,n10368);
  nor U10784(n10365,n10369,n10370);
  nor U10785(n10364,n10371,n10372);
  nor U10786(n10363,n10373,n10374);
  nand U10787(n10310,G21724,n10264);
  nand U10788(n10299,n10041,n10375);
  or U10789(n10297,n10376,n10377);
  nand U10790(G1018,n10378,n10379,n10380,n10381);
  nor U10791(n10381,n10382,n10383);
  nor U10792(n10383,n6921,n9369);
  nor U10793(n10382,n6943,n10384);
  nand U10794(n10380,n9371,n6912);
  nand U10795(n10379,n6931,n7081);
  or U10796(n7081,n10278,n10385);
  or U10797(n10385,n9953,n10277);
  nand U10798(n10277,n10386,n10387);
  nand U10799(n10387,n9953,n10388);
  or U10800(n10388,n10389,n10390);
  nand U10801(n10386,n10390,n10389);
  nand U10802(n10278,n10391,n10392,n10393,n10394);
  nor U10803(n10394,n10395,n10396);
  nor U10804(n10396,n10285,n10397);
  nor U10805(n10395,n10287,n10384);
  nand U10806(n10393,n9371,n9953);
  nand U10807(n10399,n9690,n10400);
  nand U10808(n10400,n10293,n7077);
  nand U10809(n10398,n7077,n7089);
  nand U10810(n10391,n9686,n10294);
  nand U10811(n10378,n9686,n6933);
  not U10812(n9686,n7077);
  or U10813(n7077,n10376,n10377);
  or U10814(n10377,n10401,n9110);
  nand U10815(n10401,n10402,n10403,n10404,n10405);
  nor U10816(n10405,n10406,n10407);
  nor U10817(n10407,n10248,n10384);
  not U10818(n10384,G21787);
  nor U10819(n10406,n10246,n9369);
  nand U10820(n10404,G21596,n10247);
  nand U10821(n10403,n9371,n10305);
  not U10822(n9371,n7080);
  nand U10823(n7080,n10308,n10408);
  nand U10824(n10408,n10409,n10410);
  or U10825(n10308,n10410,n10409);
  or U10826(n10409,n10411,n10248);
  nand U10827(n10411,n10412,n10413,n10414,n10415);
  nor U10828(n10415,n10416,n10417);
  nor U10829(n10417,n9110,n9369);
  not U10830(n9369,G21628);
  nor U10831(n10416,n10262,n10397);
  not U10832(n10397,G21596);
  nand U10833(n10414,G21755,n10316);
  or U10834(n10413,n7079,n7078,n9290);
  not U10835(n7078,n10322);
  nand U10836(n10322,n10418,n10419);
  nor U10837(n7079,n10419,n10418);
  not U10838(n10418,n7090);
  nand U10839(n10419,n10420,n10421);
  nand U10840(n10421,G21596,n9101);
  nand U10841(n10420,n10422,n8737);
  nand U10842(n10422,n10423,n10424,n10425,n10426);
  nor U10843(n10426,n10427,n10428,n10429,n10430);
  nor U10844(n10430,n10431,n10332);
  nor U10845(n10429,n10432,n10334);
  nor U10846(n10428,n10433,n10336);
  nor U10847(n10427,n10434,n10338);
  nor U10848(n10425,n10435,n10436,n10437,n10438);
  nor U10849(n10438,n10439,n10344);
  nor U10850(n10437,n10440,n10346);
  nor U10851(n10436,n10441,n10348);
  nor U10852(n10435,n10442,n10350);
  nor U10853(n10424,n10443,n10444,n10445,n10446);
  nor U10854(n10446,n10447,n10356);
  nor U10855(n10445,n10448,n10358);
  nor U10856(n10444,n10449,n10360);
  nor U10857(n10443,n10450,n10362);
  nor U10858(n10423,n10451,n10452,n10453,n10454);
  nor U10859(n10454,n10455,n10368);
  nor U10860(n10453,n10456,n10370);
  nor U10861(n10452,n10457,n10372);
  nor U10862(n10451,n10458,n10374);
  nand U10863(n10412,G21723,n10264);
  nand U10864(n10402,n10041,n10459);
  nand U10865(G1017,n10460,n10461,n10462,n10463);
  nor U10866(n10463,n10464,n10465);
  nor U10867(n10465,n6921,n9379);
  nor U10868(n10464,n6943,n10466);
  nand U10869(n10462,n9381,n6912);
  nand U10870(n10461,n6931,n7093);
  or U10871(n7093,n10390,n10467);
  or U10872(n10467,n9953,n10389);
  nand U10873(n10389,n10468,n10469);
  nand U10874(n10469,n9953,n10470);
  or U10875(n10470,n10471,n10472);
  nand U10876(n10468,n10472,n10471);
  nand U10877(n10390,n10473,n10474,n10475,n10476);
  nor U10878(n10476,n10477,n10478);
  nor U10879(n10478,n10287,n10466);
  nor U10880(n10477,n9936,n7092);
  nand U10881(n10475,G21595,n10250);
  nand U10882(n10474,n9690,n10294);
  nand U10883(n10473,n10293,n10290,n7089);
  nand U10884(n10460,n9690,n6933);
  not U10885(n9690,n7089);
  nand U10886(n7089,n10479,n10376);
  nand U10887(n10376,n10480,n10481,n10482);
  not U10888(n10480,n10483);
  nand U10889(n10479,n10483,n10484);
  nand U10890(n10484,n10482,n10481);
  or U10891(n10483,n10485,n9110);
  nand U10892(n10485,n10486,n10487,n10488);
  nor U10893(n10488,n10489,n10490,n10491);
  nor U10894(n10491,n10248,n10466);
  not U10895(n10466,G21786);
  nor U10896(n10490,n10246,n9379);
  and U10897(n10489,n10492,n10041);
  nand U10898(n10487,G21595,n10247);
  nand U10899(n10486,n9381,n10305);
  not U10900(n9381,n7092);
  nand U10901(n7092,n10410,n10493);
  nand U10902(n10493,n10494,n10495);
  or U10903(n10410,n10495,n10494);
  or U10904(n10494,n10496,n10248);
  nand U10905(n10496,n10497,n10498,n10499,n10500);
  nor U10906(n10500,n10501,n10502);
  nor U10907(n10502,n9110,n9379);
  not U10908(n9379,G21627);
  nor U10909(n10501,n10262,n10503);
  not U10910(n10262,n10504);
  nand U10911(n10499,G21754,n10316);
  nand U10912(n10498,n7091,n7090,n9783);
  nand U10913(n7090,n10505,n10506,n7102);
  nand U10914(n10506,n9101,n10503);
  not U10915(n10503,G21595);
  or U10916(n10505,n10507,n9101);
  nand U10917(n7091,n10508,n10509,n10510);
  nand U10918(n10509,G21595,n9101);
  nand U10919(n10508,n10507,n8737);
  nand U10920(n10507,n10511,n10512,n10513,n10514);
  nor U10921(n10514,n10515,n10516,n10517,n10518);
  nor U10922(n10518,n10519,n10332);
  nor U10923(n10517,n10520,n10334);
  nor U10924(n10516,n10521,n10336);
  nor U10925(n10515,n10522,n10338);
  nor U10926(n10513,n10523,n10524,n10525,n10526);
  nor U10927(n10526,n10527,n10344);
  nor U10928(n10525,n10528,n10346);
  nor U10929(n10524,n10529,n10348);
  nor U10930(n10523,n10530,n10350);
  nor U10931(n10512,n10531,n10532,n10533,n10534);
  nor U10932(n10534,n10535,n10356);
  nor U10933(n10533,n10536,n10358);
  nor U10934(n10532,n10537,n10360);
  nor U10935(n10531,n10538,n10362);
  nor U10936(n10511,n10539,n10540,n10541,n10542);
  nor U10937(n10542,n10543,n10368);
  nor U10938(n10541,n10544,n10370);
  nor U10939(n10540,n10545,n10372);
  nor U10940(n10539,n10546,n10374);
  nand U10941(n10497,G21722,n10264);
  nand U10942(G1016,n10547,n10548,n10549,n10550);
  nor U10943(n10550,n10551,n10552);
  nor U10944(n10552,n6921,n9389);
  nor U10945(n10551,n6943,n10553);
  nand U10946(n10549,n9391,n6912);
  nand U10947(n10548,n6931,n7105);
  or U10948(n7105,n10472,n10554);
  or U10949(n10554,n9953,n10471);
  nand U10950(n10471,n10555,n10556);
  nand U10951(n10556,n9953,n10557);
  or U10952(n10557,n10558,n10559);
  nand U10953(n10555,n10559,n10558);
  nand U10954(n10472,n10560,n10561,n10562,n10563);
  nor U10955(n10563,n10564,n10565);
  nor U10956(n10565,n10285,n10566);
  nor U10957(n10564,n10287,n10553);
  nand U10958(n10562,n9391,n9953);
  nand U10959(n10561,n10567,n9698,n10290,n10568);
  nand U10960(n10560,n9694,n10294);
  nand U10961(n10294,n10569,n10570);
  not U10962(n10568,n10293);
  nor U10963(n10293,n7101,n7113,n10571);
  not U10964(n7101,n9694);
  nand U10965(n10547,n9694,n6933);
  or U10966(n9694,n10482,n10481);
  or U10967(n10481,n10572,n9110);
  nand U10968(n10572,n10573,n10574,n10575,n10576);
  nor U10969(n10576,n10577,n10578);
  nor U10970(n10578,n10248,n10553);
  not U10971(n10553,G21785);
  nor U10972(n10577,n10246,n9389);
  not U10973(n9389,G21626);
  nand U10974(n10575,G21594,n10247);
  nand U10975(n10574,n9391,n10305);
  not U10976(n9391,n7104);
  nand U10977(n7104,n10495,n10579);
  nand U10978(n10579,n10580,n10581);
  or U10979(n10495,n10581,n10580);
  or U10980(n10580,n9284,n10582);
  nor U10981(n10582,n10583,n10584,n10585,n10586);
  and U10982(n10586,n10264,G21721);
  nor U10983(n10585,n9290,n7102,n7103);
  and U10984(n7103,n10587,n10588,n10589);
  nand U10985(n10588,G21594,n9101);
  nand U10986(n10587,n10590,n8737);
  not U10987(n7102,n10510);
  nand U10988(n10510,n10591,n10592,n7114);
  nand U10989(n10592,n9101,n10566);
  not U10990(n10566,G21594);
  or U10991(n10591,n10590,n9101);
  nand U10992(n10590,n10593,n10594,n10595,n10596);
  nor U10993(n10596,n10597,n10598,n10599,n10600);
  nor U10994(n10600,n10601,n10332);
  nor U10995(n10599,n10602,n10334);
  nor U10996(n10598,n10603,n10336);
  nor U10997(n10597,n10604,n10338);
  nor U10998(n10595,n10605,n10606,n10607,n10608);
  nor U10999(n10608,n10609,n10344);
  nor U11000(n10607,n10610,n10346);
  nor U11001(n10606,n10611,n10348);
  nor U11002(n10605,n10612,n10350);
  nor U11003(n10594,n10613,n10614,n10615,n10616);
  nor U11004(n10616,n10617,n10356);
  nor U11005(n10615,n10618,n10358);
  nor U11006(n10614,n10619,n10360);
  nor U11007(n10613,n10620,n10362);
  nor U11008(n10593,n10621,n10622,n10623,n10624);
  nor U11009(n10624,n10625,n10368);
  nor U11010(n10623,n10626,n10370);
  nor U11011(n10622,n10627,n10372);
  nor U11012(n10621,n10628,n10374);
  nor U11013(n10584,n10263,n9390);
  not U11014(n9390,G21753);
  nand U11015(n10583,n10629,n10630);
  nand U11016(n10630,G21594,n10504);
  nand U11017(n10629,G21626,n7590);
  nand U11018(n10573,n10041,n10631);
  nand U11019(G1015,n10632,n10633,n10634,n10635);
  nor U11020(n10635,n10636,n10637);
  nor U11021(n10637,n6921,n9399);
  nor U11022(n10636,n6943,n10638);
  nand U11023(n10634,n9401,n6912);
  nand U11024(n10633,n6931,n7117);
  or U11025(n7117,n10559,n10639);
  or U11026(n10639,n9953,n10558);
  nand U11027(n10558,n10640,n10641);
  nand U11028(n10641,n9953,n10642);
  or U11029(n10642,n10643,n10644);
  nand U11030(n10640,n10644,n10643);
  nand U11031(n10559,n10645,n10646,n10647,n10648);
  nor U11032(n10648,n10649,n10650);
  nor U11033(n10650,n10287,n10638);
  nor U11034(n10649,n9936,n7116);
  nand U11035(n10647,G21593,n10250);
  nand U11036(n10646,n9698,n10651);
  nand U11037(n10645,n10567,n10290,n7113);
  not U11038(n7113,n9698);
  nand U11039(n10632,n9698,n6933);
  nor U11040(n9698,n10482,n10652);
  and U11041(n10652,n10653,n10654);
  nor U11042(n10482,n10654,n10653);
  or U11043(n10653,n10655,n9110);
  nand U11044(n10655,n10656,n10657,n10658);
  nor U11045(n10658,n10659,n10660,n10661);
  nor U11046(n10661,n10248,n10638);
  not U11047(n10638,G21784);
  nor U11048(n10660,n10246,n9399);
  not U11049(n9399,G21625);
  and U11050(n10659,n10662,n10041);
  nand U11051(n10657,G21593,n10247);
  nand U11052(n10656,n9401,n10305);
  not U11053(n9401,n7116);
  nand U11054(n7116,n10581,n10663);
  nand U11055(n10663,n10664,n10665);
  or U11056(n10581,n10665,n10664);
  or U11057(n10664,n10666,n10248);
  nand U11058(n10666,n10667,n10668,n10669,n10670);
  nand U11059(n10670,G21752,n10316);
  nor U11060(n10669,n10671,n10672);
  and U11061(n10672,n10264,G21720);
  nor U11062(n10671,n9290,n7114,n7115);
  and U11063(n7115,n10673,n10674,n10675);
  nand U11064(n10674,G21593,n9101);
  nand U11065(n10673,n10676,n8737);
  not U11066(n7114,n10589);
  nand U11067(n10589,n10677,n10678,n10679);
  not U11068(n10679,n10675);
  or U11069(n10678,n8737,G21593);
  or U11070(n10677,n10676,n9101);
  nand U11071(n10676,n10680,n10681,n10682,n10683);
  nor U11072(n10683,n10684,n10685,n10686,n10687);
  nor U11073(n10687,n10688,n10332);
  nor U11074(n10686,n10689,n10334);
  nor U11075(n10685,n10690,n10336);
  nor U11076(n10684,n10691,n10338);
  nor U11077(n10682,n10692,n10693,n10694,n10695);
  nor U11078(n10695,n10696,n10344);
  nor U11079(n10694,n10697,n10346);
  nor U11080(n10693,n10698,n10348);
  nor U11081(n10692,n10699,n10350);
  nor U11082(n10681,n10700,n10701,n10702,n10703);
  nor U11083(n10703,n10704,n10356);
  nor U11084(n10702,n10705,n10358);
  nor U11085(n10701,n10706,n10360);
  nor U11086(n10700,n10707,n10362);
  nor U11087(n10680,n10708,n10709,n10710,n10711);
  nor U11088(n10711,n10712,n10368);
  nor U11089(n10710,n10713,n10370);
  nor U11090(n10709,n10714,n10372);
  nor U11091(n10708,n10715,n10374);
  nand U11092(n10668,G21593,n10504);
  nand U11093(n10667,G21625,n7590);
  nand U11094(n10654,n10716,n10717);
  not U11095(n10716,n10718);
  nand U11096(G1014,n10719,n10720,n10721,n10722);
  nor U11097(n10722,n10723,n10724);
  nor U11098(n10724,n6921,n9409);
  nor U11099(n10723,n6943,n7125);
  nand U11100(n10721,n7131,n6912);
  nand U11101(n10720,n6931,n7129);
  or U11102(n7129,n10644,n10725);
  or U11103(n10725,n9953,n10643);
  nand U11104(n10643,n10726,n10727);
  nand U11105(n10727,n9953,n10728);
  or U11106(n10728,n10729,n10730);
  nand U11107(n10726,n10730,n10729);
  nand U11108(n10644,n10731,n10732,n10733,n10734);
  nor U11109(n10734,n10735,n10736);
  nor U11110(n10736,n10285,n7127);
  nor U11111(n10735,n10287,n7125);
  nand U11112(n10733,n7131,n9953);
  nand U11113(n10732,n10737,n9705,n7153,n10571);
  nand U11114(n10731,n7130,n10651);
  nand U11115(n10651,n10569,n10738);
  nand U11116(n10738,n10290,n10571);
  not U11117(n10571,n10567);
  nor U11118(n10567,n10739,n7139,n9411,n9431);
  nand U11119(n10719,n7130,n6933);
  not U11120(n7130,n9411);
  or U11121(n9411,n10717,n10718);
  or U11122(n10717,n10740,n9110);
  nand U11123(n10740,n10741,n10742,n10743,n10744);
  nor U11124(n10744,n10745,n10746);
  nor U11125(n10746,n10248,n7125);
  not U11126(n7125,G21783);
  nor U11127(n10745,n10246,n9409);
  not U11128(n9409,G21624);
  nand U11129(n10743,G21592,n10247);
  nand U11130(n10742,n7131,n10305);
  not U11131(n7131,n9835);
  nand U11132(n9835,n10665,n10747);
  nand U11133(n10747,n10748,n10749);
  or U11134(n10665,n10749,n10748);
  or U11135(n10748,n10750,n10248);
  nand U11136(n10750,n10751,n10752,n10753,n10754);
  nand U11137(n10754,G21751,n10316);
  nor U11138(n10753,n10755,n10756);
  and U11139(n10756,n10264,G21719);
  nor U11140(n10755,n9290,n7126);
  nand U11141(n7126,n10757,n10675);
  nand U11142(n10675,n10758,n10759,n10760,n10761);
  nand U11143(n10761,n9101,n7127);
  not U11144(n7127,G21592);
  or U11145(n10760,n10762,n9101);
  nand U11146(n10757,n10763,n10764,n10765);
  nand U11147(n10765,n10758,n10759);
  nand U11148(n10764,G21592,n9101);
  nand U11149(n10763,n10762,n8737);
  nand U11150(n10762,n10766,n10767,n10768,n10769);
  nor U11151(n10769,n10770,n10771,n10772,n10773);
  nor U11152(n10773,n10774,n10332);
  nor U11153(n10772,n10775,n10334);
  nor U11154(n10771,n10776,n10336);
  nor U11155(n10770,n10777,n10338);
  nor U11156(n10768,n10778,n10779,n10780,n10781);
  nor U11157(n10781,n10782,n10344);
  nor U11158(n10780,n10783,n10346);
  nor U11159(n10779,n10784,n10348);
  nor U11160(n10778,n10785,n10350);
  nor U11161(n10767,n10786,n10787,n10788,n10789);
  nor U11162(n10789,n10790,n10356);
  nor U11163(n10788,n10791,n10358);
  nor U11164(n10787,n10792,n10360);
  nor U11165(n10786,n10793,n10362);
  nor U11166(n10766,n10794,n10795,n10796,n10797);
  nor U11167(n10797,n10798,n10368);
  nor U11168(n10796,n10799,n10370);
  nor U11169(n10795,n10800,n10372);
  nor U11170(n10794,n10801,n10374);
  nand U11171(n10752,G21592,n10504);
  nand U11172(n10751,G21624,n7590);
  nand U11173(n10741,n10041,n10802);
  nand U11174(G1013,n10803,n10804,n10805,n10806);
  nor U11175(n10806,n10807,n10808);
  nor U11176(n10808,n6921,n9419);
  nor U11177(n10807,n6943,n10809);
  nand U11178(n10805,n9421,n6912);
  nand U11179(n10804,n6931,n7142);
  or U11180(n7142,n10730,n10810);
  or U11181(n10810,n9953,n10729);
  nand U11182(n10729,n10811,n10812);
  nand U11183(n10812,n9953,n10813);
  or U11184(n10813,n10814,n10815);
  nand U11185(n10811,n10815,n10814);
  nand U11186(n10730,n10816,n10817,n10818,n10819);
  nor U11187(n10819,n10820,n10821);
  nor U11188(n10821,n10287,n10809);
  nor U11189(n10820,n9936,n7141);
  nand U11190(n10818,G21591,n10250);
  nand U11191(n10817,n9705,n10822);
  nand U11192(n10822,n10823,n10824);
  nand U11193(n10824,n10290,n9431);
  not U11194(n10823,n10825);
  nand U11195(n10816,n10737,n7153,n7139);
  nand U11196(n10803,n9705,n6933);
  not U11197(n9705,n7139);
  nand U11198(n7139,n10718,n10826);
  nand U11199(n10826,n10827,n10828,n10829);
  or U11200(n10829,n7590,n10830);
  nand U11201(n10718,n10831,n10832);
  nand U11202(n10832,n10827,n10828);
  nand U11203(n10827,n10833,n10834);
  or U11204(n10831,n10830,n9110);
  nand U11205(n10830,n10835,n10836,n10837);
  nor U11206(n10837,n10838,n10839,n10840);
  nor U11207(n10840,n10248,n10809);
  not U11208(n10809,G21782);
  nor U11209(n10839,n10246,n9419);
  not U11210(n9419,G21623);
  and U11211(n10838,n10841,n10041);
  nand U11212(n10836,G21591,n10247);
  nand U11213(n10835,n9421,n10305);
  not U11214(n9421,n7141);
  nand U11215(n7141,n10749,n10842);
  nand U11216(n10842,n10843,n10844);
  or U11217(n10749,n10844,n10843);
  or U11218(n10843,n10845,n10248);
  nand U11219(n10845,n10846,n10847,n10848);
  nor U11220(n10848,n10849,n10850,n10851);
  and U11221(n10851,n10264,G21718);
  nor U11222(n10850,n7140,n9290);
  or U11223(n7140,n10758,n10759);
  nand U11224(n10759,n10852,n10853);
  nand U11225(n10853,G21591,n9101);
  nand U11226(n10852,n10854,n8737);
  nand U11227(n10854,n10855,n10856,n10857,n10858);
  nor U11228(n10858,n10859,n10860,n10861,n10862);
  nor U11229(n10862,n10863,n10332);
  nor U11230(n10861,n10864,n10334);
  nor U11231(n10860,n10865,n10336);
  nor U11232(n10859,n10866,n10338);
  nor U11233(n10857,n10867,n10868,n10869,n10870);
  nor U11234(n10870,n10871,n10344);
  nor U11235(n10869,n10872,n10346);
  nor U11236(n10868,n10873,n10348);
  nor U11237(n10867,n10874,n10350);
  nor U11238(n10856,n10875,n10876,n10877,n10878);
  nor U11239(n10878,n10879,n10356);
  nor U11240(n10877,n10880,n10358);
  nor U11241(n10876,n10881,n10360);
  nor U11242(n10875,n10882,n10362);
  nor U11243(n10855,n10883,n10884,n10885,n10886);
  nor U11244(n10886,n10887,n10368);
  nor U11245(n10885,n10888,n10370);
  nor U11246(n10884,n10889,n10372);
  nor U11247(n10883,n10890,n10374);
  and U11248(n10758,n10891,n10892);
  nor U11249(n10849,n10263,n9420);
  not U11250(n9420,G21750);
  nand U11251(n10847,G21591,n10504);
  nand U11252(n10846,G21623,n7590);
  nand U11253(G1012,n10893,n10894,n10895,n10896);
  nor U11254(n10896,n10897,n10898);
  nor U11255(n10898,n6921,n9429);
  nor U11256(n10897,n6943,n7150);
  nand U11257(n10895,n7154,n6912);
  nand U11258(n10894,n6931,n7152);
  or U11259(n7152,n10815,n10899);
  or U11260(n10899,n9953,n10814);
  nand U11261(n10814,n10900,n10901);
  nand U11262(n10901,n9953,n10902);
  or U11263(n10902,n10903,n10904);
  nand U11264(n10900,n10904,n10903);
  nand U11265(n10815,n10905,n10906,n10907,n10908);
  nor U11266(n10908,n10909,n10910);
  nor U11267(n10910,n10287,n7150);
  nor U11268(n10909,n9936,n9850);
  nand U11269(n10907,G21590,n10250);
  nand U11270(n10906,n10737,n9431);
  nor U11271(n10737,n10739,n9216);
  nand U11272(n10905,n7153,n10825);
  nand U11273(n10893,n7153,n6933);
  not U11274(n7153,n9431);
  or U11275(n9431,n10911,n10834);
  nand U11276(n10834,n10912,n10913);
  nand U11277(n10913,n10914,n10915);
  nand U11278(n10912,n10916,n10917,n10041);
  nand U11279(n10911,n10828,n10833);
  nand U11280(n10833,n10918,n10919);
  nand U11281(n10919,n10041,n10920);
  or U11282(n10918,n7590,n10921);
  nand U11283(n10828,n10921,n10920,n10041);
  nand U11284(n10921,n10922,n10923,n10924,n10925);
  nor U11285(n10925,n10926,n10927);
  nor U11286(n10927,n10248,n7150);
  not U11287(n7150,G21781);
  nor U11288(n10926,n10246,n9429);
  not U11289(n9429,G21622);
  nand U11290(n10924,G21590,n10247);
  nand U11291(n10923,n7154,n10305);
  not U11292(n7154,n9850);
  nand U11293(n9850,n10844,n10928);
  nand U11294(n10928,n10929,n10930);
  or U11295(n10844,n10930,n10929);
  or U11296(n10929,n10931,n10248);
  nand U11297(n10931,n10932,n10933,n10934);
  nor U11298(n10934,n10935,n10936,n10937);
  and U11299(n10937,n10264,G21717);
  nor U11300(n10936,n7151,n9290);
  or U11301(n7151,n10891,n10892);
  nand U11302(n10892,n10938,n10939);
  nand U11303(n10939,G21590,n9101);
  nand U11304(n10938,n10940,n8737);
  nand U11305(n10940,n10941,n10942,n10943,n10944);
  nor U11306(n10944,n10945,n10946,n10947,n10948);
  nor U11307(n10948,n10949,n10332);
  nand U11308(n10332,n10950,n10951);
  nor U11309(n10947,n10952,n10334);
  nand U11310(n10334,n10950,n10953);
  nor U11311(n10946,n10954,n10336);
  nand U11312(n10336,n10951,n10955);
  nor U11313(n10945,n10956,n10338);
  nand U11314(n10338,n10955,n10953);
  nor U11315(n10943,n10957,n10958,n10959,n10960);
  nor U11316(n10960,n10961,n10344);
  nand U11317(n10344,n10962,n10951);
  nor U11318(n10959,n10963,n10346);
  nand U11319(n10346,n10962,n10953);
  nor U11320(n10958,n10964,n10348);
  nand U11321(n10348,n10965,n10951);
  nor U11322(n10951,n8916,n10966);
  nor U11323(n10957,n10967,n10350);
  nand U11324(n10350,n10965,n10953);
  nor U11325(n10953,G21561,n10966);
  nor U11326(n10942,n10968,n10969,n10970,n10971);
  nor U11327(n10971,n10972,n10356);
  nand U11328(n10356,n10973,n10965);
  nor U11329(n10970,n10974,n10358);
  nand U11330(n10358,n10975,n10965);
  nor U11331(n10965,n9161,n9183);
  nor U11332(n10969,n10976,n10360);
  nand U11333(n10360,n10973,n10962);
  nor U11334(n10968,n10977,n10362);
  nand U11335(n10362,n10975,n10962);
  nor U11336(n10962,n9183,n10978);
  not U11337(n9183,n10979);
  nor U11338(n10941,n10980,n10981,n10982,n10983);
  nor U11339(n10983,n10984,n10368);
  nand U11340(n10368,n10973,n10955);
  nor U11341(n10982,n10985,n10370);
  nand U11342(n10370,n10975,n10955);
  nor U11343(n10955,n9161,n10979);
  not U11344(n9161,n10978);
  nor U11345(n10981,n10986,n10372);
  nand U11346(n10372,n10973,n10950);
  nor U11347(n10973,n9228,G21561);
  nor U11348(n10980,n10987,n10374);
  nand U11349(n10374,n10975,n10950);
  nor U11350(n10950,n10979,n10978);
  nor U11351(n10978,n10988,n10989);
  nor U11352(n10988,n10990,n9101);
  or U11353(n10979,G21559,n10991);
  nor U11354(n10975,n9228,n8916);
  not U11355(n9228,n10966);
  nor U11356(n10966,n10992,n10993);
  nor U11357(n10993,n10994,G21559,n10995);
  not U11358(n10995,n10991);
  and U11359(n10992,n8896,n10996);
  nand U11360(n10996,n10994,n10991);
  nand U11361(n10991,n9101,n10997);
  nand U11362(n10891,n10998,n10999);
  nand U11363(n10999,n11000,G21589);
  nand U11364(n10998,n10375,n8737);
  nand U11365(n10375,n11001,n11002,n11003,n11004);
  nor U11366(n11004,n11005,n11006,n11007,n11008);
  nor U11367(n11008,n10357,n7623);
  nor U11368(n11007,n10359,n7703);
  nor U11369(n11006,n10361,n7783);
  nor U11370(n11005,n10369,n7945);
  nor U11371(n11003,n11009,n11010,n11011,n11012);
  nor U11372(n11012,n10371,n8023);
  nor U11373(n11011,n10373,n8101);
  nor U11374(n11010,n10347,n8261);
  nor U11375(n11009,n10345,n8339);
  nor U11376(n11002,n11013,n11014,n11015,n11016);
  nor U11377(n11016,n10343,n8417);
  nor U11378(n11015,n10335,n8577);
  nor U11379(n11014,n10333,n8655);
  nor U11380(n11013,n10331,n8732);
  nor U11381(n11001,n11017,n11018,n11019,n11020);
  nor U11382(n11020,n10355,n7513);
  nor U11383(n11019,n10367,n7865);
  nor U11384(n11018,n10349,n8181);
  nor U11385(n11017,n10337,n8495);
  nor U11386(n10935,n10263,n9430);
  not U11387(n9430,G21749);
  nand U11388(n10933,G21590,n10504);
  nand U11389(n10932,G21622,n7590);
  nand U11390(n10922,n10041,n11021);
  nand U11391(G1011,n11022,n11023,n11024,n11025);
  nor U11392(n11025,n11026,n11027);
  nor U11393(n11027,n6921,n9439);
  not U11394(n9439,G21621);
  nor U11395(n11026,n6943,n7162);
  nand U11396(n11024,n7167,n6912);
  nand U11397(n11023,n6931,n7165);
  or U11398(n7165,n10904,n11028);
  or U11399(n11028,n9953,n10903);
  nand U11400(n10903,n11029,n11030);
  nand U11401(n11030,n9953,n11031);
  or U11402(n11031,n11032,n11033);
  nand U11403(n11029,n11033,n11032);
  nand U11404(n10904,n11034,n11035,n11036,n11037);
  nor U11405(n11037,n11038,n11039);
  nor U11406(n11039,n10285,n7164);
  nor U11407(n11038,n10287,n7162);
  not U11408(n7162,G21780);
  nand U11409(n11036,n7167,n9953);
  nand U11410(n11035,n7179,n11040,n7191,n10739);
  nand U11411(n11034,n7166,n10825);
  nand U11412(n10825,n10569,n11041);
  nand U11413(n11041,n10290,n10739);
  or U11414(n10739,n9441,n11042,n9451,n9461);
  nand U11415(n11022,n7166,n6933);
  not U11416(n7166,n9441);
  or U11417(n9441,n10915,n10914);
  nand U11418(n10914,n11043,n11044);
  nand U11419(n11044,n10041,n10917);
  or U11420(n11043,n7590,n10916);
  nand U11421(n10916,n11045,n11046,n11047,n11048);
  nand U11422(n11048,n7167,n10305);
  not U11423(n7167,n9858);
  nand U11424(n9858,n10930,n11049);
  nand U11425(n11049,n11050,n11051);
  or U11426(n10930,n11051,n11050);
  or U11427(n11050,n11052,n10248);
  nand U11428(n11052,n11053,n11054,n11055);
  nor U11429(n11055,n11056,n11057,n11058);
  and U11430(n11058,n10264,G21716);
  nor U11431(n11057,n7163,n9290);
  and U11432(n7163,n11059,n11060);
  nand U11433(n11060,n10459,n8737);
  nand U11434(n10459,n11061,n11062,n11063,n11064);
  nor U11435(n11064,n11065,n11066,n11067,n11068);
  nor U11436(n11068,n10448,n7623);
  nor U11437(n11067,n10449,n7703);
  nor U11438(n11066,n10450,n7783);
  nor U11439(n11065,n10456,n7945);
  nor U11440(n11063,n11069,n11070,n11071,n11072);
  nor U11441(n11072,n10457,n8023);
  nor U11442(n11071,n10458,n8101);
  nor U11443(n11070,n10441,n8261);
  nor U11444(n11069,n10440,n8339);
  nor U11445(n11062,n11073,n11074,n11075,n11076);
  nor U11446(n11076,n10439,n8417);
  nor U11447(n11075,n10433,n8577);
  nor U11448(n11074,n10432,n8655);
  nor U11449(n11073,n10431,n8732);
  nor U11450(n11061,n11077,n11078,n11079,n11080);
  nor U11451(n11080,n10447,n7513);
  nor U11452(n11079,n10455,n7865);
  nor U11453(n11078,n10442,n8181);
  nor U11454(n11077,n10434,n8495);
  nand U11455(n11059,n11081,n9101);
  or U11456(n11081,n7164,n11000);
  nor U11457(n11000,n11082,n7177);
  not U11458(n7177,G21588);
  not U11459(n7164,G21589);
  nor U11460(n11056,n10263,n9440);
  not U11461(n9440,G21748);
  nand U11462(n11054,G21589,n10504);
  nand U11463(n11053,G21621,n7590);
  nand U11464(n11047,G21589,n10247);
  nand U11465(n11046,G21621,n11083);
  nand U11466(n11045,G21780,n9284);
  and U11467(n10915,n11084,n11085);
  nand U11468(G1010,n11086,n11087,n11088,n11089);
  nor U11469(n11089,n11090,n11091);
  nor U11470(n11091,n6921,n9449);
  not U11471(n9449,G21620);
  nor U11472(n11090,n6943,n7175);
  nand U11473(n11088,n7180,n6912);
  nand U11474(n11087,n6931,n7178);
  or U11475(n7178,n11033,n11092);
  or U11476(n11092,n9953,n11032);
  nand U11477(n11032,n11093,n11094);
  nand U11478(n11094,n9953,n11095);
  or U11479(n11095,n11096,n11097);
  nand U11480(n11093,n11097,n11096);
  nand U11481(n11033,n11098,n11099,n11100,n11101);
  nor U11482(n11101,n11102,n11103);
  nor U11483(n11103,n10287,n7175);
  not U11484(n7175,G21779);
  nor U11485(n11102,n9936,n9866);
  nand U11486(n11100,G21588,n10250);
  nand U11487(n11099,n7179,n11104);
  nand U11488(n11104,n11105,n11106);
  nand U11489(n11106,n10290,n9461);
  not U11490(n11105,n11107);
  nand U11491(n11098,n11040,n7191,n9451);
  not U11492(n9451,n7179);
  nand U11493(n11086,n7179,n6933);
  or U11494(n7179,n11085,n11084);
  nand U11495(n11084,n11108,n11109);
  nand U11496(n11109,n10041,n11110);
  or U11497(n11108,n7590,n11111);
  nand U11498(n11111,n11112,n11113,n11114,n11115);
  nand U11499(n11115,n7180,n10305);
  not U11500(n7180,n9866);
  nand U11501(n9866,n11051,n11116);
  nand U11502(n11116,n11117,n11118);
  or U11503(n11051,n11118,n11117);
  or U11504(n11117,n11119,n10248);
  nand U11505(n11119,n11120,n11121,n11122);
  nor U11506(n11122,n11123,n11124,n11125);
  and U11507(n11125,n10264,G21715);
  nor U11508(n11124,n7176,n9290);
  and U11509(n7176,n11126,n11127,n11128);
  or U11510(n11128,n11082,G21588);
  nand U11511(n11127,G21588,n11082,n9101);
  nand U11512(n11082,n11129,G21587);
  nand U11513(n11126,n10492,n8737);
  nand U11514(n10492,n11130,n11131,n11132,n11133);
  nor U11515(n11133,n11134,n11135,n11136,n11137);
  nor U11516(n11137,n10536,n7623);
  nor U11517(n11136,n10537,n7703);
  nor U11518(n11135,n10538,n7783);
  nor U11519(n11134,n10544,n7945);
  nor U11520(n11132,n11138,n11139,n11140,n11141);
  nor U11521(n11141,n10545,n8023);
  nor U11522(n11140,n10546,n8101);
  nor U11523(n11139,n10529,n8261);
  nor U11524(n11138,n10528,n8339);
  nor U11525(n11131,n11142,n11143,n11144,n11145);
  nor U11526(n11145,n10527,n8417);
  nor U11527(n11144,n10521,n8577);
  nor U11528(n11143,n10520,n8655);
  nor U11529(n11142,n10519,n8732);
  nor U11530(n11130,n11146,n11147,n11148,n11149);
  nor U11531(n11149,n10535,n7513);
  nor U11532(n11148,n10543,n7865);
  nor U11533(n11147,n10530,n8181);
  nor U11534(n11146,n10522,n8495);
  nor U11535(n11123,n10263,n9450);
  not U11536(n9450,G21747);
  nand U11537(n11121,G21588,n10504);
  nand U11538(n11120,G21620,n7590);
  nand U11539(n11114,G21588,n10247);
  nand U11540(n11113,G21620,n11083);
  nand U11541(n11112,G21779,n9284);
  nand U11542(n11085,n11150,n11151);
  nand U11543(n11151,n11152,n11153);
  nand U11544(n11150,n11154,n11155,n10041);
  or U11545(n11154,n11156,n7590);
  nand U11546(G1009,n11157,n11158,n11159,n11160);
  nor U11547(n11160,n11161,n11162);
  nor U11548(n11162,n6921,n9459);
  not U11549(n9459,G21619);
  nor U11550(n11161,n6943,n7188);
  nand U11551(n11159,n7192,n6912);
  nand U11552(n11158,n6931,n7190);
  or U11553(n7190,n11097,n11163);
  or U11554(n11163,n9953,n11096);
  nand U11555(n11096,n11164,n11165);
  nand U11556(n11165,n9953,n11166);
  or U11557(n11166,n11167,n11168);
  nand U11558(n11164,n11168,n11167);
  nand U11559(n11097,n11169,n11170,n11171,n11172);
  nor U11560(n11172,n11173,n11174);
  nor U11561(n11174,n10287,n7188);
  not U11562(n7188,G21778);
  nor U11563(n11173,n9936,n9874);
  nand U11564(n11171,G21587,n10250);
  nand U11565(n11170,n9461,n11040);
  nor U11566(n11040,n11042,n9216);
  not U11567(n9461,n7191);
  nand U11568(n11169,n7191,n11107);
  nand U11569(n11157,n7191,n6933);
  or U11570(n7191,n11153,n11152);
  nand U11571(n11152,n11175,n11176);
  nand U11572(n11176,n10041,n11155);
  or U11573(n11175,n7590,n11156);
  nand U11574(n11156,n11177,n11178,n11179,n11180);
  nand U11575(n11180,n7192,n10305);
  not U11576(n7192,n9874);
  nand U11577(n9874,n11118,n11181);
  nand U11578(n11181,n11182,n11183);
  or U11579(n11118,n11183,n11182);
  or U11580(n11182,n11184,n10248);
  nand U11581(n11184,n11185,n11186,n11187);
  nor U11582(n11187,n11188,n11189,n11190);
  and U11583(n11190,n10264,G21714);
  nor U11584(n11189,n7189,n9290);
  and U11585(n7189,n11191,n11192);
  nand U11586(n11192,n10631,n8737);
  nand U11587(n10631,n11193,n11194,n11195,n11196);
  nor U11588(n11196,n11197,n11198,n11199,n11200);
  nor U11589(n11200,n10618,n7623);
  nor U11590(n11199,n10619,n7703);
  nor U11591(n11198,n10620,n7783);
  nor U11592(n11197,n10626,n7945);
  nor U11593(n11195,n11201,n11202,n11203,n11204);
  nor U11594(n11204,n10627,n8023);
  nor U11595(n11203,n10628,n8101);
  nor U11596(n11202,n10611,n8261);
  nor U11597(n11201,n10610,n8339);
  nor U11598(n11194,n11205,n11206,n11207,n11208);
  nor U11599(n11208,n10609,n8417);
  nor U11600(n11207,n10603,n8577);
  nor U11601(n11206,n10602,n8655);
  nor U11602(n11205,n10601,n8732);
  nor U11603(n11193,n11209,n11210,n11211,n11212);
  nor U11604(n11212,n10617,n7513);
  nor U11605(n11211,n10625,n7865);
  nor U11606(n11210,n10612,n8181);
  nor U11607(n11209,n10604,n8495);
  nand U11608(n11191,n11213,n9101);
  or U11609(n11213,G21587,n11129);
  nor U11610(n11129,n11214,n7202);
  nor U11611(n11188,n10263,n9460);
  not U11612(n9460,G21746);
  nand U11613(n11186,G21587,n10504);
  nand U11614(n11185,G21619,n7590);
  nand U11615(n11179,G21587,n10247);
  nand U11616(n11178,G21619,n11083);
  nand U11617(n11177,G21778,n9284);
  nand U11618(n11153,n11215,n11216);
  nand U11619(n11216,n11217,n11218);
  nand U11620(n11215,n10041,n11219,n11220);
  or U11621(n11220,n11221,n9110);
  nand U11622(G1008,n11222,n11223,n11224,n11225);
  nor U11623(n11225,n11226,n11227);
  nor U11624(n11227,n6921,n9471);
  not U11625(n9471,G21618);
  nor U11626(n11226,n6943,n7200);
  nand U11627(n11224,n7205,n6912);
  nand U11628(n11223,n6931,n7203);
  or U11629(n7203,n11168,n11228);
  or U11630(n11228,n9953,n11167);
  nand U11631(n11167,n11229,n11230);
  nand U11632(n11230,n9953,n11231);
  or U11633(n11231,n11232,n11233);
  nand U11634(n11229,n11233,n11232);
  nand U11635(n11168,n11234,n11235,n11236,n11237);
  nor U11636(n11237,n11238,n11239);
  nor U11637(n11239,n10285,n7202);
  not U11638(n7202,G21586);
  nor U11639(n11238,n10287,n7200);
  not U11640(n7200,G21777);
  nand U11641(n11236,n7205,n9953);
  nand U11642(n11235,n7229,n11240,n7216,n11042);
  nand U11643(n11234,n7204,n11107);
  nand U11644(n11107,n10569,n11241);
  nand U11645(n11241,n10290,n11042);
  nand U11646(n11042,n7242,n11242,n7216,n11243);
  nor U11647(n11243,n9470,n9490);
  not U11648(n9470,n7204);
  nand U11649(n11222,n7204,n6933);
  or U11650(n7204,n11218,n11217);
  nand U11651(n11217,n11244,n11245);
  nand U11652(n11245,n10041,n11219);
  or U11653(n11244,n7590,n11221);
  nand U11654(n11221,n11246,n11247,n11248,n11249);
  nand U11655(n11249,n7205,n10305);
  not U11656(n7205,n9882);
  nand U11657(n9882,n11183,n11250);
  nand U11658(n11250,n11251,n11252);
  or U11659(n11183,n11252,n11251);
  or U11660(n11251,n11253,n10248);
  nand U11661(n11253,n11254,n11255,n11256);
  nor U11662(n11256,n11257,n11258,n11259);
  and U11663(n11259,n10264,G21713);
  nor U11664(n11258,n7201,n9290);
  and U11665(n7201,n11260,n11261,n11262);
  or U11666(n11262,n11214,G21586);
  nand U11667(n11261,G21586,n11214,n9101);
  nand U11668(n11214,n11263,G21585);
  nand U11669(n11260,n10662,n8737);
  nand U11670(n10662,n11264,n11265,n11266,n11267);
  nor U11671(n11267,n11268,n11269,n11270,n11271);
  nor U11672(n11271,n10705,n7623);
  nor U11673(n11270,n10706,n7703);
  nor U11674(n11269,n10707,n7783);
  nor U11675(n11268,n10713,n7945);
  nor U11676(n11266,n11272,n11273,n11274,n11275);
  nor U11677(n11275,n10714,n8023);
  nor U11678(n11274,n10715,n8101);
  nor U11679(n11273,n10698,n8261);
  nor U11680(n11272,n10697,n8339);
  nor U11681(n11265,n11276,n11277,n11278,n11279);
  nor U11682(n11279,n10696,n8417);
  nor U11683(n11278,n10690,n8577);
  nor U11684(n11277,n10689,n8655);
  nor U11685(n11276,n10688,n8732);
  nor U11686(n11264,n11280,n11281,n11282,n11283);
  nor U11687(n11283,n10704,n7513);
  nor U11688(n11282,n10712,n7865);
  nor U11689(n11281,n10699,n8181);
  nor U11690(n11280,n10691,n8495);
  nor U11691(n11257,n10263,n9472);
  not U11692(n9472,G21745);
  nand U11693(n11255,G21586,n10504);
  nand U11694(n11254,G21618,n7590);
  nand U11695(n11248,G21586,n10247);
  nand U11696(n11247,G21618,n11083);
  nand U11697(n11246,G21777,n9284);
  nand U11698(n11218,n11284,n11285);
  nand U11699(n11285,n11286,n11287);
  nand U11700(G1007,n11288,n11289,n11290,n11291);
  nor U11701(n11291,n11292,n11293);
  nor U11702(n11293,n6921,n9481);
  not U11703(n9481,G21617);
  nor U11704(n11292,n6943,n7213);
  nand U11705(n11290,n7217,n6912);
  nand U11706(n11289,n6931,n7215);
  or U11707(n7215,n11233,n11294);
  or U11708(n11294,n9953,n11232);
  nand U11709(n11232,n11295,n11296);
  nand U11710(n11296,n9953,n11297);
  or U11711(n11297,n11298,n11299);
  nand U11712(n11295,n11299,n11298);
  nand U11713(n11233,n11300,n11301,n11302,n11303);
  nor U11714(n11303,n11304,n11305);
  nor U11715(n11305,n10287,n7213);
  not U11716(n7213,G21776);
  nor U11717(n11304,n9936,n9890);
  nand U11718(n11302,G21585,n10250);
  nand U11719(n11301,n7216,n11306);
  nand U11720(n11306,n11307,n11308);
  nand U11721(n11308,n10290,n9490);
  nand U11722(n11300,n11240,n7229,n9480);
  nand U11723(n11288,n7216,n6933);
  not U11724(n7216,n9480);
  or U11725(n9480,n11287,n11309);
  and U11726(n11309,n11286,n11284);
  nand U11727(n11284,n10041,n11310,n11311);
  or U11728(n11311,n11312,n7590);
  nand U11729(n11286,n11313,n11314);
  nand U11730(n11314,n10041,n11310);
  or U11731(n11313,n9110,n11312);
  and U11732(n11312,n11315,n11316,n11317,n11318);
  nand U11733(n11318,n7217,n10305);
  not U11734(n7217,n9890);
  nand U11735(n9890,n11252,n11319);
  nand U11736(n11319,n11320,n11321);
  or U11737(n11252,n11321,n11320);
  or U11738(n11320,n11322,n10248);
  nand U11739(n11322,n11323,n11324,n11325);
  nor U11740(n11325,n11326,n11327,n11328);
  and U11741(n11328,n10264,G21712);
  nor U11742(n11327,n7214,n9290);
  and U11743(n7214,n11329,n11330);
  nand U11744(n11330,n10802,n8737);
  nand U11745(n10802,n11331,n11332,n11333,n11334);
  nor U11746(n11334,n11335,n11336,n11337,n11338);
  nor U11747(n11338,n10791,n7623);
  nor U11748(n11337,n10792,n7703);
  nor U11749(n11336,n10793,n7783);
  nor U11750(n11335,n10799,n7945);
  nor U11751(n11333,n11339,n11340,n11341,n11342);
  nor U11752(n11342,n10800,n8023);
  nor U11753(n11341,n10801,n8101);
  nor U11754(n11340,n10784,n8261);
  nor U11755(n11339,n10783,n8339);
  nor U11756(n11332,n11343,n11344,n11345,n11346);
  nor U11757(n11346,n10782,n8417);
  nor U11758(n11345,n10776,n8577);
  nor U11759(n11344,n10775,n8655);
  nor U11760(n11343,n10774,n8732);
  nor U11761(n11331,n11347,n11348,n11349,n11350);
  nor U11762(n11350,n10790,n7513);
  nor U11763(n11349,n10798,n7865);
  nor U11764(n11348,n10785,n8181);
  nor U11765(n11347,n10777,n8495);
  nand U11766(n11329,n11351,n9101);
  or U11767(n11351,G21585,n11263);
  nor U11768(n11263,n11352,n7227);
  not U11769(n7227,G21584);
  nor U11770(n11326,n10263,n9482);
  not U11771(n9482,G21744);
  nand U11772(n11324,G21585,n10504);
  nand U11773(n11323,G21617,n7590);
  nand U11774(n11317,G21585,n10247);
  nand U11775(n11316,G21617,n11083);
  nand U11776(n11315,G21776,n9284);
  nand U11777(n11287,n11353,n11354);
  nand U11778(n11354,n11355,n11356);
  nand U11779(G1006,n11357,n11358,n11359,n11360);
  nor U11780(n11360,n11361,n11362);
  nor U11781(n11362,n6921,n9491);
  not U11782(n9491,G21616);
  nand U11783(n11359,n7230,n6912);
  nand U11784(n11358,n6931,n7228);
  or U11785(n7228,n11299,n11363);
  or U11786(n11363,n9953,n11298);
  nand U11787(n11298,n11364,n11365);
  nand U11788(n11365,n9953,n11366);
  or U11789(n11366,n11367,n11368);
  nand U11790(n11364,n11368,n11367);
  nand U11791(n11299,n11369,n11370,n11371,n11372);
  nor U11792(n11372,n11373,n11374);
  nor U11793(n11374,n10287,n7225);
  not U11794(n7225,G21775);
  nor U11795(n11373,n9936,n9898);
  nand U11796(n11371,G21584,n10250);
  nand U11797(n11370,n11240,n9490);
  nor U11798(n11240,n9500,n11375,n9216);
  or U11799(n11369,n9490,n11307);
  nor U11800(n11307,n11376,n11377);
  nor U11801(n11377,n7242,n9216);
  nand U11802(n11357,n7229,n6933);
  not U11803(n7229,n9490);
  or U11804(n9490,n11356,n11378);
  and U11805(n11378,n11355,n11353);
  nand U11806(n11353,n10041,n11379,n11380);
  or U11807(n11380,n11381,n9110);
  nand U11808(n11355,n11382,n11383);
  nand U11809(n11383,n10041,n11379);
  or U11810(n11382,n7590,n11381);
  nand U11811(n11381,n11384,n11385,n11386,n11387);
  nand U11812(n11387,n7230,n10305);
  not U11813(n7230,n9898);
  nand U11814(n9898,n11321,n11388);
  nand U11815(n11388,n11389,n11390);
  or U11816(n11321,n11390,n11389);
  or U11817(n11389,n11391,n10248);
  nand U11818(n11391,n11392,n11393,n11394);
  nor U11819(n11394,n11395,n11396,n11397);
  and U11820(n11397,n10264,G21711);
  nor U11821(n11396,n7226,n9290);
  and U11822(n7226,n11398,n11399,n11400);
  or U11823(n11400,n11352,G21584);
  nand U11824(n11399,G21584,n11352,n9101);
  nand U11825(n11352,n11401,G21583);
  nand U11826(n11398,n10841,n8737);
  nand U11827(n10841,n11402,n11403,n11404,n11405);
  nor U11828(n11405,n11406,n11407,n11408,n11409);
  nor U11829(n11409,n10880,n7623);
  nor U11830(n11408,n10881,n7703);
  nor U11831(n11407,n10882,n7783);
  nor U11832(n11406,n10888,n7945);
  nor U11833(n11404,n11410,n11411,n11412,n11413);
  nor U11834(n11413,n10889,n8023);
  nor U11835(n11412,n10890,n8101);
  nor U11836(n11411,n10873,n8261);
  nor U11837(n11410,n10872,n8339);
  nor U11838(n11403,n11414,n11415,n11416,n11417);
  nor U11839(n11417,n10871,n8417);
  nor U11840(n11416,n10865,n8577);
  nor U11841(n11415,n10864,n8655);
  nor U11842(n11414,n10863,n8732);
  nor U11843(n11402,n11418,n11419,n11420,n11421);
  nor U11844(n11421,n10879,n7513);
  nor U11845(n11420,n10887,n7865);
  nor U11846(n11419,n10874,n8181);
  nor U11847(n11418,n10866,n8495);
  nor U11848(n11395,n10263,n9492);
  not U11849(n9492,G21743);
  nand U11850(n11393,G21584,n10504);
  nand U11851(n11392,G21616,n7590);
  nand U11852(n11386,G21584,n10247);
  nand U11853(n11385,G21616,n11083);
  nand U11854(n11384,G21775,n9284);
  nand U11855(n11356,n11422,n11423);
  nand U11856(n11423,n11424,n11425);
  not U11857(n11424,n11426);
  nand U11858(G1005,n11427,n11428,n11429,n11430);
  nor U11859(n11430,n11431,n11432);
  nor U11860(n11432,n6921,n9501);
  not U11861(n9501,G21615);
  nor U11862(n11431,n6943,n7238);
  nand U11863(n11429,n7243,n6912);
  nand U11864(n11428,n6931,n7241);
  or U11865(n7241,n11368,n11433);
  or U11866(n11433,n9953,n11367);
  nand U11867(n11367,n11434,n11435);
  nand U11868(n11435,n9953,n11436);
  or U11869(n11436,n11437,n11438);
  nand U11870(n11434,n11438,n11437);
  nand U11871(n11368,n11439,n11440,n11441,n11442);
  nor U11872(n11442,n11443,n11444);
  nor U11873(n11444,n10287,n7238);
  not U11874(n7238,G21774);
  nor U11875(n11443,n9936,n9906);
  nand U11876(n11441,G21583,n10250);
  nand U11877(n11440,n7242,n11376);
  nand U11878(n11376,n10569,n11445);
  not U11879(n11375,n11242);
  nand U11880(n11439,n10290,n11242,n9500);
  not U11881(n9500,n7242);
  nand U11882(n11242,n11446,n11447);
  nand U11883(n11447,n11448,n11449);
  nand U11884(n11448,n9510,n11450);
  or U11885(n11446,n9510,n11450);
  nand U11886(n11427,n6933,n7242);
  or U11887(n7242,n11451,n11426);
  nand U11888(n11451,n11422,n11425);
  nand U11889(n11425,n11452,n11453);
  nand U11890(n11453,n10041,n11454);
  or U11891(n11452,n9110,n11455);
  nand U11892(n11422,n10041,n11454,n11456);
  or U11893(n11456,n7590,n11455);
  and U11894(n11455,n11457,n11458,n11459,n11460);
  nand U11895(n11460,n7243,n10305);
  not U11896(n7243,n9906);
  nand U11897(n9906,n11390,n11461);
  nand U11898(n11461,n11462,n11463,n11464);
  or U11899(n11464,n9284,n11465);
  nand U11900(n11390,n11466,n11467);
  nand U11901(n11467,n11462,n11463);
  nand U11902(n11462,n11468,n11469);
  or U11903(n11466,n11465,n10248);
  nand U11904(n11465,n11470,n11471,n11472);
  nor U11905(n11472,n11473,n11474,n11475);
  and U11906(n11475,n10264,G21710);
  nor U11907(n11474,n7239,n9290);
  and U11908(n7239,n11476,n11477);
  nand U11909(n11477,n11401,n7240);
  not U11910(n7240,G21583);
  nand U11911(n11476,n11478,n11479);
  not U11912(n11479,n11401);
  nor U11913(n11401,n7251,n7254,n7252);
  or U11914(n7252,n7283,n7280,n7281);
  nand U11915(n7281,G21578,G21577,n7328);
  nor U11916(n7328,n7338,n7339);
  nand U11917(n7339,n7349,G21575);
  nor U11918(n7349,n7362,n7359,n7360);
  nand U11919(n7360,G21572,G21571,n7403);
  nor U11920(n7403,n7401,n7404);
  and U11921(n7404,n7417,n7416);
  nand U11922(n7416,G21569,n9101);
  nand U11923(n7417,n7427,G21568);
  nor U11924(n7427,n8737,n11480);
  not U11925(n7401,G21570);
  not U11926(n7359,G21573);
  not U11927(n7362,G21574);
  nand U11928(n7338,G21576,n9101);
  nand U11929(n11478,n11481,n11482);
  nand U11930(n11482,G21583,n9101);
  nand U11931(n11481,n11021,n8737);
  nand U11932(n11021,n11483,n11484,n11485,n11486);
  nor U11933(n11486,n11487,n11488,n11489,n11490);
  nor U11934(n11490,n10974,n7623);
  nand U11935(n7623,n11491,n11492);
  nor U11936(n11489,n10976,n7703);
  nand U11937(n7703,n11493,n11494);
  nor U11938(n11488,n10977,n7783);
  nand U11939(n7783,n11491,n11494);
  nor U11940(n11487,n10985,n7945);
  nand U11941(n7945,n11492,n11495);
  nor U11942(n11485,n11496,n11497,n11498,n11499);
  nor U11943(n11499,n10986,n8023);
  nand U11944(n8023,n11500,n11494);
  nor U11945(n11498,n10987,n8101);
  nand U11946(n8101,n11494,n11495);
  nor U11947(n11494,n9157,n11501);
  nor U11948(n11497,n10964,n8261);
  nand U11949(n8261,n11502,n11491);
  nor U11950(n11496,n10963,n8339);
  nand U11951(n8339,n11503,n11493);
  nor U11952(n11484,n11504,n11505,n11506,n11507);
  nor U11953(n11507,n10961,n8417);
  nand U11954(n8417,n11503,n11491);
  nor U11955(n11491,n11508,n9135);
  nor U11956(n11506,n10954,n8577);
  nand U11957(n8577,n11502,n11495);
  nor U11958(n11505,n10952,n8655);
  nand U11959(n8655,n11500,n11503);
  nor U11960(n11504,n10949,n8732);
  nand U11961(n8732,n11503,n11495);
  nor U11962(n11495,n9135,n9180);
  nor U11963(n11503,n9198,n9157);
  nor U11964(n11483,n11509,n11510,n11511,n11512);
  nor U11965(n11512,n10972,n7513);
  nand U11966(n7513,n11493,n11492);
  nor U11967(n11511,n10984,n7865);
  nand U11968(n7865,n11500,n11492);
  nor U11969(n11492,n11501,n11513);
  not U11970(n11501,n9198);
  nor U11971(n11510,n10967,n8181);
  nand U11972(n8181,n11502,n11493);
  nor U11973(n11493,n11508,n11514);
  nor U11974(n11509,n10956,n8495);
  nand U11975(n8495,n11500,n11502);
  nor U11976(n11502,n9198,n11513);
  not U11977(n11513,n9157);
  nor U11978(n11500,n9180,n11514);
  not U11979(n11514,n9135);
  nor U11980(n11473,n10263,n9502);
  not U11981(n9502,G21742);
  not U11982(n10263,n10316);
  nand U11983(n11471,G21583,n10504);
  nand U11984(n11470,G21615,n7590);
  nand U11985(n11459,G21583,n10247);
  nand U11986(n11458,G21615,n11083);
  nand U11987(n11457,G21774,n9284);
  nand U11988(G1004,n11515,n11516,n11517,n11518);
  nor U11989(n11518,n11519,n11520);
  nor U11990(n11520,n6921,n9511);
  not U11991(n9511,G21614);
  nor U11992(n11519,n6943,n7257);
  nand U11993(n11517,n7260,n6912);
  nand U11994(n11516,n6931,n7258);
  or U11995(n7258,n11438,n11521);
  or U11996(n11521,n9953,n11437);
  nand U11997(n11437,n11522,n11523);
  nand U11998(n11523,n9953,n11524);
  or U11999(n11524,n11525,n11526);
  nand U12000(n11522,n11526,n11525);
  nand U12001(n11438,n11527,n11528,n11529,n11530);
  nor U12002(n11530,n11531,n11532);
  nor U12003(n11532,n10285,n7254);
  not U12004(n7254,G21582);
  nor U12005(n11531,n10287,n7257);
  not U12006(n7257,G21773);
  nand U12007(n11529,n7260,n9953);
  or U12008(n11533,n11450,n11534);
  or U12009(n11534,n11449,n7259);
  nand U12010(n11450,n11535,n11536);
  nand U12011(n11536,n11537,n11538);
  or U12012(n11538,n9520,n11539);
  nand U12013(n11535,n11539,n9520);
  nand U12014(n11527,n7259,n10239);
  nand U12015(n11515,n7259,n6933);
  not U12016(n7259,n9510);
  nand U12017(n9510,n11426,n11540);
  nand U12018(n11540,n11541,n11542);
  or U12019(n11541,n7590,n11543);
  nand U12020(n11426,n11544,n11545);
  or U12021(n11544,n11543,n9110);
  nand U12022(n11543,n11546,n11547,n11548,n11549);
  nand U12023(n11549,n7260,n10305);
  or U12024(n7260,n11469,n11550);
  and U12025(n11550,n11468,n11463);
  nand U12026(n11463,n11551,n11449,n9783);
  nand U12027(n11468,n11552,n11553);
  nand U12028(n11553,n9783,n11449);
  nand U12029(n11449,n11554,n11555,n11556,n11557);
  nor U12030(n11557,n11558,n11559,n11560,n11561);
  nor U12031(n11561,n10333,n11562);
  nor U12032(n11560,n10335,n11563);
  nor U12033(n11559,n10337,n11564);
  nor U12034(n11558,n10345,n11565);
  nor U12035(n11556,n11566,n11567,n11568,n11569);
  nor U12036(n11569,n10347,n11570);
  nor U12037(n11568,n10349,n11571);
  nor U12038(n11567,n10357,n11572);
  nor U12039(n11566,n10359,n11573);
  nor U12040(n11555,n11574,n11575,n11576,n11577);
  nor U12041(n11577,n10361,n11578);
  nor U12042(n11576,n10369,n11579);
  nor U12043(n11575,n10371,n11580);
  nor U12044(n11574,n10373,n11581);
  nor U12045(n11554,n11582,n11583,n11584,n11585);
  nor U12046(n11585,n10331,n11586);
  nor U12047(n11584,n10343,n11587);
  nor U12048(n11583,n10355,n11588);
  nor U12049(n11582,n10367,n11589);
  or U12050(n11552,n9284,n11551);
  nand U12051(n11551,n11590,n11591,n11592,n11593);
  nand U12052(n11593,G21709,n10264);
  nand U12053(n11592,G21741,n10316);
  nand U12054(n11591,G21582,n10504);
  nand U12055(n11590,G21614,n7590);
  nand U12056(n11469,n11594,n11595);
  nand U12057(n11595,n11596,n11597);
  nand U12058(n11548,G21582,n10247);
  nand U12059(n11547,G21614,n11083);
  nand U12060(n11546,G21773,n9284);
  nand U12061(G1003,n11598,n11599,n11600,n11601);
  nor U12062(n11601,n11602,n11603);
  nor U12063(n11603,n6921,n9521);
  not U12064(n9521,G21613);
  nor U12065(n11602,n6943,n7269);
  nand U12066(n11600,n7272,n6912);
  nand U12067(n11599,n6931,n7270);
  or U12068(n7270,n11526,n11604);
  or U12069(n11604,n9953,n11525);
  nand U12070(n11525,n11605,n11606);
  nand U12071(n11606,n9953,n11607);
  or U12072(n11607,n11608,n11609);
  nand U12073(n11605,n11609,n11608);
  nand U12074(n11526,n11610,n11611,n11612,n11613);
  nor U12075(n11613,n11614,n11615);
  nor U12076(n11615,n10285,n7251);
  not U12077(n7251,G21581);
  nor U12078(n11614,n10287,n7269);
  not U12079(n7269,G21772);
  nand U12080(n11612,n7272,n9953);
  or U12081(n11616,n11539,n11617);
  or U12082(n11617,n11537,n9520);
  not U12083(n11537,n11618);
  nand U12084(n11539,n11619,n11620);
  nand U12085(n11620,n11621,n11622);
  or U12086(n11622,n11623,n9530);
  not U12087(n11621,n11624);
  nand U12088(n11619,n9530,n11623);
  nand U12089(n11610,n7271,n10239);
  nand U12090(n11598,n7271,n6933);
  not U12091(n7271,n9520);
  nand U12092(n9520,n11542,n11625);
  nand U12093(n11625,n11626,n11627);
  not U12094(n11542,n11545);
  nor U12095(n11545,n11627,n11626);
  or U12096(n11626,n11628,n9110);
  nand U12097(n11628,n11629,n11630,n11631,n11632);
  nand U12098(n11632,n7272,n10305);
  or U12099(n7272,n11597,n11633);
  and U12100(n11633,n11594,n11596);
  nand U12101(n11596,n11634,n11635);
  nand U12102(n11635,n9783,n11618);
  or U12103(n11634,n9284,n11636);
  nand U12104(n11594,n11636,n11618,n9783);
  nand U12105(n11618,n11637,n11638,n11639,n11640);
  nor U12106(n11640,n11641,n11642,n11643,n11644);
  nor U12107(n11644,n10456,n11579);
  nor U12108(n11643,n10455,n11589);
  nor U12109(n11642,n10447,n11588);
  nor U12110(n11641,n10439,n11587);
  nor U12111(n11639,n11645,n11646,n11647,n11648);
  nor U12112(n11648,n10448,n11572);
  nor U12113(n11647,n10442,n11571);
  nor U12114(n11646,n10458,n11581);
  nor U12115(n11645,n10457,n11580);
  nor U12116(n11638,n11649,n11650,n11651,n11652);
  nor U12117(n11652,n10440,n11565);
  nor U12118(n11651,n10434,n11564);
  nor U12119(n11650,n10433,n11563);
  nor U12120(n11649,n10449,n11573);
  nor U12121(n11637,n11653,n11654,n11655,n11656);
  nor U12122(n11656,n10431,n11586);
  nor U12123(n11655,n10432,n11562);
  nor U12124(n11654,n10441,n11570);
  nor U12125(n11653,n10450,n11578);
  nand U12126(n11636,n11657,n11658,n11659,n11660);
  nand U12127(n11660,G21708,n10264);
  nand U12128(n11659,G21740,n10316);
  nand U12129(n11658,G21581,n10504);
  nand U12130(n11657,G21613,n7590);
  nand U12131(n11597,n11661,n11662);
  nand U12132(n11662,n11663,n11664);
  nand U12133(n11631,G21581,n10247);
  nand U12134(n11630,G21613,n11083);
  nand U12135(n11629,G21772,n9284);
  or U12136(n11627,n11665,n11666);
  nand U12137(G1002,n11667,n11668,n11669,n11670);
  nor U12138(n11670,n11671,n11672);
  nor U12139(n11672,n6921,n9531);
  not U12140(n9531,G21612);
  nor U12141(n11671,n6943,n7286);
  nand U12142(n11669,n7289,n6912);
  nand U12143(n11668,n6931,n7287);
  or U12144(n7287,n11609,n11673);
  or U12145(n11673,n9953,n11608);
  nand U12146(n11608,n11674,n11675);
  nand U12147(n11675,n9953,n11676);
  or U12148(n11676,n11677,n11678);
  nand U12149(n11674,n11678,n11677);
  nand U12150(n11609,n11679,n11680,n11681,n11682);
  nor U12151(n11682,n11683,n11684);
  nor U12152(n11684,n10285,n7283);
  not U12153(n7283,G21580);
  nor U12154(n11683,n10287,n7286);
  not U12155(n7286,G21771);
  nand U12156(n11681,n7289,n9953);
  nand U12157(n11680,n10290,n11685);
  or U12158(n11685,n9530,n11686);
  or U12159(n11686,n11623,n11624);
  nand U12160(n11623,n11687,n11688);
  nand U12161(n11688,n11689,n11690);
  or U12162(n11690,n9540,n11691);
  nand U12163(n11687,n11691,n9540);
  nand U12164(n11679,n7288,n10239);
  nand U12165(n11667,n7288,n6933);
  not U12166(n7288,n9530);
  or U12167(n9530,n11665,n11666);
  or U12168(n11666,n11692,n9110);
  nand U12169(n11692,n11693,n11694,n11695,n11696);
  nand U12170(n11696,n7289,n10305);
  or U12171(n7289,n11664,n11697);
  and U12172(n11697,n11663,n11661);
  nand U12173(n11661,n11698,n11624,n9783);
  nand U12174(n11663,n11699,n11700);
  nand U12175(n11700,n9783,n11624);
  nand U12176(n11624,n11701,n11702,n11703,n11704);
  nor U12177(n11704,n11705,n11706,n11707,n11708);
  nor U12178(n11708,n10544,n11579);
  nor U12179(n11707,n10543,n11589);
  nor U12180(n11706,n10535,n11588);
  nor U12181(n11705,n10527,n11587);
  nor U12182(n11703,n11709,n11710,n11711,n11712);
  nor U12183(n11712,n10536,n11572);
  nor U12184(n11711,n10530,n11571);
  nor U12185(n11710,n10546,n11581);
  nor U12186(n11709,n10545,n11580);
  nor U12187(n11702,n11713,n11714,n11715,n11716);
  nor U12188(n11716,n10528,n11565);
  nor U12189(n11715,n10522,n11564);
  nor U12190(n11714,n10521,n11563);
  nor U12191(n11713,n10537,n11573);
  nor U12192(n11701,n11717,n11718,n11719,n11720);
  nor U12193(n11720,n10519,n11586);
  nor U12194(n11719,n10520,n11562);
  nor U12195(n11718,n10529,n11570);
  nor U12196(n11717,n10538,n11578);
  or U12197(n11699,n9284,n11698);
  nand U12198(n11698,n11721,n11722,n11723,n11724);
  nand U12199(n11724,G21707,n10264);
  nand U12200(n11723,G21739,n10316);
  nand U12201(n11722,G21580,n10504);
  nand U12202(n11721,G21612,n7590);
  nand U12203(n11664,n11725,n11726);
  nand U12204(n11726,n11727,n11728);
  nand U12205(n11695,G21580,n10247);
  nand U12206(n11694,G21612,n11083);
  nand U12207(n11693,G21771,n9284);
  nand U12208(G1001,n11729,n11730,n11731,n11732);
  nor U12209(n11732,n11733,n11734);
  nor U12210(n11734,n6921,n9541);
  not U12211(n9541,G21611);
  nor U12212(n11733,n6943,n7298);
  nand U12213(n11731,n7301,n6912);
  nand U12214(n11730,n6931,n7299);
  or U12215(n7299,n11678,n11735);
  or U12216(n11735,n9953,n11677);
  nand U12217(n11677,n11736,n11737);
  nand U12218(n11737,n9953,n11738);
  nand U12219(n11738,n11739,n11740);
  nand U12220(n11736,n11741,n11742);
  nand U12221(n11678,n11743,n11744,n11745,n11746);
  nor U12222(n11746,n11747,n11748);
  nor U12223(n11748,n10285,n7280);
  not U12224(n7280,G21579);
  nor U12225(n11747,n10287,n7298);
  not U12226(n7298,G21770);
  nand U12227(n11745,n7301,n9953);
  or U12228(n11749,n11691,n11750);
  or U12229(n11750,n11689,n9540);
  not U12230(n11689,n11751);
  nand U12231(n11691,n11752,n11753);
  nand U12232(n11753,n11754,n11755);
  or U12233(n11755,n9550,n11756);
  nand U12234(n11752,n11756,n9550);
  nand U12235(n11743,n7300,n10239);
  not U12236(n10239,n10569);
  nand U12237(n11729,n7300,n6933);
  not U12238(n7300,n9540);
  nand U12239(n9540,n11757,n11665);
  or U12240(n11665,n11758,n11759);
  nand U12241(n11757,n11759,n11758);
  or U12242(n11759,n11760,n9110);
  nand U12243(n11760,n11761,n11762,n11763,n11764);
  nand U12244(n11764,n7301,n10305);
  or U12245(n7301,n11727,n11765);
  and U12246(n11765,n11728,n11725);
  nand U12247(n11725,n11766,n11751,n9783);
  nand U12248(n11728,n11767,n11768);
  nand U12249(n11768,n9783,n11751);
  nand U12250(n11751,n11769,n11770,n11771,n11772);
  nor U12251(n11772,n11773,n11774,n11775,n11776);
  nor U12252(n11776,n10626,n11579);
  nor U12253(n11775,n10625,n11589);
  nor U12254(n11774,n10617,n11588);
  nor U12255(n11773,n10609,n11587);
  nor U12256(n11771,n11777,n11778,n11779,n11780);
  nor U12257(n11780,n10618,n11572);
  nor U12258(n11779,n10612,n11571);
  nor U12259(n11778,n10628,n11581);
  nor U12260(n11777,n10627,n11580);
  nor U12261(n11770,n11781,n11782,n11783,n11784);
  nor U12262(n11784,n10610,n11565);
  nor U12263(n11783,n10604,n11564);
  nor U12264(n11782,n10603,n11563);
  nor U12265(n11781,n10619,n11573);
  nor U12266(n11769,n11785,n11786,n11787,n11788);
  nor U12267(n11788,n10601,n11586);
  nor U12268(n11787,n10602,n11562);
  nor U12269(n11786,n10611,n11570);
  nor U12270(n11785,n10620,n11578);
  or U12271(n11767,n9284,n11766);
  nand U12272(n11766,n11789,n11790,n11791,n11792);
  nand U12273(n11792,G21706,n10264);
  nand U12274(n11791,G21738,n10316);
  nand U12275(n11790,G21579,n10504);
  nand U12276(n11789,G21611,n7590);
  nand U12277(n11727,n11793,n11794);
  nand U12278(n11794,n11795,n11796);
  nand U12279(n11763,G21579,n10247);
  nand U12280(n11762,G21611,n11083);
  nand U12281(n11761,G21770,n9284);
  nand U12282(G1000,n11797,n11798,n11799,n11800);
  nor U12283(n11800,n11801,n11802);
  nor U12284(n11802,n6921,n9551);
  not U12285(n9551,G21610);
  nor U12286(n11801,n6917,n9550);
  nand U12287(n11799,G21769,n6920);
  not U12288(n6920,n6943);
  nand U12289(n6943,n8824,n6921);
  nand U12290(n11798,n7315,n6931);
  nand U12291(n6919,G21428,n6921);
  and U12292(n7315,n11803,n11804);
  nand U12293(n11804,n11805,n9936);
  or U12294(n11805,n9937,n11739);
  not U12295(n11739,n11742);
  nand U12296(n11803,n11806,n9953);
  or U12297(n11806,n11742,n11740);
  nor U12298(n11740,n9939,n11741);
  not U12299(n11741,n9937);
  nand U12300(n9937,n11807,n11808);
  nand U12301(n11808,n11809,n9936);
  nand U12302(n11809,n9940,n9939);
  nor U12303(n9940,n9952,n11810);
  nand U12304(n11807,n9952,n11810);
  not U12305(n11810,n9949);
  nand U12306(n9949,n11811,n11812);
  nand U12307(n11812,n9953,n11813);
  or U12308(n11813,n9960,n9958);
  nand U12309(n11811,n9958,n9960);
  nand U12310(n9960,n9967,n11814);
  nand U12311(n11814,n9965,n9968);
  or U12312(n9968,n11815,n11816);
  nand U12313(n9965,n9977,n9976);
  nand U12314(n9976,n11817,n11818);
  or U12315(n11817,n11819,n9936);
  nand U12316(n9977,n9981,n11820);
  nand U12317(n11820,n9980,n9979);
  nand U12318(n9979,n11821,n11822);
  nand U12319(n9980,n9988,n9986);
  nand U12320(n9986,n9995,n11823);
  nand U12321(n11823,n9996,n9993);
  nand U12322(n9993,n10005,n11824);
  nand U12323(n11824,n10007,n10006);
  nand U12324(n10006,n11825,n11826);
  or U12325(n11826,n9953,n11827);
  not U12326(n11825,n11828);
  nand U12327(n10007,n10020,n10017);
  nand U12328(n10017,n11829,n11830);
  or U12329(n11829,n11831,n9936);
  nand U12330(n10020,n10018,n11832);
  nand U12331(n11832,n10016,n10015);
  nand U12332(n10015,n11833,n11834);
  nand U12333(n10016,n10027,n10025);
  nand U12334(n10025,n10034,n11835);
  nand U12335(n11835,n9953,n10033);
  nand U12336(n10033,n11836,n11837);
  or U12337(n11837,n9953,n11838);
  not U12338(n11836,n11839);
  nand U12339(n10034,n11840,n11839);
  nand U12340(n11839,n11841,n11842,n11843,n11844);
  nor U12341(n11844,n11845,n7482);
  nor U12342(n11845,n7447,n9936);
  nand U12343(n11843,G21567,n10250);
  nand U12344(n11842,n7033,n11846);
  nand U12345(n11841,n10249,G21758);
  or U12346(n11840,n11838,n9936);
  nand U12347(n11838,n11847,n11848,n11849,n11850);
  nor U12348(n11850,n9217,n11851,n11852,n11853);
  nor U12349(n11853,n11854,n9216);
  nor U12350(n11854,n11855,n11856,n11857,n11858);
  nand U12351(n11858,n11859,n11860,n11861,n11862);
  nand U12352(n11862,n11863,G21556);
  nand U12353(n11861,n11864,G21548);
  nand U12354(n11860,n11865,G21540);
  nand U12355(n11859,n11866,G21532);
  nand U12356(n11857,n11867,n11868,n11869,n11870);
  nand U12357(n11870,n11871,G21524);
  nand U12358(n11869,n11872,G21516);
  nand U12359(n11868,n11873,G21508);
  nand U12360(n11867,n11874,G21500);
  nand U12361(n11856,n11875,n11876,n11877,n11878);
  nand U12362(n11878,n11879,G21492);
  nand U12363(n11877,n11880,G21484);
  nand U12364(n11876,n11881,G21476);
  nand U12365(n11875,n11882,G21468);
  nand U12366(n11855,n11883,n11884,n11885,n11886);
  nand U12367(n11886,n11887,G21460);
  nand U12368(n11885,n11888,G21452);
  nand U12369(n11884,n11889,G21444);
  nand U12370(n11883,n11890,G21436);
  nor U12371(n11852,n11891,n11892,n11893,n11894);
  nand U12372(n11894,n9953,n11895,n11896,n11897);
  nand U12373(n11897,n11898,G21524);
  nand U12374(n11896,n11899,G21468);
  nand U12375(n11895,n11900,G21436);
  nand U12376(n11893,n11901,n11902,n11903,n11904);
  nand U12377(n11904,n11905,G21556);
  nand U12378(n11903,n11906,G21492);
  nand U12379(n11902,n11907,G21484);
  nand U12380(n11901,n11908,G21476);
  nand U12381(n11892,n11909,n11910,n11911,n11912);
  nand U12382(n11912,n11913,G21460);
  nand U12383(n11911,n11914,G21452);
  nand U12384(n11910,n11915,G21444);
  nand U12385(n11909,n11916,G21500);
  nand U12386(n11891,n11917,n11918,n11919,n11920);
  nor U12387(n11920,n11921,n11922);
  nor U12388(n11922,n10986,n11923);
  nor U12389(n11921,n10985,n11924);
  nand U12390(n11919,n11925,G21532);
  nand U12391(n11918,n11926,G21540);
  nand U12392(n11917,n11927,G21548);
  nand U12393(n11849,G21561,n7482);
  nand U12394(n11848,n11928,n11929);
  nand U12395(n11929,n11930,n11931,n11932,n11933);
  nor U12396(n11933,n11934,n11935,n11936,n11937);
  nor U12397(n11937,n10952,n8714);
  nor U12398(n11936,n10954,n8636);
  nor U12399(n11935,n10956,n8554);
  nor U12400(n11934,n10963,n8398);
  nor U12401(n11932,n11938,n11939,n11940,n11941);
  nor U12402(n11941,n10964,n8320);
  nor U12403(n11940,n10967,n8240);
  nor U12404(n11939,n10986,n8082);
  nor U12405(n11938,n10985,n8004);
  nor U12406(n11931,n11942,n11943,n11944,n11945);
  nor U12407(n11945,n10984,n7924);
  nor U12408(n11944,n10976,n7762);
  nor U12409(n11943,n10974,n7682);
  nor U12410(n11942,n10972,n7596);
  nor U12411(n11930,n11946,n11947,n11948,n11949);
  nor U12412(n11949,n10949,n8829);
  nor U12413(n11948,n10961,n8476);
  nor U12414(n11947,n10987,n8160);
  nor U12415(n11946,n10977,n7842);
  nand U12416(n11847,n11950,n11454);
  nand U12417(n11454,n11951,n11952,n11953,n11954);
  nor U12418(n11954,n11955,n11956,n11957,n11958);
  nor U12419(n11958,n10952,n11959);
  nor U12420(n11957,n10954,n11960);
  nor U12421(n11956,n10956,n11961);
  nor U12422(n11955,n10963,n11962);
  nor U12423(n11953,n11963,n11964,n11965,n11966);
  nor U12424(n11966,n10964,n11967);
  nor U12425(n11965,n10967,n11968);
  nor U12426(n11964,n10986,n11969);
  nor U12427(n11963,n10985,n11970);
  nor U12428(n11952,n11971,n11972,n11973,n11974);
  nor U12429(n11974,n10984,n11975);
  nor U12430(n11973,n10976,n11976);
  nor U12431(n11972,n10974,n11977);
  nor U12432(n11971,n10972,n11978);
  nor U12433(n11951,n11979,n11980,n11981,n11982);
  nor U12434(n11982,n10949,n11983);
  nor U12435(n11981,n10961,n11984);
  nor U12436(n11980,n10987,n11985);
  nor U12437(n11979,n10977,n11986);
  or U12438(n10027,n11834,n11833);
  or U12439(n11833,n11987,n9936);
  nand U12440(n11987,n11988,n11989,n11990,n11991);
  nor U12441(n11991,n9219,n11992,n11993,n11994);
  nor U12442(n11994,n11995,n9216);
  nor U12443(n11995,n11996,n11997,n11998,n11999);
  nand U12444(n11999,n12000,n12001,n12002,n12003);
  nand U12445(n12003,n11863,G21555);
  nand U12446(n12002,n11864,G21547);
  nand U12447(n12001,n11865,G21539);
  nand U12448(n12000,n11866,G21531);
  nand U12449(n11998,n12004,n12005,n12006,n12007);
  nand U12450(n12007,n11871,G21523);
  nand U12451(n12006,n11872,G21515);
  nand U12452(n12005,n11873,G21507);
  nand U12453(n12004,n11874,G21499);
  nand U12454(n11997,n12008,n12009,n12010,n12011);
  nand U12455(n12011,n11879,G21491);
  nand U12456(n12010,n11880,G21483);
  nand U12457(n12009,n11881,G21475);
  nand U12458(n12008,n11882,G21467);
  nand U12459(n11996,n12012,n12013,n12014,n12015);
  nand U12460(n12015,n11887,G21459);
  nand U12461(n12014,n11888,G21451);
  nand U12462(n12013,n11889,G21443);
  nand U12463(n12012,n11890,G21435);
  nor U12464(n11993,n12016,n12017,n12018,n12019);
  nand U12465(n12019,n9953,n12020,n12021,n12022);
  nand U12466(n12022,n11898,G21523);
  not U12467(n11898,n12023);
  nand U12468(n12021,n11899,G21467);
  not U12469(n11899,n12024);
  nand U12470(n12020,n11900,G21435);
  not U12471(n11900,n12025);
  nand U12472(n12018,n12026,n12027,n12028,n12029);
  nand U12473(n12029,n11905,G21555);
  not U12474(n11905,n12030);
  nand U12475(n12028,n11906,G21491);
  not U12476(n11906,n12031);
  nand U12477(n12027,n11907,G21483);
  not U12478(n11907,n12032);
  nand U12479(n12026,n11908,G21475);
  not U12480(n11908,n12033);
  nand U12481(n12017,n12034,n12035,n12036,n12037);
  nand U12482(n12037,n11913,G21459);
  not U12483(n11913,n12038);
  nand U12484(n12036,n11914,G21451);
  not U12485(n11914,n12039);
  nand U12486(n12035,n11915,G21443);
  not U12487(n11915,n12040);
  nand U12488(n12034,n11916,G21499);
  not U12489(n11916,n12041);
  nand U12490(n12016,n12042,n12043,n12044,n12045);
  nor U12491(n12045,n12046,n12047);
  nor U12492(n12047,n10889,n11923);
  nor U12493(n12046,n10888,n11924);
  nand U12494(n12044,n11925,G21531);
  not U12495(n11925,n12048);
  nand U12496(n12043,n11926,G21539);
  not U12497(n11926,n12049);
  nand U12498(n12042,n11927,G21547);
  not U12499(n11927,n12050);
  nand U12500(n11990,G21560,n7482);
  nand U12501(n11989,n11928,n12051);
  nand U12502(n12051,n12052,n12053,n12054,n12055);
  nor U12503(n12055,n12056,n12057,n12058,n12059);
  nor U12504(n12059,n10864,n8714);
  nor U12505(n12058,n10865,n8636);
  nor U12506(n12057,n10866,n8554);
  nor U12507(n12056,n10872,n8398);
  nor U12508(n12054,n12060,n12061,n12062,n12063);
  nor U12509(n12063,n10873,n8320);
  nor U12510(n12062,n10874,n8240);
  nor U12511(n12061,n10889,n8082);
  nor U12512(n12060,n10888,n8004);
  nor U12513(n12053,n12064,n12065,n12066,n12067);
  nor U12514(n12067,n10887,n7924);
  nor U12515(n12066,n10881,n7762);
  nor U12516(n12065,n10880,n7682);
  nor U12517(n12064,n10879,n7596);
  nor U12518(n12052,n12068,n12069,n12070,n12071);
  nor U12519(n12071,n10863,n8829);
  nor U12520(n12070,n10871,n8476);
  nor U12521(n12069,n10890,n8160);
  nor U12522(n12068,n10882,n7842);
  nand U12523(n11988,n11950,n11379);
  nand U12524(n11379,n12072,n12073,n12074,n12075);
  nor U12525(n12075,n12076,n12077,n12078,n12079);
  nor U12526(n12079,n10864,n11959);
  nor U12527(n12078,n10865,n11960);
  nor U12528(n12077,n10866,n11961);
  nor U12529(n12076,n10872,n11962);
  nor U12530(n12074,n12080,n12081,n12082,n12083);
  nor U12531(n12083,n10873,n11967);
  nor U12532(n12082,n10874,n11968);
  nor U12533(n12081,n10889,n11969);
  nor U12534(n12080,n10888,n11970);
  nor U12535(n12073,n12084,n12085,n12086,n12087);
  nor U12536(n12087,n10887,n11975);
  nor U12537(n12086,n10881,n11976);
  nor U12538(n12085,n10880,n11977);
  nor U12539(n12084,n10879,n11978);
  nor U12540(n12072,n12088,n12089,n12090,n12091);
  nor U12541(n12091,n10863,n11983);
  nor U12542(n12090,n10871,n11984);
  nor U12543(n12089,n10890,n11985);
  nor U12544(n12088,n10882,n11986);
  nand U12545(n11834,n12092,n12093,n12094,n12095);
  nand U12546(n12095,n7022,n11846);
  nand U12547(n12094,n10249,G21759);
  nand U12548(n12093,G21568,n10250);
  nand U12549(n12092,n9953,n7020);
  nand U12550(n10018,n12096,n12097);
  or U12551(n12097,n9953,n11831);
  nand U12552(n11831,n12098,n12099,n12100,n12101);
  nor U12553(n12101,n12102,n12103,n12104);
  and U12554(n12104,n11310,n11950);
  nand U12555(n11310,n12105,n12106,n12107,n12108);
  nor U12556(n12108,n12109,n12110,n12111,n12112);
  nor U12557(n12112,n10775,n11959);
  nor U12558(n12111,n10776,n11960);
  nor U12559(n12110,n10777,n11961);
  nor U12560(n12109,n10783,n11962);
  nor U12561(n12107,n12113,n12114,n12115,n12116);
  nor U12562(n12116,n10784,n11967);
  nor U12563(n12115,n10785,n11968);
  nor U12564(n12114,n10800,n11969);
  nor U12565(n12113,n10799,n11970);
  nor U12566(n12106,n12117,n12118,n12119,n12120);
  nor U12567(n12120,n10798,n11975);
  nor U12568(n12119,n10792,n11976);
  nor U12569(n12118,n10791,n11977);
  nor U12570(n12117,n10790,n11978);
  nor U12571(n12105,n12121,n12122,n12123,n12124);
  nor U12572(n12124,n10774,n11983);
  nor U12573(n12123,n10782,n11984);
  nor U12574(n12122,n10801,n11985);
  nor U12575(n12121,n10793,n11986);
  nor U12576(n12103,n12125,n9216);
  nor U12577(n12125,n12126,n12127,n12128,n12129);
  nand U12578(n12129,n12130,n12131,n12132,n12133);
  nand U12579(n12133,n11863,G21554);
  nand U12580(n12132,n11864,G21546);
  nand U12581(n12131,n11865,G21538);
  nand U12582(n12130,n11866,G21530);
  nand U12583(n12128,n12134,n12135,n12136,n12137);
  nand U12584(n12137,n11871,G21522);
  nand U12585(n12136,n11872,G21514);
  nand U12586(n12135,n11873,G21506);
  nand U12587(n12134,n11874,G21498);
  nand U12588(n12127,n12138,n12139,n12140,n12141);
  nand U12589(n12141,n11879,G21490);
  nand U12590(n12140,n11880,G21482);
  nand U12591(n12139,n11881,G21474);
  nand U12592(n12138,n11882,G21466);
  nand U12593(n12126,n12142,n12143,n12144,n12145);
  nand U12594(n12145,n11887,G21458);
  nand U12595(n12144,n11888,G21450);
  nand U12596(n12143,n11889,G21442);
  nand U12597(n12142,n11890,G21434);
  nor U12598(n12102,n7465,n8919);
  nand U12599(n12100,n11928,n12146);
  nand U12600(n12146,n12147,n12148,n12149,n12150);
  nor U12601(n12150,n12151,n12152,n12153,n12154);
  nor U12602(n12154,n10775,n8714);
  nor U12603(n12153,n10776,n8636);
  nor U12604(n12152,n10777,n8554);
  nor U12605(n12151,n10783,n8398);
  nor U12606(n12149,n12155,n12156,n12157,n12158);
  nor U12607(n12158,n10784,n8320);
  nor U12608(n12157,n10785,n8240);
  nor U12609(n12156,n10800,n8082);
  nor U12610(n12155,n10799,n8004);
  nor U12611(n12148,n12159,n12160,n12161,n12162);
  nor U12612(n12162,n10798,n7924);
  nor U12613(n12161,n10792,n7762);
  nor U12614(n12160,n10791,n7682);
  nor U12615(n12159,n10790,n7596);
  nor U12616(n12147,n12163,n12164,n12165,n12166);
  nor U12617(n12166,n10774,n8829);
  nor U12618(n12165,n10782,n8476);
  nor U12619(n12164,n10801,n8160);
  nor U12620(n12163,n10793,n7842);
  nand U12621(n12098,n12167,n12168,n12169,n12170);
  nor U12622(n12170,n12171,n12172,n12173,n12174);
  nor U12623(n12174,n10791,n12050);
  nor U12624(n12173,n10792,n12049);
  nor U12625(n12172,n10793,n12048);
  nand U12626(n12171,n12175,n12176);
  nand U12627(n12176,n12177,G21514);
  nand U12628(n12175,n12178,G21506);
  nor U12629(n12169,n12179,n12180,n12181,n12182);
  nor U12630(n12182,n10801,n12041);
  nor U12631(n12181,n10775,n12040);
  nor U12632(n12180,n10776,n12039);
  nor U12633(n12179,n10777,n12038);
  nor U12634(n12168,n12183,n12184,n12185,n12186);
  nor U12635(n12186,n10783,n12033);
  nor U12636(n12185,n10784,n12032);
  nor U12637(n12184,n10785,n12031);
  nor U12638(n12183,n10790,n12030);
  nor U12639(n12167,n12187,n12188,n12189,n9936);
  nor U12640(n12189,n10774,n12025);
  nor U12641(n12188,n10782,n12024);
  nor U12642(n12187,n10798,n12023);
  not U12643(n12096,n11830);
  nand U12644(n11830,n12190,n12191,n12192,n12193);
  nand U12645(n12193,n11846,n7011);
  nand U12646(n12192,n10249,G21760);
  nand U12647(n12191,G21569,n10250);
  nand U12648(n12190,n9953,n7009);
  nand U12649(n10005,n12194,n11828);
  nand U12650(n11828,n12195,n12196,n12197,n12198);
  nand U12651(n12198,n7001,n11846);
  nand U12652(n12197,n10249,G21761);
  nand U12653(n12196,G21570,n10250);
  nand U12654(n12195,n9953,n6999);
  or U12655(n12194,n11827,n9936);
  nand U12656(n11827,n12199,n12200,n12201,n12202);
  nor U12657(n12202,n12203,n12204);
  nor U12658(n12204,n7465,n8896);
  and U12659(n12203,n11219,n11950);
  nand U12660(n11219,n12205,n12206,n12207,n12208);
  nor U12661(n12208,n12209,n12210,n12211,n12212);
  nor U12662(n12212,n10689,n11959);
  nor U12663(n12211,n10690,n11960);
  nor U12664(n12210,n10691,n11961);
  nor U12665(n12209,n10697,n11962);
  nor U12666(n12207,n12213,n12214,n12215,n12216);
  nor U12667(n12216,n10698,n11967);
  nor U12668(n12215,n10699,n11968);
  nor U12669(n12214,n10714,n11969);
  nor U12670(n12213,n10713,n11970);
  nor U12671(n12206,n12217,n12218,n12219,n12220);
  nor U12672(n12220,n10712,n11975);
  nor U12673(n12219,n10706,n11976);
  nor U12674(n12218,n10705,n11977);
  nor U12675(n12217,n10704,n11978);
  nor U12676(n12205,n12221,n12222,n12223,n12224);
  nor U12677(n12224,n10688,n11983);
  nor U12678(n12223,n10696,n11984);
  nor U12679(n12222,n10715,n11985);
  nor U12680(n12221,n10707,n11986);
  nand U12681(n12201,n10290,n12225);
  nand U12682(n12225,n12226,n12227,n12228,n12229);
  nor U12683(n12229,n12230,n12231,n12232,n12233);
  nor U12684(n12233,n10688,n12234);
  nor U12685(n12232,n10689,n12235);
  nor U12686(n12231,n10690,n12236);
  nor U12687(n12230,n10691,n12237);
  nor U12688(n12228,n12238,n12239,n12240,n12241);
  nor U12689(n12241,n10696,n12242);
  nor U12690(n12240,n10697,n12243);
  nor U12691(n12239,n10698,n12244);
  nor U12692(n12238,n10699,n12245);
  nor U12693(n12227,n12246,n12247,n12248,n12249);
  nor U12694(n12249,n10715,n12250);
  nor U12695(n12248,n10714,n12251);
  nor U12696(n12247,n10713,n12252);
  nor U12697(n12246,n10712,n12253);
  nor U12698(n12226,n12254,n12255,n12256,n12257);
  nor U12699(n12257,n10707,n12258);
  nor U12700(n12256,n10706,n12259);
  nor U12701(n12255,n10705,n12260);
  nor U12702(n12254,n10704,n12261);
  nand U12703(n12200,n12262,n12263,n12264,n12265);
  nor U12704(n12265,n12266,n12267,n12268,n12269);
  nor U12705(n12269,n10705,n12050);
  nor U12706(n12268,n10706,n12049);
  nor U12707(n12267,n10707,n12048);
  nand U12708(n12266,n12270,n12271);
  nand U12709(n12271,n12177,G21513);
  nand U12710(n12270,n12178,G21505);
  nor U12711(n12264,n12272,n12273,n12274,n12275);
  nor U12712(n12275,n10715,n12041);
  nor U12713(n12274,n10689,n12040);
  nor U12714(n12273,n10690,n12039);
  nor U12715(n12272,n10691,n12038);
  nor U12716(n12263,n12276,n12277,n12278,n12279);
  nor U12717(n12279,n10697,n12033);
  nor U12718(n12278,n10698,n12032);
  nor U12719(n12277,n10699,n12031);
  nor U12720(n12276,n10704,n12030);
  nor U12721(n12262,n12280,n12281,n12282,n9936);
  nor U12722(n12282,n10688,n12025);
  nor U12723(n12281,n10696,n12024);
  nor U12724(n12280,n10712,n12023);
  nand U12725(n12199,n11928,n12283);
  nand U12726(n12283,n12284,n12285,n12286,n12287);
  nor U12727(n12287,n12288,n12289,n12290,n12291);
  nor U12728(n12291,n10689,n8714);
  nor U12729(n12290,n10690,n8636);
  nor U12730(n12289,n10691,n8554);
  nor U12731(n12288,n10697,n8398);
  nor U12732(n12286,n12292,n12293,n12294,n12295);
  nor U12733(n12295,n10698,n8320);
  nor U12734(n12294,n10699,n8240);
  nor U12735(n12293,n10714,n8082);
  nor U12736(n12292,n10713,n8004);
  nor U12737(n12285,n12296,n12297,n12298,n12299);
  nor U12738(n12299,n10712,n7924);
  nor U12739(n12298,n10706,n7762);
  nor U12740(n12297,n10705,n7682);
  nor U12741(n12296,n10704,n7596);
  nor U12742(n12284,n12300,n12301,n12302,n12303);
  nor U12743(n12303,n10688,n8829);
  nor U12744(n12302,n10696,n8476);
  nor U12745(n12301,n10715,n8160);
  nor U12746(n12300,n10707,n7842);
  or U12747(n9996,n12304,n12305);
  nand U12748(n9995,n12305,n12304);
  nand U12749(n12304,n12306,n12307,n12308,n12309);
  nand U12750(n12309,n6990,n11846);
  not U12751(n6990,n8873);
  or U12752(n8873,n12310,n12311);
  and U12753(n12311,n12312,n12313);
  nand U12754(n12308,n10249,G21762);
  nand U12755(n12307,G21571,n10250);
  nand U12756(n12306,n9953,n6988);
  or U12757(n12305,n9936,n12314);
  nand U12758(n12314,n12315,n12316,n12317,n12318);
  nor U12759(n12318,n12319,n12320);
  nor U12760(n12320,n7465,n8874);
  nor U12761(n12319,n12321,n9216);
  nor U12762(n12321,n12322,n12323,n12324,n12325);
  nand U12763(n12325,n12326,n12327,n12328,n12329);
  nand U12764(n12329,n11863,G21552);
  not U12765(n11863,n12261);
  nand U12766(n12328,n11864,G21544);
  not U12767(n11864,n12260);
  nand U12768(n12327,n11865,G21536);
  not U12769(n11865,n12259);
  nand U12770(n12326,n11866,G21528);
  not U12771(n11866,n12258);
  nand U12772(n12324,n12330,n12331,n12332,n12333);
  nand U12773(n12333,n11871,G21520);
  not U12774(n11871,n12253);
  nand U12775(n12332,n11872,G21512);
  not U12776(n11872,n12252);
  nand U12777(n12331,n11873,G21504);
  not U12778(n11873,n12251);
  nand U12779(n12330,n11874,G21496);
  not U12780(n11874,n12250);
  nand U12781(n12323,n12334,n12335,n12336,n12337);
  nand U12782(n12337,n11879,G21488);
  not U12783(n11879,n12245);
  nand U12784(n12336,n11880,G21480);
  not U12785(n11880,n12244);
  nand U12786(n12335,n11881,G21472);
  not U12787(n11881,n12243);
  nand U12788(n12334,n11882,G21464);
  not U12789(n11882,n12242);
  nand U12790(n12322,n12338,n12339,n12340,n12341);
  nand U12791(n12341,n11887,G21456);
  not U12792(n11887,n12237);
  nand U12793(n12340,n11888,G21448);
  not U12794(n11888,n12236);
  nand U12795(n12339,n11889,G21440);
  not U12796(n11889,n12235);
  nand U12797(n12338,n11890,G21432);
  not U12798(n11890,n12234);
  nand U12799(n12317,n11950,n11155);
  nand U12800(n11155,n12342,n12343,n12344,n12345);
  nor U12801(n12345,n12346,n12347,n12348,n12349);
  nor U12802(n12349,n10602,n11959);
  nor U12803(n12348,n10603,n11960);
  nor U12804(n12347,n10604,n11961);
  nor U12805(n12346,n10610,n11962);
  nor U12806(n12344,n12350,n12351,n12352,n12353);
  nor U12807(n12353,n10611,n11967);
  nor U12808(n12352,n10612,n11968);
  nor U12809(n12351,n10627,n11969);
  nor U12810(n12350,n10626,n11970);
  nor U12811(n12343,n12354,n12355,n12356,n12357);
  nor U12812(n12357,n10625,n11975);
  nor U12813(n12356,n10619,n11976);
  nor U12814(n12355,n10618,n11977);
  nor U12815(n12354,n10617,n11978);
  nor U12816(n12342,n12358,n12359,n12360,n12361);
  nor U12817(n12361,n10601,n11983);
  nor U12818(n12360,n10609,n11984);
  nor U12819(n12359,n10628,n11985);
  nor U12820(n12358,n10620,n11986);
  nand U12821(n12316,n12362,n12363,n12364,n12365);
  nor U12822(n12365,n12366,n12367,n12368,n12369);
  nor U12823(n12369,n10618,n12050);
  nor U12824(n12368,n10619,n12049);
  nor U12825(n12367,n10620,n12048);
  nand U12826(n12366,n12370,n12371);
  nand U12827(n12371,n12177,G21512);
  nand U12828(n12370,n12178,G21504);
  nor U12829(n12364,n12372,n12373,n12374,n12375);
  nor U12830(n12375,n10628,n12041);
  nor U12831(n12374,n10602,n12040);
  nor U12832(n12373,n10603,n12039);
  nor U12833(n12372,n10604,n12038);
  nor U12834(n12363,n12376,n12377,n12378,n12379);
  nor U12835(n12379,n10610,n12033);
  nor U12836(n12378,n10611,n12032);
  nor U12837(n12377,n10612,n12031);
  nor U12838(n12376,n10617,n12030);
  nor U12839(n12362,n12380,n12381,n12382,n9936);
  nor U12840(n12382,n10601,n12025);
  nor U12841(n12381,n10609,n12024);
  nor U12842(n12380,n10625,n12023);
  nand U12843(n12315,n11928,n12383);
  nand U12844(n12383,n12384,n12385,n12386,n12387);
  nor U12845(n12387,n12388,n12389,n12390,n12391);
  nor U12846(n12391,n10602,n8714);
  nor U12847(n12390,n10603,n8636);
  nor U12848(n12389,n10604,n8554);
  nor U12849(n12388,n10610,n8398);
  nor U12850(n12386,n12392,n12393,n12394,n12395);
  nor U12851(n12395,n10611,n8320);
  nor U12852(n12394,n10612,n8240);
  nor U12853(n12393,n10627,n8082);
  nor U12854(n12392,n10626,n8004);
  nor U12855(n12385,n12396,n12397,n12398,n12399);
  nor U12856(n12399,n10625,n7924);
  nor U12857(n12398,n10619,n7762);
  nor U12858(n12397,n10618,n7682);
  nor U12859(n12396,n10617,n7596);
  nor U12860(n12384,n12400,n12401,n12402,n12403);
  nor U12861(n12403,n10601,n8829);
  nor U12862(n12402,n10609,n8476);
  nor U12863(n12401,n10628,n8160);
  nor U12864(n12400,n10620,n7842);
  or U12865(n9988,n11822,n11821);
  or U12866(n11821,n12404,n9936);
  nand U12867(n12404,n12405,n12406,n12407,n12408);
  nand U12868(n12408,n12409,n12410,n12411,n12412);
  nor U12869(n12412,n12413,n12414,n12415,n12416);
  nor U12870(n12416,n10536,n12050);
  nor U12871(n12415,n10537,n12049);
  nor U12872(n12414,n10538,n12048);
  nand U12873(n12413,n12417,n12418);
  nand U12874(n12418,n12177,G21511);
  nand U12875(n12417,n12178,G21503);
  nor U12876(n12411,n12419,n12420,n12421,n12422);
  nor U12877(n12422,n10546,n12041);
  nor U12878(n12421,n10520,n12040);
  nor U12879(n12420,n10521,n12039);
  nor U12880(n12419,n10522,n12038);
  nor U12881(n12410,n12423,n12424,n12425,n12426);
  nor U12882(n12426,n10528,n12033);
  nor U12883(n12425,n10529,n12032);
  nor U12884(n12424,n10530,n12031);
  nor U12885(n12423,n10535,n12030);
  nor U12886(n12409,n12427,n12428,n12429,n9936);
  nor U12887(n12429,n10519,n12025);
  nor U12888(n12428,n10527,n12024);
  nor U12889(n12427,n10543,n12023);
  nand U12890(n12407,n11950,n11110);
  nand U12891(n11110,n12430,n12431,n12432,n12433);
  nor U12892(n12433,n12434,n12435,n12436,n12437);
  nor U12893(n12437,n10520,n11959);
  nor U12894(n12436,n10521,n11960);
  nor U12895(n12435,n10522,n11961);
  nor U12896(n12434,n10528,n11962);
  nor U12897(n12432,n12438,n12439,n12440,n12441);
  nor U12898(n12441,n10529,n11967);
  nor U12899(n12440,n10530,n11968);
  nor U12900(n12439,n10545,n11969);
  nor U12901(n12438,n10544,n11970);
  nor U12902(n12431,n12442,n12443,n12444,n12445);
  nor U12903(n12445,n10543,n11975);
  nor U12904(n12444,n10537,n11976);
  nor U12905(n12443,n10536,n11977);
  nor U12906(n12442,n10535,n11978);
  nor U12907(n12430,n12446,n12447,n12448,n12449);
  nor U12908(n12449,n10519,n11983);
  nor U12909(n12448,n10527,n11984);
  nor U12910(n12447,n10546,n11985);
  nor U12911(n12446,n10538,n11986);
  nand U12912(n12406,n10290,n12450);
  nand U12913(n12450,n12451,n12452,n12453,n12454);
  nor U12914(n12454,n12455,n12456,n12457,n12458);
  nor U12915(n12458,n10519,n12234);
  nor U12916(n12457,n10520,n12235);
  nor U12917(n12456,n10521,n12236);
  nor U12918(n12455,n10522,n12237);
  nor U12919(n12453,n12459,n12460,n12461,n12462);
  nor U12920(n12462,n10527,n12242);
  nor U12921(n12461,n10528,n12243);
  nor U12922(n12460,n10529,n12244);
  nor U12923(n12459,n10530,n12245);
  nor U12924(n12452,n12463,n12464,n12465,n12466);
  nor U12925(n12466,n10546,n12250);
  nor U12926(n12465,n10545,n12251);
  nor U12927(n12464,n10544,n12252);
  nor U12928(n12463,n10543,n12253);
  nor U12929(n12451,n12467,n12468,n12469,n12470);
  nor U12930(n12470,n10538,n12258);
  nor U12931(n12469,n10537,n12259);
  nor U12932(n12468,n10536,n12260);
  nor U12933(n12467,n10535,n12261);
  nand U12934(n12405,n11928,n12471);
  nand U12935(n12471,n12472,n12473,n12474,n12475);
  nor U12936(n12475,n12476,n12477,n12478,n12479);
  nor U12937(n12479,n10520,n8714);
  nor U12938(n12478,n10521,n8636);
  nor U12939(n12477,n10522,n8554);
  nor U12940(n12476,n10528,n8398);
  nor U12941(n12474,n12480,n12481,n12482,n12483);
  nor U12942(n12483,n10529,n8320);
  nor U12943(n12482,n10530,n8240);
  nor U12944(n12481,n10545,n8082);
  nor U12945(n12480,n10544,n8004);
  nor U12946(n12473,n12484,n12485,n12486,n12487);
  nor U12947(n12487,n10543,n7924);
  nor U12948(n12486,n10537,n7762);
  nor U12949(n12485,n10536,n7682);
  nor U12950(n12484,n10535,n7596);
  nor U12951(n12472,n12488,n12489,n12490,n12491);
  nor U12952(n12491,n10519,n8829);
  nor U12953(n12490,n10527,n8476);
  nor U12954(n12489,n10546,n8160);
  nor U12955(n12488,n10538,n7842);
  nand U12956(n11822,n12492,n12493,n12494,n12495);
  nand U12957(n12495,n6979,n11846);
  not U12958(n6979,n9606);
  or U12959(n9606,n12496,n12497);
  and U12960(n12497,n12498,n12499);
  nand U12961(n12494,n10249,G21763);
  nand U12962(n12493,G21572,n10250);
  nand U12963(n12492,n9953,n6977);
  nand U12964(n9981,n12500,n12501);
  or U12965(n12501,n9953,n11819);
  nand U12966(n11819,n12502,n12503,n12504,n12505);
  nand U12967(n12505,n12506,n12507,n12508,n12509);
  nor U12968(n12509,n12510,n12511,n12512,n12513);
  nor U12969(n12513,n10448,n12050);
  nor U12970(n12512,n10449,n12049);
  nor U12971(n12511,n10450,n12048);
  nand U12972(n12510,n12514,n12515);
  nand U12973(n12515,n12177,G21510);
  nand U12974(n12514,n12178,G21502);
  nor U12975(n12508,n12516,n12517,n12518,n12519);
  nor U12976(n12519,n10458,n12041);
  nor U12977(n12518,n10432,n12040);
  nor U12978(n12517,n10433,n12039);
  nor U12979(n12516,n10434,n12038);
  nor U12980(n12507,n12520,n12521,n12522,n12523);
  nor U12981(n12523,n10440,n12033);
  nor U12982(n12522,n10441,n12032);
  nor U12983(n12521,n10442,n12031);
  nor U12984(n12520,n10447,n12030);
  nor U12985(n12506,n12524,n12525,n12526,n9936);
  nor U12986(n12526,n10431,n12025);
  nor U12987(n12525,n10439,n12024);
  nor U12988(n12524,n10455,n12023);
  nand U12989(n12504,n11950,n10917);
  nand U12990(n10917,n12527,n12528,n12529,n12530);
  nor U12991(n12530,n12531,n12532,n12533,n12534);
  nor U12992(n12534,n10432,n11959);
  nor U12993(n12533,n10433,n11960);
  nor U12994(n12532,n10434,n11961);
  nor U12995(n12531,n10440,n11962);
  nor U12996(n12529,n12535,n12536,n12537,n12538);
  nor U12997(n12538,n10441,n11967);
  nor U12998(n12537,n10442,n11968);
  nor U12999(n12536,n10457,n11969);
  nor U13000(n12535,n10456,n11970);
  nor U13001(n12528,n12539,n12540,n12541,n12542);
  nor U13002(n12542,n10455,n11975);
  nor U13003(n12541,n10449,n11976);
  nor U13004(n12540,n10448,n11977);
  nor U13005(n12539,n10447,n11978);
  nor U13006(n12527,n12543,n12544,n12545,n12546);
  nor U13007(n12546,n10431,n11983);
  nor U13008(n12545,n10439,n11984);
  nor U13009(n12544,n10458,n11985);
  nor U13010(n12543,n10450,n11986);
  nand U13011(n12503,n10290,n12547);
  nand U13012(n12547,n12548,n12549,n12550,n12551);
  nor U13013(n12551,n12552,n12553,n12554,n12555);
  nor U13014(n12555,n10431,n12234);
  nor U13015(n12554,n10432,n12235);
  nor U13016(n12553,n10433,n12236);
  nor U13017(n12552,n10434,n12237);
  nor U13018(n12550,n12556,n12557,n12558,n12559);
  nor U13019(n12559,n10439,n12242);
  nor U13020(n12558,n10440,n12243);
  nor U13021(n12557,n10441,n12244);
  nor U13022(n12556,n10442,n12245);
  nor U13023(n12549,n12560,n12561,n12562,n12563);
  nor U13024(n12563,n10458,n12250);
  nor U13025(n12562,n10457,n12251);
  nor U13026(n12561,n10456,n12252);
  nor U13027(n12560,n10455,n12253);
  nor U13028(n12548,n12564,n12565,n12566,n12567);
  nor U13029(n12567,n10450,n12258);
  nor U13030(n12566,n10449,n12259);
  nor U13031(n12565,n10448,n12260);
  nor U13032(n12564,n10447,n12261);
  nand U13033(n12502,n11928,n12568);
  nand U13034(n12568,n12569,n12570,n12571,n12572);
  nor U13035(n12572,n12573,n12574,n12575,n12576);
  nor U13036(n12576,n10432,n8714);
  nor U13037(n12575,n10433,n8636);
  nor U13038(n12574,n10434,n8554);
  nor U13039(n12573,n10440,n8398);
  nor U13040(n12571,n12577,n12578,n12579,n12580);
  nor U13041(n12580,n10441,n8320);
  nor U13042(n12579,n10442,n8240);
  nor U13043(n12578,n10457,n8082);
  nor U13044(n12577,n10456,n8004);
  nor U13045(n12570,n12581,n12582,n12583,n12584);
  nor U13046(n12584,n10455,n7924);
  nor U13047(n12583,n10449,n7762);
  nor U13048(n12582,n10448,n7682);
  nor U13049(n12581,n10447,n7596);
  nor U13050(n12569,n12585,n12586,n12587,n12588);
  nor U13051(n12588,n10431,n8829);
  nor U13052(n12587,n10439,n8476);
  nor U13053(n12586,n10458,n8160);
  nor U13054(n12585,n10450,n7842);
  not U13055(n12500,n11818);
  nand U13056(n11818,n12589,n12590,n12591,n12592);
  nand U13057(n12592,n6968,n11846);
  not U13058(n6968,n9595);
  nand U13059(n9595,n12593,n12594);
  nand U13060(n12594,n12595,n12596);
  not U13061(n12595,n12597);
  nand U13062(n12593,n12598,n12498,n12599);
  nand U13063(n12598,n12596,n12600);
  nand U13064(n12591,n10249,G21764);
  nand U13065(n12590,G21573,n10250);
  nand U13066(n12589,n9953,n6966);
  nand U13067(n9967,n11816,n11815);
  nand U13068(n11815,n12601,n12602,n12603,n12604);
  nand U13069(n12604,n6957,n11846);
  nand U13070(n11846,n10569,n9216);
  not U13071(n6957,n9586);
  or U13072(n9586,n12605,n12606);
  and U13073(n12606,n12607,n12608);
  nand U13074(n12603,n10249,G21765);
  nand U13075(n12602,G21574,n10250);
  nand U13076(n12601,n9953,n6955);
  or U13077(n11816,n9936,n12609);
  nand U13078(n12609,n12610,n12611,n12612,n12613);
  nand U13079(n12613,n12614,n12615,n12616,n12617);
  nor U13080(n12617,n12618,n12619,n12620,n12621);
  nor U13081(n12621,n10357,n12050);
  nand U13082(n12050,n12622,n12623);
  nor U13083(n12620,n10359,n12049);
  nand U13084(n12049,n12624,n12623);
  nor U13085(n12619,n10361,n12048);
  nand U13086(n12048,n12625,n12623);
  nand U13087(n12618,n12626,n12627);
  nand U13088(n12627,n12177,G21509);
  not U13089(n12177,n11924);
  nand U13090(n11924,n12628,n12622);
  nand U13091(n12626,n12178,G21501);
  not U13092(n12178,n11923);
  nand U13093(n11923,n12628,n12624);
  nor U13094(n12616,n12629,n12630,n12631,n12632);
  nor U13095(n12632,n10373,n12041);
  nand U13096(n12041,n12628,n12625);
  nor U13097(n12631,n10333,n12040);
  nand U13098(n12040,n12633,n12624);
  nor U13099(n12630,n10335,n12039);
  nand U13100(n12039,n12633,n12622);
  nor U13101(n12629,n10337,n12038);
  nand U13102(n12038,n12633,n12634);
  nor U13103(n12615,n12635,n12636,n12637,n12638);
  nor U13104(n12638,n10345,n12033);
  nand U13105(n12033,n12639,n12624);
  nor U13106(n12624,n7033,n9641);
  nor U13107(n12637,n10347,n12032);
  nand U13108(n12032,n12639,n12622);
  nor U13109(n12622,n7022,n7436);
  nor U13110(n12636,n10349,n12031);
  nand U13111(n12031,n12639,n12634);
  nor U13112(n12635,n10355,n12030);
  nand U13113(n12030,n12634,n12623);
  nor U13114(n12623,n7011,n7001);
  nor U13115(n12614,n12640,n12641,n12642,n9936);
  nor U13116(n12642,n10331,n12025);
  nand U13117(n12025,n12633,n12625);
  nor U13118(n12633,n7405,n7413);
  nor U13119(n12641,n10343,n12024);
  nand U13120(n12024,n12639,n12625);
  nor U13121(n12625,n9641,n7436);
  not U13122(n7436,n7033);
  nor U13123(n12639,n7405,n7011);
  nor U13124(n12640,n10367,n12023);
  nand U13125(n12023,n12634,n12628);
  nor U13126(n12628,n7001,n7413);
  not U13127(n7413,n7011);
  nand U13128(n7011,n12643,n12644);
  nand U13129(n12644,n12645,n12646);
  nand U13130(n12645,n12647,n12648);
  nand U13131(n12643,n12649,n12647);
  not U13132(n7001,n7405);
  or U13133(n7405,n12649,n12650);
  and U13134(n12650,n12651,n12652);
  not U13135(n12649,n12653);
  nor U13136(n12634,n7033,n7022);
  not U13137(n7022,n9641);
  or U13138(n9641,n12654,n12655);
  and U13139(n12655,n12656,n12657);
  or U13140(n7033,n12658,n9110);
  nand U13141(n12658,n12659,n12660);
  nand U13142(n12612,n11950,n10920);
  nand U13143(n10920,n12661,n12662,n12663,n12664);
  nor U13144(n12664,n12665,n12666,n12667,n12668);
  nor U13145(n12668,n10333,n11959);
  nand U13146(n11959,n12669,n12670);
  nor U13147(n12667,n10335,n11960);
  nand U13148(n11960,n12671,n12669);
  nor U13149(n12666,n10337,n11961);
  nand U13150(n11961,n12669,n12672);
  nor U13151(n12665,n10345,n11962);
  nand U13152(n11962,n12673,n12670);
  nor U13153(n12663,n12674,n12675,n12676,n12677);
  nor U13154(n12677,n10347,n11967);
  nand U13155(n11967,n12671,n12673);
  nor U13156(n12676,n10349,n11968);
  nand U13157(n11968,n12672,n12673);
  nor U13158(n12675,n10371,n11969);
  nand U13159(n11969,n12678,n12670);
  nor U13160(n12674,n10369,n11970);
  nand U13161(n11970,n12678,n12671);
  nor U13162(n12662,n12679,n12680,n12681,n12682);
  nor U13163(n12682,n10367,n11975);
  nand U13164(n11975,n12678,n12672);
  nor U13165(n12681,n10359,n11976);
  nand U13166(n11976,n12683,n12670);
  nor U13167(n12670,n7031,n12684);
  nor U13168(n12680,n10357,n11977);
  nand U13169(n11977,n12683,n12671);
  nor U13170(n12671,n7447,n7020);
  nor U13171(n12679,n10355,n11978);
  nand U13172(n11978,n12683,n12672);
  nor U13173(n12672,n7031,n7020);
  nor U13174(n12661,n12685,n12686,n12687,n12688);
  nor U13175(n12688,n10331,n11983);
  nand U13176(n11983,n12689,n12669);
  nor U13177(n12669,n7418,n9201);
  nor U13178(n12687,n10343,n11984);
  nand U13179(n11984,n12689,n12673);
  nor U13180(n12673,n9201,n7009);
  nor U13181(n12686,n10373,n11985);
  nand U13182(n11985,n12689,n12678);
  nor U13183(n12678,n7418,n6999);
  nor U13184(n12685,n10361,n11986);
  nand U13185(n11986,n12689,n12683);
  nor U13186(n12683,n6999,n7009);
  nor U13187(n12689,n12684,n7447);
  not U13188(n7447,n7031);
  nand U13189(n12611,n10290,n12690);
  nand U13190(n12690,n12691,n12692,n12693,n12694);
  nor U13191(n12694,n12695,n12696,n12697,n12698);
  nor U13192(n12698,n10331,n12234);
  nand U13193(n12234,n12699,n12700);
  nor U13194(n12697,n10333,n12235);
  nand U13195(n12235,n12699,n12701);
  nor U13196(n12696,n10335,n12236);
  nand U13197(n12236,n12700,n12702);
  nor U13198(n12695,n10337,n12237);
  nand U13199(n12237,n12702,n12701);
  nor U13200(n12693,n12703,n12704,n12705,n12706);
  nor U13201(n12706,n10343,n12242);
  nand U13202(n12242,n12707,n12700);
  nor U13203(n12705,n10345,n12243);
  nand U13204(n12243,n12707,n12701);
  nor U13205(n12704,n10347,n12244);
  nand U13206(n12244,n12708,n12700);
  nor U13207(n12700,n12709,G21561);
  nor U13208(n12703,n10349,n12245);
  nand U13209(n12245,n12708,n12701);
  nor U13210(n12701,n12709,n8916);
  not U13211(n12709,n9220);
  nor U13212(n12692,n12710,n12711,n12712,n12713);
  nor U13213(n12713,n10373,n12250);
  nand U13214(n12250,n12714,n12699);
  nor U13215(n12712,n10371,n12251);
  nand U13216(n12251,n12715,n12699);
  and U13217(n12699,n9182,n9164);
  nor U13218(n12711,n10369,n12252);
  nand U13219(n12252,n12714,n12702);
  nor U13220(n12710,n10367,n12253);
  nand U13221(n12253,n12715,n12702);
  and U13222(n12702,n12716,n9182);
  nor U13223(n12691,n12717,n12718,n12719,n12720);
  nor U13224(n12720,n10361,n12258);
  nand U13225(n12258,n12714,n12707);
  nor U13226(n12719,n10359,n12259);
  nand U13227(n12259,n12715,n12707);
  nor U13228(n12707,n9182,n12716);
  nor U13229(n12718,n10357,n12260);
  nand U13230(n12260,n12714,n12708);
  nor U13231(n12714,n9220,G21561);
  nor U13232(n12717,n10355,n12261);
  nand U13233(n12261,n12715,n12708);
  nor U13234(n12708,n9182,n9164);
  not U13235(n9164,n12716);
  nor U13236(n12716,n9160,n10989);
  nand U13237(n9182,n12721,n12722);
  nand U13238(n12722,n12723,n12724);
  nand U13239(n12724,n9101,n8919);
  nand U13240(n12721,n10997,n12725);
  nor U13241(n12715,n8916,n9220);
  or U13242(n9220,n12723,n8896);
  and U13243(n12723,n12726,n12725);
  nand U13244(n12725,n12727,n10997);
  or U13245(n12727,n9101,G21559);
  nand U13246(n12726,G21559,n8737);
  nand U13247(n12610,n11928,n12728);
  nand U13248(n9958,n12729,n12730,n12731,n12732);
  nor U13249(n12732,n12733,n12734);
  and U13250(n12734,n6944,n9953);
  nor U13251(n12733,n10569,n9577);
  nand U13252(n12731,G21575,n10250);
  or U13253(n12735,n12737,n6946);
  nand U13254(n12729,n10249,G21766);
  not U13255(n9952,n9950);
  nand U13256(n9950,n12738,n12739,n12740,n12741);
  nor U13257(n12741,n12742,n12743);
  nor U13258(n12743,n7340,n9936);
  nor U13259(n12742,n10569,n7336);
  nand U13260(n12740,G21576,n10250);
  or U13261(n12744,n12745,n7336);
  or U13262(n12745,n12746,n12747);
  nand U13263(n12738,n10249,G21767);
  nand U13264(n9939,n12748,n12749,n12750,n12751);
  nor U13265(n12751,n12752,n12753);
  nor U13266(n12753,n7325,n9936);
  not U13267(n7325,n6913);
  nor U13268(n12752,n10569,n6916);
  nand U13269(n12750,G21577,n10250);
  or U13270(n12754,n12755,n12756);
  or U13271(n12756,n12757,n6916);
  nand U13272(n12748,n10249,G21768);
  nand U13273(n11742,n12758,n12759,n12760,n12761);
  nor U13274(n12761,n12762,n12763);
  and U13275(n12763,n9953,n7317);
  nor U13276(n12762,n10569,n9550);
  nor U13277(n10569,n11928,n11950);
  nor U13278(n11950,n9117,n7477,n12765);
  nand U13279(n12760,G21578,n10250);
  not U13280(n10250,n10285);
  nor U13281(n10285,n9219,n9217,n11851);
  or U13282(n12766,n11756,n12767);
  or U13283(n12767,n11754,n9550);
  nand U13284(n9550,n11758,n12768);
  nand U13285(n12768,n12769,n12770);
  or U13286(n11758,n12770,n12769);
  or U13287(n12769,n12771,n9110);
  nand U13288(n12771,n12772,n12773,n12774,n12775);
  nand U13289(n12775,G21578,n10247);
  nand U13290(n12774,n7317,n10305);
  nand U13291(n12773,G21610,n11083);
  nand U13292(n12772,G21769,n9284);
  nand U13293(n11756,n12776,n12777);
  nand U13294(n12777,n12757,n12778);
  or U13295(n12778,n12755,n6916);
  not U13296(n12757,n12779);
  nand U13297(n12776,n12755,n6916);
  nand U13298(n6916,n12780,n12770);
  or U13299(n12770,n12781,n12782);
  nand U13300(n12780,n12782,n12781);
  or U13301(n12782,n12783,n9110);
  nand U13302(n12783,n12784,n12785,n12786,n12787);
  nand U13303(n12787,n6913,n10305);
  nand U13304(n6913,n12788,n12789);
  nand U13305(n12789,n12790,n12791);
  nand U13306(n12791,n12792,n12793);
  not U13307(n12792,n12794);
  nand U13308(n12788,n12795,n12796);
  nand U13309(n12786,G21577,n10247);
  nand U13310(n12785,G21609,n11083);
  nand U13311(n12784,G21768,n9284);
  nand U13312(n12755,n12797,n12798);
  nand U13313(n12798,n12746,n12799);
  nand U13314(n12799,n12747,n6934);
  not U13315(n6934,n7336);
  not U13316(n12747,n12736);
  not U13317(n12746,n12800);
  nand U13318(n12797,n7336,n12736);
  nand U13319(n12736,n6946,n12737);
  not U13320(n6946,n9577);
  nand U13321(n9577,n12801,n12802);
  or U13322(n12801,n12803,n12804);
  nand U13323(n7336,n12781,n12805);
  nand U13324(n12805,n12806,n12802);
  or U13325(n12781,n12802,n12806);
  or U13326(n12806,n12807,n9110);
  nand U13327(n12807,n12808,n12809,n12810,n12811);
  nand U13328(n12811,n6930,n10305);
  not U13329(n6930,n7340);
  or U13330(n7340,n12812,n12813);
  nand U13331(n12812,n12814,n12815);
  nand U13332(n12810,G21576,n10247);
  nand U13333(n12809,G21608,n11083);
  nand U13334(n12808,G21767,n9284);
  nand U13335(n12802,n12804,n12803);
  nand U13336(n12803,n12816,n12607);
  nand U13337(n12607,n9783,G21549,n12817);
  or U13338(n12817,n12818,n9110);
  nand U13339(n12816,n12608,n12605);
  nand U13340(n12605,n12597,n12596);
  nand U13341(n12596,n9783,G21550,n12819);
  or U13342(n12819,n12820,n9110);
  nand U13343(n12597,n12600,n12821);
  nand U13344(n12821,n12599,n12498);
  nand U13345(n12498,n9783,G21551,n12822);
  or U13346(n12822,n12823,n9110);
  nand U13347(n12599,n12499,n12496);
  nand U13348(n12496,n12312,n12824);
  nand U13349(n12824,n12313,n12310);
  nand U13350(n12310,n12651,n12825);
  nand U13351(n12825,n12653,n12652);
  nand U13352(n12652,n12826,n12827);
  nand U13353(n12827,n9783,G21553);
  or U13354(n12826,n7590,n12828);
  nand U13355(n12653,n12648,n12829);
  nand U13356(n12829,n12646,n12647);
  nand U13357(n12647,n12830,n12831,n12832,n8830);
  or U13358(n12830,n7590,n12833);
  nand U13359(n12646,n12656,n12834);
  nand U13360(n12834,n12654,n12657);
  or U13361(n12657,n12835,n12836);
  nand U13362(n12654,n12660,n12837);
  nand U13363(n12837,n7590,n12659);
  nand U13364(n12659,n12838,n12839);
  or U13365(n12839,n7590,n12840);
  not U13366(n12838,n12841);
  nand U13367(n12660,n12842,n12841);
  nand U13368(n12841,n12843,n12844,n12832,n8809);
  nand U13369(n12844,G21428,n12845);
  nand U13370(n12845,n12846,n12847,n12848,n12849);
  nor U13371(n12849,n9210,n12850,n12851,n12852);
  nor U13372(n12852,n9779,n9218);
  nor U13373(n12851,n12765,n9302);
  nor U13374(n12848,n12853,n12854);
  nand U13375(n12847,n9779,n7468);
  nand U13376(n12846,n12855,n8798);
  nand U13377(n12843,n9783,G21556);
  or U13378(n12842,n12840,n9110);
  nand U13379(n12840,n12856,n12857,n12858,n12859);
  nor U13380(n12859,n12860,n12861);
  nor U13381(n12861,n10248,n7030);
  not U13382(n7030,G21758);
  nor U13383(n12860,n10246,n7029);
  nand U13384(n12858,G21567,n10247);
  nand U13385(n12857,n7031,n10305);
  or U13386(n7031,n12862,n10248);
  nand U13387(n12862,n12863,n12864);
  nand U13388(n12856,G21561,n12865);
  nand U13389(n12656,n12836,n12835);
  nand U13390(n12835,n10248,n8855,n12866,n12867);
  nor U13391(n12867,n12868,n12869,n12870);
  nor U13392(n12870,n10879,n9290);
  nor U13393(n12869,n7477,n12871);
  not U13394(n12868,n12872);
  nand U13395(n12866,n11992,n9305,n12873,G21428);
  or U13396(n12836,n9110,n12874);
  nand U13397(n12874,n12875,n12876,n12877,n12878);
  nor U13398(n12878,n12879,n12880);
  nor U13399(n12880,n10248,n7019);
  not U13400(n7019,G21759);
  nor U13401(n12879,n10246,n7018);
  nand U13402(n12877,G21568,n10247);
  nand U13403(n12876,n7020,n10305);
  not U13404(n7020,n12684);
  or U13405(n12684,n12881,n12882);
  and U13406(n12882,n12883,n12884);
  nand U13407(n12875,G21560,n12865);
  nand U13408(n12648,n12885,n12886);
  nand U13409(n12886,n12832,n8830,n12831);
  nand U13410(n12831,n9783,G21554);
  or U13411(n12885,n12833,n9110);
  nand U13412(n12833,n12887,n12888,n12889,n12890);
  nand U13413(n12890,G21569,n10247);
  nor U13414(n12889,n12891,n12892);
  and U13415(n12892,n12865,G21559);
  and U13416(n12891,n10305,n7009);
  not U13417(n7009,n7418);
  nand U13418(n7418,n12893,n12894);
  nand U13419(n12894,n12895,n12883,n12896);
  or U13420(n12896,n9284,n12897);
  nand U13421(n12888,G21601,n11083);
  nand U13422(n12887,G21760,n9284);
  nand U13423(n12651,n9783,G21553,n12898);
  or U13424(n12898,n12828,n9110);
  nand U13425(n12828,n12899,n12900,n12901,n12902);
  nor U13426(n12902,n12903,n12904);
  nor U13427(n12904,n10248,n6998);
  not U13428(n6998,G21761);
  nor U13429(n12903,n10246,n6997);
  nand U13430(n12901,G21570,n10247);
  nand U13431(n12900,G21558,n12865);
  nand U13432(n12865,n12905,n12906,n8809,n10039);
  not U13433(n10039,n10264);
  nand U13434(n12905,G21428,n12907);
  nand U13435(n12907,n7449,n12908);
  nand U13436(n12908,n12855,n8887);
  not U13437(n12855,n12764);
  nand U13438(n12764,n9117,n7470);
  and U13439(n7449,n9221,n9240,n12909);
  nand U13440(n9221,n12910,n9101);
  nand U13441(n12899,n6999,n10305);
  not U13442(n6999,n9201);
  nand U13443(n9201,n12911,n12912);
  nand U13444(n12912,n12913,n12893);
  nand U13445(n12313,n12914,n12915);
  nand U13446(n12915,n9783,G21552);
  or U13447(n12914,n7590,n12916);
  nand U13448(n12312,n9783,G21552,n12917);
  or U13449(n12917,n12916,n9110);
  nand U13450(n12916,n12918,n12919,n12920,n12921);
  nor U13451(n12921,n12922,n12923);
  nor U13452(n12923,n10248,n6987);
  not U13453(n6987,G21762);
  nor U13454(n12922,n10246,n6986);
  not U13455(n6986,G21603);
  nand U13456(n12920,G21571,n10247);
  nand U13457(n12919,G21557,n12924);
  nand U13458(n12924,n12906,n12925);
  nand U13459(n12925,n9200,G21428);
  not U13460(n9200,n9240);
  nand U13461(n9240,n9671,n9210);
  not U13462(n9671,n8884);
  nand U13463(n12918,n6988,n10305);
  and U13464(n6988,n12926,n12927);
  nand U13465(n12927,n12928,n12911);
  nand U13466(n12499,n12929,n12930);
  nand U13467(n12930,n9783,G21551);
  or U13468(n12929,n7590,n12823);
  nand U13469(n12823,n12931,n12932,n12933,n12934);
  nand U13470(n12934,n6977,n10305);
  and U13471(n6977,n12935,n12936);
  nand U13472(n12936,n12937,n12926);
  nand U13473(n12933,G21572,n10247);
  nand U13474(n12932,G21604,n11083);
  nand U13475(n12931,G21763,n9284);
  nand U13476(n12600,n12938,n12939);
  nand U13477(n12939,n9783,G21550);
  or U13478(n12938,n7590,n12820);
  nand U13479(n12820,n12940,n12941,n12942,n12943);
  nand U13480(n12943,n6966,n10305);
  and U13481(n6966,n12944,n12945);
  nand U13482(n12945,n12946,n12935);
  nand U13483(n12942,G21573,n10247);
  nand U13484(n12941,G21605,n11083);
  nand U13485(n12940,G21764,n9284);
  nand U13486(n12608,n12947,n12948);
  nand U13487(n12948,n9783,G21549);
  or U13488(n12947,n7590,n12818);
  nand U13489(n12818,n12949,n12950,n12951,n12952);
  nand U13490(n12952,n6955,n10305);
  nor U13491(n6955,n12953,n12954);
  and U13492(n12954,n12955,n12944);
  nand U13493(n12951,G21574,n10247);
  nand U13494(n12950,G21606,n11083);
  nand U13495(n12949,G21765,n9284);
  or U13496(n12804,n12956,n7590);
  nand U13497(n12956,n12957,n12958,n12959,n12960);
  nand U13498(n12960,n6944,n10305);
  or U13499(n6944,n12953,n12961);
  and U13500(n12961,n12962,n12963);
  nand U13501(n12959,G21575,n10247);
  nand U13502(n12832,G21428,n8798,n7472,n12966);
  and U13503(n12966,n12873,n11928);
  nor U13504(n11928,n12967,n9101);
  nand U13505(n12965,G21428,n7443);
  nand U13506(n7443,n9197,n12968);
  and U13507(n9197,n12969,n12970);
  nand U13508(n12970,n12850,n12971);
  nand U13509(n12969,n12910,n8737);
  not U13510(n12910,n12972);
  nand U13511(n12958,G21607,n11083);
  nand U13512(n12957,G21766,n9284);
  nand U13513(n12758,G21769,n10249);
  not U13514(n10249,n10287);
  nand U13515(n10287,n11992,n7477);
  and U13516(n11992,n10143,n8737,n7481);
  nand U13517(n11797,n7317,n6912);
  nand U13518(n12973,n9085,n8843,n8923);
  or U13519(n9293,n9281,n9282);
  nand U13520(n9282,n8887,G21426,n9672);
  not U13521(n9281,n7467);
  nor U13522(n7467,n12974,n12975);
  and U13523(n12975,n12976,n12977,n12978,n12979);
  nand U13524(n12979,n12980,n12981,n12982);
  or U13525(n12982,n12983,n7470);
  nand U13526(n12981,n12984,n12985,n12986);
  not U13527(n12986,n12987);
  nand U13528(n12984,n9087,n12988);
  or U13529(n12980,n12988,n9087);
  nand U13530(n12978,n12983,n7470);
  nand U13531(n12977,n12989,n12990);
  or U13532(n7317,n12795,n12991);
  and U13533(n12991,n11793,n11795);
  nand U13534(n11795,n12992,n12993);
  nand U13535(n12993,n9783,n12994);
  or U13536(n11793,n9290,n11754,n12992);
  or U13537(n12992,n12995,n10248);
  nand U13538(n12995,n12996,n12997,n12998,n12999);
  nand U13539(n12999,G21705,n10264);
  nand U13540(n12998,G21737,n10316);
  nand U13541(n12997,G21578,n10504);
  nand U13542(n12996,G21610,n7590);
  not U13543(n11754,n12994);
  nand U13544(n12994,n13000,n13001,n13002,n13003);
  nor U13545(n13003,n13004,n13005,n13006,n13007);
  nor U13546(n13007,n10713,n11579);
  nor U13547(n13006,n10712,n11589);
  nor U13548(n13005,n10704,n11588);
  nor U13549(n13004,n10696,n11587);
  nor U13550(n13002,n13008,n13009,n13010,n13011);
  nor U13551(n13011,n10705,n11572);
  nor U13552(n13010,n10699,n11571);
  nor U13553(n13009,n10715,n11581);
  nor U13554(n13008,n10714,n11580);
  nor U13555(n13001,n13012,n13013,n13014,n13015);
  nor U13556(n13015,n10697,n11565);
  nor U13557(n13014,n10691,n11564);
  nor U13558(n13013,n10690,n11563);
  nor U13559(n13012,n10706,n11573);
  nor U13560(n13000,n13016,n13017,n13018,n13019);
  nor U13561(n13019,n10688,n11586);
  nor U13562(n13018,n10689,n11562);
  nor U13563(n13017,n10698,n11570);
  nor U13564(n13016,n10707,n11578);
  not U13565(n9290,n9783);
  not U13566(n12795,n11796);
  nand U13567(n11796,n12793,n12794);
  nand U13568(n12794,n12796,n12790);
  nand U13569(n12790,n12815,n13020);
  nand U13570(n13020,n12814,n12813);
  nand U13571(n12813,n12962,n13021);
  nand U13572(n13021,n12953,n12963);
  nand U13573(n12963,n13022,n13023);
  nand U13574(n13023,n9783,n12737);
  or U13575(n13022,n9284,n13024);
  nor U13576(n12953,n12944,n12955);
  or U13577(n12955,n13025,n10248);
  nand U13578(n13025,n13026,n13027,n13028,n13029);
  nand U13579(n13029,G21701,n10264);
  nand U13580(n13028,G21733,n10316);
  nand U13581(n13027,G21574,n10504);
  nand U13582(n13026,G21606,n7590);
  or U13583(n12944,n12935,n12946);
  or U13584(n12946,n13030,n10248);
  nand U13585(n13030,n13031,n13032,n13033,n13034);
  nand U13586(n13034,G21700,n10264);
  nand U13587(n13033,G21732,n10316);
  nand U13588(n13032,G21573,n10504);
  nand U13589(n13031,G21605,n7590);
  or U13590(n12935,n12926,n12937);
  or U13591(n12937,n13035,n10248);
  nand U13592(n13035,n13036,n13037,n13038,n13039);
  nand U13593(n13039,G21699,n10264);
  nand U13594(n13038,G21731,n10316);
  nand U13595(n13037,G21572,n10504);
  nand U13596(n13036,G21604,n7590);
  or U13597(n12926,n12911,n12928);
  or U13598(n12928,n13040,n10248);
  nand U13599(n13040,n13041,n13042,n13043,n13044);
  nand U13600(n13044,G21698,n10264);
  nand U13601(n13043,G21730,n10316);
  nand U13602(n13042,G21571,n10504);
  nand U13603(n13041,G21603,n7590);
  or U13604(n12911,n12893,n12913);
  or U13605(n12913,n13045,n10248);
  nand U13606(n13045,n13046,n13047,n13048,n13049);
  nor U13607(n13049,n13050,n13051,n13052,n13053);
  and U13608(n13053,n10264,G21697);
  nor U13609(n13052,n13054,n8896);
  nor U13610(n13051,n8825,n8809);
  nor U13611(n13050,n8830,n9198);
  or U13612(n9198,n13055,n13056);
  nor U13613(n13056,n7499,n13057);
  and U13614(n13057,n13058,G21558);
  nor U13615(n7499,n9196,G21426);
  nand U13616(n13055,n13059,n13060);
  nand U13617(n13060,n13061,n13062);
  or U13618(n13061,n13063,n13064);
  nand U13619(n13059,n13063,n13064);
  nor U13620(n13048,n13065,n13066);
  nor U13621(n13066,n9110,n6997);
  not U13622(n6997,G21602);
  nor U13623(n13065,n8855,n9196);
  nand U13624(n13047,G21729,n10316);
  nand U13625(n13046,G21570,n10504);
  nand U13626(n12893,n13067,n13068);
  nand U13627(n13068,n12895,n12883);
  nand U13628(n12883,n13069,n13070);
  nand U13629(n12895,n12884,n12881);
  nand U13630(n12881,n12864,n13071);
  nand U13631(n13071,n9284,n12863);
  nand U13632(n12863,n13072,n13073);
  or U13633(n13073,n9284,n13074);
  not U13634(n13072,n13075);
  nand U13635(n12864,n13076,n13075);
  nand U13636(n13075,n10246,n13077,n8809,n9291);
  nand U13637(n13077,G21428,n13078);
  nand U13638(n13078,n9243,n13079,n13080,n13081);
  nor U13639(n13081,n13082,n13083,n13084);
  nor U13640(n13084,n9779,n13085);
  nor U13641(n13083,n7472,n13086,n13087);
  nor U13642(n13087,n7481,n9779);
  nor U13643(n13082,n12765,n7482);
  not U13644(n13080,n12854);
  nand U13645(n12854,n13088,n13089,n13090);
  nand U13646(n13090,n7481,n7482);
  nand U13647(n13088,n9305,n9101);
  nand U13648(n13079,n12850,n7477);
  and U13649(n9243,n13091,n13092);
  nand U13650(n13092,n9248,n7470);
  not U13651(n10246,n11083);
  nand U13652(n11083,n8830,n8855);
  or U13653(n13076,n13074,n10248);
  nand U13654(n13074,n13093,n13094,n13095,n13096);
  nor U13655(n13096,n13097,n13098,n13099,n13100);
  and U13656(n13100,n10264,G21694);
  nor U13657(n13099,n13054,n8916);
  nor U13658(n13098,n8566,n8809);
  nor U13659(n13097,n8830,n9135);
  nand U13660(n9135,n13101,n13102);
  nand U13661(n13102,n9673,n13103);
  nor U13662(n13095,n13104,n13105);
  nor U13663(n13105,n9110,n7029);
  not U13664(n7029,G21599);
  nor U13665(n13104,n8855,n9137);
  nand U13666(n13094,G21726,n10316);
  nand U13667(n13093,G21567,n10504);
  or U13668(n12884,n13070,n13069);
  or U13669(n13069,n13106,n10248);
  nand U13670(n13106,n13107,n13108,n13109,n13110);
  nor U13671(n13110,n13111,n13112,n13113,n13114);
  and U13672(n13114,n10264,G21695);
  nor U13673(n13113,n13054,n10990);
  nor U13674(n13112,n8906,n8809);
  nor U13675(n13111,n9157,n8830);
  or U13676(n9157,n13115,n13101);
  or U13677(n13115,n13116,n13117);
  nor U13678(n13109,n13118,n13119);
  nor U13679(n13119,n9110,n7018);
  not U13680(n7018,G21600);
  nor U13681(n13118,n9162,n8855);
  nand U13682(n13108,G21727,n10316);
  nand U13683(n13107,G21568,n10504);
  nand U13684(n13070,n12872,n13120,n13121,n13122);
  nor U13685(n13121,n7590,n10041);
  nor U13686(n12872,n10040,n13123);
  nor U13687(n13123,n8843,n7468,n9224);
  or U13688(n13067,n12897,n10248);
  nand U13689(n12897,n13124,n13125,n13126,n13127);
  nor U13690(n13127,n13128,n13129,n13130,n13131);
  and U13691(n13131,n10264,G21696);
  nor U13692(n13130,n13054,n8919);
  and U13693(n13054,n9291,n12871,n12964);
  and U13694(n12964,n13122,n13132);
  nand U13695(n13132,G21428,n13133);
  nand U13696(n13133,n9205,n13134,n13135,n13136);
  nor U13697(n13136,n7444,n13137,n13138,n13139);
  nor U13698(n13139,n9102,n9307);
  nor U13699(n9102,n9210,n13140);
  nor U13700(n13140,n7470,n9101);
  nor U13701(n13138,n13141,n9302);
  not U13702(n9302,n9248);
  nor U13703(n9248,n8737,n7482);
  nor U13704(n13141,n13142,n9305);
  nor U13705(n13142,n7468,n12967);
  nor U13706(n13137,n9218,n9101,n12850);
  not U13707(n9218,n13086);
  nor U13708(n7444,n9224,n7484);
  nor U13709(n13135,n13143,n13144);
  nor U13710(n13144,n7481,n13089);
  not U13711(n13089,n9209);
  and U13712(n13143,n13145,n9657);
  or U13713(n13134,n9216,n9204);
  and U13714(n9205,n13146,n13147,n13148,n13149);
  nand U13715(n13149,n12850,n13150);
  nand U13716(n13150,n7472,n12967,n9779);
  nand U13717(n13148,n7468,n7482,n8808);
  nand U13718(n13147,n13086,n9307);
  not U13719(n13146,n12853);
  nand U13720(n12853,n13151,n13091,n13152);
  nand U13721(n13152,n13153,n8788);
  nand U13722(n13153,n9242,n9247);
  nand U13723(n13091,n11851,n7477);
  nand U13724(n13151,n13154,n8769);
  nand U13725(n13154,n7465,n13155);
  nand U13726(n13155,n7481,n7484);
  nand U13727(n13122,G21428,n10143,n8882);
  not U13728(n8882,n9211);
  nand U13729(n9211,n7481,n8737,n7472,n13156);
  nor U13730(n13156,n13157,n9658);
  nand U13731(n12871,G21428,n7483,n8887);
  not U13732(n9291,n10041);
  nor U13733(n10041,n9159,n8843);
  nand U13734(n9159,n10290,n13085,n9087,n7484);
  nor U13735(n13085,n7482,n12850,n8798);
  nor U13736(n10290,n8737,n9779);
  nor U13737(n13129,n9180,n8830);
  nand U13738(n8830,G21797,G21427);
  not U13739(n9180,n11508);
  or U13740(n11508,n13063,n13158);
  or U13741(n13158,n13062,n13064);
  nor U13742(n13064,n13159,n7495);
  nor U13743(n7495,n9179,G21426);
  and U13744(n13159,G21559,n13058);
  and U13745(n13063,n13160,n13161);
  nand U13746(n13161,n13117,n13162);
  nand U13747(n13162,n13116,n13101);
  not U13748(n13117,n13163);
  or U13749(n13160,n13101,n13116);
  nor U13750(n13116,n13164,n7490);
  nor U13751(n7490,n9162,G21426);
  and U13752(n13164,G21560,n13058);
  nand U13753(n13101,n9078,n13165);
  nand U13754(n13165,n13166,n13103);
  nand U13755(n13103,G21561,n13058);
  nand U13756(n13058,n13163,n13062,n13167);
  nand U13757(n13167,n9209,G21426);
  nor U13758(n9209,n8769,n9101);
  not U13759(n13062,n9667);
  nor U13760(n9667,n7470,n7456);
  nand U13761(n13163,G21426,n13168);
  nand U13762(n13168,n13169,n13145);
  nand U13763(n13169,n9210,n10143);
  nand U13764(n13166,n9109,n7456);
  not U13765(n9078,n9673);
  nor U13766(n9673,n8737,n7456);
  nor U13767(n13128,n8826,n8809);
  not U13768(n8809,n8824);
  nor U13769(n8824,G21426,G21427);
  nor U13770(n13126,n13170,n13171);
  nor U13771(n13171,n9110,n7008);
  not U13772(n7008,G21601);
  nor U13773(n13170,n8855,n9179);
  nand U13774(n13125,G21728,n10316);
  nand U13775(n13124,G21569,n10504);
  nand U13776(n12962,n13024,n12737,n9783);
  nand U13777(n12737,n13172,n13173,n13174,n13175);
  nor U13778(n13175,n13176,n13177,n13178,n13179);
  nor U13779(n13179,n10985,n11579);
  nor U13780(n13178,n10984,n11589);
  nor U13781(n13177,n10972,n11588);
  nor U13782(n13176,n10961,n11587);
  nor U13783(n13174,n13180,n13181,n13182,n13183);
  nor U13784(n13183,n10974,n11572);
  nor U13785(n13182,n10967,n11571);
  nor U13786(n13181,n10987,n11581);
  nor U13787(n13180,n10986,n11580);
  nor U13788(n13173,n13184,n13185,n13186,n13187);
  nor U13789(n13187,n10963,n11565);
  nor U13790(n13186,n10956,n11564);
  nor U13791(n13185,n10954,n11563);
  nor U13792(n13184,n10976,n11573);
  nor U13793(n13172,n13188,n13189,n13190,n13191);
  nor U13794(n13191,n10949,n11586);
  nor U13795(n13190,n10952,n11562);
  nor U13796(n13189,n10964,n11570);
  nor U13797(n13188,n10977,n11578);
  nand U13798(n13024,n13192,n13193,n13194,n13195);
  nand U13799(n13195,G21702,n10264);
  nand U13800(n13194,G21734,n10316);
  nand U13801(n13193,G21575,n10504);
  nand U13802(n13192,G21607,n7590);
  nand U13803(n12814,n13196,n13197);
  nand U13804(n13197,n9783,n12800);
  or U13805(n13196,n9284,n13198);
  nand U13806(n12815,n12800,n13198,n9783);
  nand U13807(n13198,n13199,n13200,n13201,n13202);
  nand U13808(n13202,G21703,n10264);
  nand U13809(n13201,G21735,n10316);
  nand U13810(n13200,G21576,n10504);
  nand U13811(n13199,G21608,n7590);
  nand U13812(n12800,n13203,n13204,n13205,n13206);
  nor U13813(n13206,n13207,n13208,n13209,n13210);
  nor U13814(n13210,n10864,n11562);
  nor U13815(n13209,n10865,n11563);
  nor U13816(n13208,n10866,n11564);
  nor U13817(n13207,n10872,n11565);
  nor U13818(n13205,n13211,n13212,n13213,n13214);
  nor U13819(n13214,n10873,n11570);
  nor U13820(n13213,n10874,n11571);
  nor U13821(n13212,n10880,n11572);
  nor U13822(n13211,n10881,n11573);
  nor U13823(n13204,n13215,n13216,n13217,n13218);
  nor U13824(n13218,n10882,n11578);
  nor U13825(n13217,n10888,n11579);
  nor U13826(n13216,n10889,n11580);
  nor U13827(n13215,n10890,n11581);
  nor U13828(n13203,n13219,n13220,n13221,n13222);
  nor U13829(n13222,n10863,n11586);
  nor U13830(n13221,n10871,n11587);
  nor U13831(n13220,n10879,n11588);
  nor U13832(n13219,n10887,n11589);
  nand U13833(n12796,n13223,n13224);
  nand U13834(n13224,n9783,n12779);
  or U13835(n13223,n9284,n13225);
  nand U13836(n12793,n13225,n12779,n9783);
  not U13837(n7454,n9163);
  nor U13838(n9163,n13226,n12099,n13157,n7481);
  not U13839(n12099,n11851);
  nor U13840(n11851,n7472,n9101);
  nand U13841(n12779,n13227,n13228,n13229,n13230);
  nor U13842(n13230,n13231,n13232,n13233,n13234);
  nor U13843(n13234,n10799,n11579);
  nand U13844(n11579,n13235,n10997);
  nor U13845(n13233,n10798,n11589);
  nand U13846(n11589,n13235,n10989);
  nor U13847(n13232,n10790,n11588);
  nand U13848(n11588,n13236,n10989);
  nor U13849(n13231,n10782,n11587);
  nand U13850(n11587,n13237,n9160);
  nor U13851(n13229,n13238,n13239,n13240,n13241);
  nor U13852(n13241,n10791,n11572);
  nand U13853(n11572,n13236,n10997);
  nor U13854(n13240,n10785,n11571);
  nand U13855(n11571,n13237,n10989);
  nor U13856(n13239,n10801,n11581);
  nand U13857(n11581,n13235,n9160);
  nor U13858(n13238,n10800,n11580);
  nand U13859(n11580,n13235,n8915);
  nor U13860(n13235,n13242,n13243);
  nor U13861(n13228,n13244,n13245,n13246,n13247);
  nor U13862(n13247,n10783,n11565);
  nand U13863(n11565,n13237,n8915);
  nor U13864(n13246,n10777,n11564);
  nand U13865(n11564,n13248,n10989);
  nor U13866(n13245,n10776,n11563);
  nand U13867(n11563,n13248,n10997);
  nor U13868(n13244,n10792,n11573);
  nand U13869(n11573,n13236,n8915);
  nor U13870(n13227,n13249,n13250,n13251,n13252);
  nor U13871(n13252,n10774,n11586);
  nand U13872(n11586,n13248,n9160);
  nor U13873(n13251,n10775,n11562);
  nand U13874(n11562,n13248,n8915);
  and U13875(n13248,n13253,n13242);
  nor U13876(n13250,n10784,n11570);
  nand U13877(n11570,n13237,n10997);
  and U13878(n13237,n13243,n13242);
  not U13879(n13243,n13253);
  nor U13880(n13249,n10793,n11578);
  nand U13881(n11578,n13236,n9160);
  nor U13882(n13236,n13242,n13253);
  or U13883(n13253,G21560,n8919);
  nand U13884(n13242,n13254,n13255,n13256);
  not U13885(n13256,n13257);
  nand U13886(n13255,G21558,n10990);
  nand U13887(n13254,n13258,G21560);
  nand U13888(n13225,n13259,n13260,n13261,n13262);
  nand U13889(n13262,G21704,n10264);
  nor U13890(n10264,n7452,n8843);
  nand U13891(n7452,n13263,n13086,n9101,n7477);
  nor U13892(n13086,n7468,n8788);
  nand U13893(n13261,G21736,n10316);
  nand U13894(n10316,n10248,n9781);
  nand U13895(n9781,n9199,G21428);
  not U13896(n9199,n12968);
  nand U13897(n12968,n13263,n9219,n8798,n8737);
  nor U13898(n13263,n9307,n7484,n8808);
  not U13899(n7455,n9236);
  nor U13900(n9236,n9247,n13157,n12985,n9101);
  not U13901(n13157,n12873);
  nor U13902(n12873,n9779,n12850,n7482);
  not U13903(n9247,n9305);
  nor U13904(n9305,n8798,n7484);
  nand U13905(n13260,G21577,n10504);
  nand U13906(n10504,n13120,n12906,n13264);
  nand U13907(n13264,G21428,n13265);
  nand U13908(n13265,n13266,n12972,n12909);
  and U13909(n12909,n13267,n13268);
  nand U13910(n13268,n13269,n7484,n9226);
  nand U13911(n13269,n13270,n9658);
  not U13912(n9658,n9227);
  nand U13913(n13270,n7468,n9087);
  or U13914(n13267,n9242,n9224);
  nand U13915(n9224,n7477,n7481,n9226);
  nor U13916(n9226,n8737,n12850,n9307);
  not U13917(n9307,n9217);
  nor U13918(n9217,n8769,n7482);
  nand U13919(n9242,n7484,n8798);
  nand U13920(n12972,n9779,n9227,n12850,n13271);
  nor U13921(n13271,n7484,n7465,n8788);
  nor U13922(n9227,n8798,n7470);
  nand U13923(n13266,n9117,n8887);
  nor U13924(n8887,n9204,n13145);
  nand U13925(n13145,n8737,n8769);
  nand U13926(n9204,n13272,n7465);
  not U13927(n9117,n7483);
  nand U13928(n7483,n13273,n13274);
  nand U13929(n13274,n13275,n12728,n13276);
  not U13930(n13275,n13277);
  nand U13931(n13273,n13278,n13279);
  nand U13932(n13279,n13280,n13281,n13282);
  or U13933(n13282,n13277,n13283);
  nand U13934(n13281,n13284,n13277);
  nand U13935(n13284,n13285,n13286);
  nand U13936(n13286,n12989,n12990,n13287);
  nand U13937(n12990,n13288,n13289);
  or U13938(n13288,n7500,G21557);
  nand U13939(n12989,n13290,n13291);
  or U13940(n13290,G21562,G21557);
  nand U13941(n13285,n13292,n13293);
  nand U13942(n13293,n13294,n13295,n13296,n13297);
  nand U13943(n13297,n13298,n13299);
  nand U13944(n13298,n8853,n13300);
  nand U13945(n13296,n13301,n13302,n13303);
  nand U13946(n13303,n13304,n13305);
  nand U13947(n13305,n7468,n13306,n8853);
  not U13948(n13304,n13307);
  nand U13949(n13302,n8853,n13300,n13308);
  not U13950(n13308,n13299);
  nand U13951(n13299,n13309,n13310,n13277,n9085);
  not U13952(n9085,G21425);
  nand U13953(n13310,G21427,n13311);
  nand U13954(n13311,G21559,n13312);
  nand U13955(n13309,n13287,n12983);
  or U13956(n12983,n13313,n13314);
  or U13957(n13314,n8826,G21559);
  nand U13958(n13300,n13226,n13315);
  nand U13959(n13301,n13316,n13317,n13318,n13319);
  nand U13960(n13319,G21427,n8916);
  nand U13961(n13318,n13315,n13226,n9118);
  nand U13962(n13315,n7468,n8788);
  nand U13963(n13317,n13306,n13307,n8853);
  nand U13964(n13307,n13320,n13321);
  nand U13965(n13321,n13322,n13323,G21427);
  nand U13966(n13323,G21560,n13312);
  nand U13967(n13322,G21567,n9149,G21795);
  nand U13968(n13320,n13287,n12988);
  nand U13969(n12988,n13324,n13325,n13326);
  or U13970(n13326,n8913,n13327);
  nand U13971(n13325,n13327,G21560,G21565);
  not U13972(n13327,n13328);
  nand U13973(n13324,n13329,n8906);
  or U13974(n13329,G21560,n13328);
  nand U13975(n13306,n12967,n13330);
  nand U13976(n13330,n8769,n8788);
  not U13977(n12967,n9087);
  nor U13978(n9087,n7470,n7481);
  nand U13979(n13316,n13287,n12987);
  nand U13980(n12987,n13328,n13331);
  nand U13981(n13331,G21566,n8916);
  nand U13982(n13295,G21427,n8896);
  nand U13983(n13294,n13332,n13287);
  not U13984(n13332,n12976);
  or U13985(n12976,n13333,n13334);
  or U13986(n13334,n8825,G21558);
  nand U13987(n13292,G21425,G21557);
  or U13988(n13280,n12728,n13277);
  nand U13989(n13277,n8769,n8798,n8853);
  nand U13990(n12728,n13335,n13336,n13337,n13338);
  nor U13991(n13338,n13339,n13340,n13341,n13342);
  nor U13992(n13342,n10333,n8714);
  nand U13993(n8714,n13343,n13344);
  nor U13994(n13341,n10335,n8636);
  nand U13995(n8636,n13345,n13343);
  nor U13996(n13340,n10337,n8554);
  nand U13997(n8554,n13343,n13346);
  nor U13998(n13339,n10345,n8398);
  nand U13999(n8398,n13347,n13344);
  nor U14000(n13337,n13348,n13349,n13350,n13351);
  nor U14001(n13351,n10347,n8320);
  nand U14002(n8320,n13345,n13347);
  nor U14003(n13350,n10349,n8240);
  nand U14004(n8240,n13346,n13347);
  nor U14005(n13349,n10371,n8082);
  nand U14006(n8082,n13352,n13344);
  nor U14007(n13348,n10369,n8004);
  nand U14008(n8004,n13352,n13345);
  nor U14009(n13336,n13353,n13354,n13355,n13356);
  nor U14010(n13356,n10367,n7924);
  nand U14011(n7924,n13352,n13346);
  nor U14012(n13355,n10359,n7762);
  nand U14013(n7762,n13357,n13344);
  nor U14014(n13344,n9162,n9109);
  nor U14015(n13354,n10357,n7682);
  nand U14016(n7682,n13357,n13345);
  nor U14017(n13345,n9137,n9149);
  nor U14018(n13353,n10355,n7596);
  nand U14019(n7596,n13357,n13346);
  nor U14020(n13346,n9149,n9109);
  not U14021(n9109,n9137);
  nor U14022(n13335,n13358,n13359,n13360,n13361);
  nor U14023(n13361,n10331,n8829);
  nand U14024(n8829,n13362,n13343);
  nor U14025(n13343,n9179,n9196);
  nor U14026(n13360,n10343,n8476);
  nand U14027(n8476,n13362,n13347);
  nor U14028(n13347,n9196,n9171);
  nor U14029(n13359,n10373,n8160);
  nand U14030(n8160,n13362,n13352);
  nor U14031(n13352,n9179,n13363);
  nor U14032(n13358,n10361,n7842);
  nand U14033(n7842,n13362,n13357);
  nor U14034(n13357,n13363,n9171);
  not U14035(n9171,n9179);
  nand U14036(n9179,n13364,n13365);
  nand U14037(n13365,n13366,n13367);
  not U14038(n13363,n9196);
  or U14039(n9196,n13364,n13368);
  nor U14040(n13368,n13369,n13370,n13371);
  nor U14041(n13371,n8825,n8855);
  not U14042(n8855,n9096);
  nor U14043(n13370,G21426,n8170);
  nor U14044(n8170,n8248,n8163,n13372);
  nor U14045(n13372,n8825,n7850);
  not U14046(n8163,n8099);
  nand U14047(n8099,n7932,n7850);
  nor U14048(n7932,n8826,G21563);
  nor U14049(n8248,n8825,G21564);
  and U14050(n13369,G21558,n9672);
  or U14051(n13364,n13367,n13366);
  and U14052(n13366,n13373,n13374,n13375);
  nand U14053(n13375,n9672,G21559);
  nand U14054(n13374,n7854,n7456);
  not U14055(n7854,n8169);
  or U14056(n8169,n7850,n8826);
  nor U14057(n7850,n8566,n8906);
  nand U14058(n13373,n9096,G21564);
  nand U14059(n13367,n13376,n13377);
  nand U14060(n13377,n13378,n13379);
  nand U14061(n13378,n13380,n13381);
  or U14062(n13376,n13380,n13381);
  nor U14063(n13362,n9137,n9162);
  not U14064(n9162,n9149);
  or U14065(n9149,n13382,n13381);
  nand U14066(n13381,n13383,n13384);
  nand U14067(n13384,n8841,n13385);
  or U14068(n13385,n7426,n13386);
  nor U14069(n13386,n11480,n9655);
  nand U14070(n9655,n13387,n13388);
  nand U14071(n13388,G21427,n7044);
  not U14072(n7044,G21598);
  nand U14073(n13387,n9118,n9345);
  not U14074(n9345,G21757);
  not U14075(n7426,G21568);
  nand U14076(n13383,n9219,n9672);
  or U14077(n13382,n13380,n13379);
  nand U14078(n13380,n13389,n13390,n13391);
  nand U14079(n13391,n9672,G21560);
  nand U14080(n13390,n8565,n7456);
  not U14081(n8565,n8723);
  nor U14082(n8723,n7690,n7770);
  nor U14083(n7770,n8906,G21566);
  nor U14084(n7690,n8566,G21565);
  nand U14085(n13389,n9096,G21565);
  nand U14086(n9137,n13392,n13379);
  nand U14087(n13379,n13393,n13394);
  or U14088(n13392,n13394,n13393);
  nand U14089(n13393,n13395,n8923,n13396,n13397);
  nand U14090(n13397,n7456,n8566);
  nand U14091(n13396,n9096,G21566);
  nor U14092(n9096,n7456,G21428);
  nand U14093(n13395,n9672,G21561);
  nor U14094(n9672,n8843,G21427);
  or U14095(n13394,n13398,n9148,n8843);
  nor U14096(n9148,n11480,n9118);
  not U14097(n11480,G21567);
  and U14098(n13398,n8923,n13399);
  nand U14099(n13399,n9086,G21426);
  nor U14100(n9086,n7482,n9101,n12985);
  not U14101(n12985,n9219);
  nor U14102(n9219,n8788,n7477);
  not U14103(n8923,n8841);
  nor U14104(n8841,n9118,n7456);
  not U14105(n7456,G21426);
  not U14106(n13278,n13276);
  nand U14107(n13276,n13400,n13401);
  nand U14108(n13401,G21427,n13312,G21557);
  not U14109(n13312,G21795);
  nand U14110(n13400,n13287,n12974);
  nand U14111(n12974,n13402,n13403);
  nand U14112(n13403,n13404,n7500);
  not U14113(n7500,G21562);
  nand U14114(n13404,n13291,n8874);
  not U14115(n8874,G21557);
  not U14116(n13291,n13289);
  nand U14117(n13402,G21557,n13289);
  nand U14118(n13289,n13405,n13406);
  nand U14119(n13406,n13407,n8825);
  not U14120(n8825,G21563);
  or U14121(n13407,n13333,G21558);
  nand U14122(n13405,G21558,n13333);
  nand U14123(n13333,n13408,n13409);
  nand U14124(n13409,n13410,n8826);
  not U14125(n8826,G21564);
  nand U14126(n13410,n8919,n13313);
  or U14127(n13408,n8919,n13313);
  nand U14128(n13313,n8913,n13411);
  nand U14129(n13411,n13412,n13328);
  nand U14130(n13328,G21561,n8566);
  not U14131(n8566,G21566);
  nand U14132(n13412,G21560,n8906);
  not U14133(n8906,G21565);
  nand U14134(n8913,G21565,n10990);
  and U14135(n13287,n8853,n13413);
  nand U14136(n13413,n13283,n13226);
  not U14137(n13226,n9657);
  nor U14138(n9657,n8798,n7477);
  nor U14139(n13283,n7481,n7477,n9779);
  not U14140(n7481,n8788);
  nor U14141(n8853,G21425,G21427);
  not U14142(n12906,n10040);
  nor U14143(n10040,n7450,n8843);
  not U14144(n8843,G21428);
  not U14145(n7450,n9231);
  nor U14146(n9231,n8737,n7470,n8884);
  nand U14147(n8884,n9310,n7482);
  and U14148(n9310,n9779,n13272);
  nor U14149(n13272,n12850,n7468,n12765);
  not U14150(n12850,n8808);
  nand U14151(n8808,n13414,n13415,n13416,n13417);
  nor U14152(n13417,n13418,n13419,n13420,n13421);
  nor U14153(n13421,n13422,n10333);
  not U14154(n10333,G21437);
  nor U14155(n13420,n13423,n10335);
  not U14156(n10335,G21445);
  nor U14157(n13419,n13424,n10337);
  not U14158(n10337,G21453);
  nor U14159(n13418,n13425,n10345);
  not U14160(n10345,G21469);
  nor U14161(n13416,n13426,n13427,n13428,n13429);
  nor U14162(n13429,n13430,n10347);
  not U14163(n10347,G21477);
  nor U14164(n13428,n13431,n10349);
  not U14165(n10349,G21485);
  nor U14166(n13427,n13432,n10371);
  not U14167(n10371,G21501);
  nor U14168(n13426,n13433,n10369);
  not U14169(n10369,G21509);
  nor U14170(n13415,n13434,n13435,n13436,n13437);
  nor U14171(n13437,n13438,n10367);
  not U14172(n10367,G21517);
  nor U14173(n13436,n13439,n10359);
  not U14174(n10359,G21533);
  nor U14175(n13435,n13440,n10357);
  not U14176(n10357,G21541);
  nor U14177(n13434,n13441,n10355);
  not U14178(n10355,G21549);
  nor U14179(n13414,n13442,n13443,n13444,n13445);
  nor U14180(n13445,n13446,n10331);
  not U14181(n10331,G21429);
  nor U14182(n13444,n13447,n10343);
  not U14183(n10343,G21461);
  nor U14184(n13443,n13448,n10373);
  not U14185(n10373,G21493);
  nor U14186(n13442,n13449,n10361);
  not U14187(n10361,G21525);
  nand U14188(n13120,G21428,n10143,n12971);
  and U14189(n12971,n9210,n9779,n13450);
  nor U14190(n13450,n12765,n7468,n7465);
  not U14191(n7465,n7482);
  nand U14192(n7482,n13451,n13452,n13453,n13454);
  nor U14193(n13454,n13455,n13456,n13457,n13458);
  nor U14194(n13458,n13422,n10775);
  not U14195(n10775,G21442);
  nor U14196(n13457,n13423,n10776);
  not U14197(n10776,G21450);
  nor U14198(n13456,n13424,n10777);
  not U14199(n10777,G21458);
  nor U14200(n13455,n13425,n10783);
  not U14201(n10783,G21474);
  nor U14202(n13453,n13459,n13460,n13461,n13462);
  nor U14203(n13462,n13430,n10784);
  not U14204(n10784,G21482);
  nor U14205(n13461,n13431,n10785);
  not U14206(n10785,G21490);
  nor U14207(n13460,n13432,n10800);
  not U14208(n10800,G21506);
  nor U14209(n13459,n13433,n10799);
  not U14210(n10799,G21514);
  nor U14211(n13452,n13463,n13464,n13465,n13466);
  nor U14212(n13466,n13438,n10798);
  not U14213(n10798,G21522);
  nor U14214(n13465,n13439,n10792);
  not U14215(n10792,G21538);
  nor U14216(n13464,n13440,n10791);
  not U14217(n10791,G21546);
  nor U14218(n13463,n13441,n10790);
  not U14219(n10790,G21554);
  nor U14220(n13451,n13467,n13468,n13469,n13470);
  nor U14221(n13470,n13446,n10774);
  not U14222(n10774,G21434);
  nor U14223(n13469,n13447,n10782);
  not U14224(n10782,G21466);
  nor U14225(n13468,n13448,n10801);
  not U14226(n10801,G21498);
  nor U14227(n13467,n13449,n10793);
  not U14228(n10793,G21530);
  not U14229(n7468,n8798);
  nand U14230(n8798,n13471,n13472,n13473,n13474);
  nor U14231(n13474,n13475,n13476,n13477,n13478);
  nor U14232(n13478,n13422,n10432);
  not U14233(n10432,G21438);
  nor U14234(n13477,n13423,n10433);
  not U14235(n10433,G21446);
  nor U14236(n13476,n13424,n10434);
  not U14237(n10434,G21454);
  nor U14238(n13475,n13425,n10440);
  not U14239(n10440,G21470);
  nor U14240(n13473,n13479,n13480,n13481,n13482);
  nor U14241(n13482,n13430,n10441);
  not U14242(n10441,G21478);
  nor U14243(n13481,n13431,n10442);
  not U14244(n10442,G21486);
  nor U14245(n13480,n13432,n10457);
  not U14246(n10457,G21502);
  nor U14247(n13479,n13433,n10456);
  not U14248(n10456,G21510);
  nor U14249(n13472,n13483,n13484,n13485,n13486);
  nor U14250(n13486,n13438,n10455);
  not U14251(n10455,G21518);
  nor U14252(n13485,n13439,n10449);
  not U14253(n10449,G21534);
  nor U14254(n13484,n13440,n10448);
  not U14255(n10448,G21542);
  nor U14256(n13483,n13441,n10447);
  not U14257(n10447,G21550);
  nor U14258(n13471,n13487,n13488,n13489,n13490);
  nor U14259(n13490,n13446,n10431);
  not U14260(n10431,G21430);
  nor U14261(n13489,n13447,n10439);
  not U14262(n10439,G21462);
  nor U14263(n13488,n13448,n10458);
  not U14264(n10458,G21494);
  nor U14265(n13487,n13449,n10450);
  not U14266(n10450,G21526);
  nand U14267(n12765,n7472,n8788);
  nand U14268(n8788,n13491,n13492,n13493,n13494);
  nor U14269(n13494,n13495,n13496,n13497,n13498);
  nor U14270(n13498,n13422,n10520);
  not U14271(n10520,G21439);
  nor U14272(n13497,n13423,n10521);
  not U14273(n10521,G21447);
  nor U14274(n13496,n13424,n10522);
  not U14275(n10522,G21455);
  nor U14276(n13495,n13425,n10528);
  not U14277(n10528,G21471);
  nor U14278(n13493,n13499,n13500,n13501,n13502);
  nor U14279(n13502,n13430,n10529);
  not U14280(n10529,G21479);
  nor U14281(n13501,n13431,n10530);
  not U14282(n10530,G21487);
  nor U14283(n13500,n13432,n10545);
  not U14284(n10545,G21503);
  nor U14285(n13499,n13433,n10544);
  not U14286(n10544,G21511);
  nor U14287(n13492,n13503,n13504,n13505,n13506);
  nor U14288(n13506,n13438,n10543);
  not U14289(n10543,G21519);
  nor U14290(n13505,n13439,n10537);
  not U14291(n10537,G21535);
  nor U14292(n13504,n13440,n10536);
  not U14293(n10536,G21543);
  nor U14294(n13503,n13441,n10535);
  not U14295(n10535,G21551);
  nor U14296(n13491,n13507,n13508,n13509,n13510);
  nor U14297(n13510,n13446,n10519);
  not U14298(n10519,G21431);
  nor U14299(n13509,n13447,n10527);
  not U14300(n10527,G21463);
  nor U14301(n13508,n13448,n10546);
  not U14302(n10546,G21495);
  nor U14303(n13507,n13449,n10538);
  not U14304(n10538,G21527);
  not U14305(n7472,n7484);
  nand U14306(n7484,n13511,n13512,n13513,n13514);
  nor U14307(n13514,n13515,n13516,n13517,n13518);
  nor U14308(n13518,n13422,n10602);
  not U14309(n10602,G21440);
  nor U14310(n13517,n13423,n10603);
  not U14311(n10603,G21448);
  nor U14312(n13516,n13424,n10604);
  not U14313(n10604,G21456);
  nor U14314(n13515,n13425,n10610);
  not U14315(n10610,G21472);
  nor U14316(n13513,n13519,n13520,n13521,n13522);
  nor U14317(n13522,n13430,n10611);
  not U14318(n10611,G21480);
  nor U14319(n13521,n13431,n10612);
  not U14320(n10612,G21488);
  nor U14321(n13520,n13432,n10627);
  not U14322(n10627,G21504);
  nor U14323(n13519,n13433,n10626);
  not U14324(n10626,G21512);
  nor U14325(n13512,n13523,n13524,n13525,n13526);
  nor U14326(n13526,n13438,n10625);
  not U14327(n10625,G21520);
  nor U14328(n13525,n13439,n10619);
  not U14329(n10619,G21536);
  nor U14330(n13524,n13440,n10618);
  not U14331(n10618,G21544);
  nor U14332(n13523,n13441,n10617);
  not U14333(n10617,G21552);
  nor U14334(n13511,n13527,n13528,n13529,n13530);
  nor U14335(n13530,n13446,n10601);
  not U14336(n10601,G21432);
  nor U14337(n13529,n13447,n10609);
  not U14338(n10609,G21464);
  nor U14339(n13528,n13448,n10628);
  not U14340(n10628,G21496);
  nor U14341(n13527,n13449,n10620);
  not U14342(n10620,G21528);
  not U14343(n9779,n8769);
  nand U14344(n8769,n13531,n13532,n13533,n13534);
  nor U14345(n13534,n13535,n13536,n13537,n13538);
  nor U14346(n13538,n13422,n10689);
  not U14347(n10689,G21441);
  nor U14348(n13537,n13423,n10690);
  not U14349(n10690,G21449);
  nor U14350(n13536,n13424,n10691);
  not U14351(n10691,G21457);
  nor U14352(n13535,n13425,n10697);
  not U14353(n10697,G21473);
  nor U14354(n13533,n13539,n13540,n13541,n13542);
  nor U14355(n13542,n13430,n10698);
  not U14356(n10698,G21481);
  nor U14357(n13541,n13431,n10699);
  not U14358(n10699,G21489);
  nor U14359(n13540,n13432,n10714);
  not U14360(n10714,G21505);
  nor U14361(n13539,n13433,n10713);
  not U14362(n10713,G21513);
  nor U14363(n13532,n13543,n13544,n13545,n13546);
  nor U14364(n13546,n13438,n10712);
  not U14365(n10712,G21521);
  nor U14366(n13545,n13439,n10706);
  not U14367(n10706,G21537);
  nor U14368(n13544,n13440,n10705);
  not U14369(n10705,G21545);
  nor U14370(n13543,n13441,n10704);
  not U14371(n10704,G21553);
  nor U14372(n13531,n13547,n13548,n13549,n13550);
  nor U14373(n13550,n13446,n10688);
  not U14374(n10688,G21433);
  nor U14375(n13549,n13447,n10696);
  not U14376(n10696,G21465);
  nor U14377(n13548,n13448,n10715);
  not U14378(n10715,G21497);
  nor U14379(n13547,n13449,n10707);
  not U14380(n10707,G21529);
  nor U14381(n9210,n8737,n7477);
  not U14382(n7477,n7470);
  nand U14383(n7470,n13551,n13552,n13553,n13554);
  nor U14384(n13554,n13555,n13556,n13557,n13558);
  nor U14385(n13558,n13422,n10864);
  not U14386(n10864,G21443);
  nor U14387(n13557,n13423,n10865);
  not U14388(n10865,G21451);
  nor U14389(n13556,n13424,n10866);
  not U14390(n10866,G21459);
  nor U14391(n13555,n13425,n10872);
  not U14392(n10872,G21475);
  nor U14393(n13553,n13559,n13560,n13561,n13562);
  nor U14394(n13562,n13430,n10873);
  not U14395(n10873,G21483);
  nor U14396(n13561,n13431,n10874);
  not U14397(n10874,G21491);
  nor U14398(n13560,n13432,n10889);
  not U14399(n10889,G21507);
  nor U14400(n13559,n13433,n10888);
  not U14401(n10888,G21515);
  nor U14402(n13552,n13563,n13564,n13565,n13566);
  nor U14403(n13566,n13438,n10887);
  not U14404(n10887,G21523);
  nor U14405(n13565,n13439,n10881);
  not U14406(n10881,G21539);
  nor U14407(n13564,n13440,n10880);
  not U14408(n10880,G21547);
  nor U14409(n13563,n13441,n10879);
  not U14410(n10879,G21555);
  nor U14411(n13551,n13567,n13568,n13569,n13570);
  nor U14412(n13570,n13446,n10863);
  not U14413(n10863,G21435);
  nor U14414(n13569,n13447,n10871);
  not U14415(n10871,G21467);
  nor U14416(n13568,n13448,n10890);
  not U14417(n10890,G21499);
  nor U14418(n13567,n13449,n10882);
  not U14419(n10882,G21531);
  nor U14420(n13574,n13575,n13576,n13577,n13578);
  nor U14421(n13578,n13422,n10952);
  not U14422(n10952,G21444);
  nand U14423(n13422,n13579,n10989);
  nor U14424(n13577,n13423,n10954);
  not U14425(n10954,G21452);
  nand U14426(n13423,n9160,n13579);
  nor U14427(n13576,n13424,n10956);
  not U14428(n10956,G21460);
  nand U14429(n13424,n8915,n13579);
  nor U14430(n13575,n13425,n10963);
  not U14431(n10963,G21476);
  nand U14432(n13425,n13257,n10989);
  nor U14433(n13573,n13580,n13581,n13582,n13583);
  nor U14434(n13583,n13430,n10964);
  not U14435(n10964,G21484);
  nand U14436(n13430,n9160,n13257);
  nor U14437(n13582,n13431,n10967);
  not U14438(n10967,G21492);
  nand U14439(n13431,n8915,n13257);
  nor U14440(n13581,n13432,n10986);
  not U14441(n10986,G21508);
  nand U14442(n13432,n13258,n10989);
  nor U14443(n13580,n13433,n10985);
  not U14444(n10985,G21516);
  nand U14445(n13433,n13258,n9160);
  nor U14446(n13572,n13584,n13585,n13586,n13587);
  nor U14447(n13587,n13438,n10984);
  not U14448(n10984,G21524);
  nand U14449(n13438,n13258,n8915);
  nor U14450(n13586,n13439,n10976);
  not U14451(n10976,G21540);
  nand U14452(n13439,n10994,n10989);
  nor U14453(n10989,n10990,G21561);
  nor U14454(n13585,n13440,n10974);
  not U14455(n10974,G21548);
  nand U14456(n13440,n10994,n9160);
  nor U14457(n9160,n8916,G21560);
  nor U14458(n13584,n13441,n10972);
  not U14459(n10972,G21556);
  nand U14460(n13441,n10994,n8915);
  nor U14461(n8915,G21560,G21561);
  nor U14462(n13571,n13588,n13589,n13590,n13591);
  nor U14463(n13591,n13446,n10949);
  not U14464(n10949,G21436);
  nand U14465(n13446,n10997,n13579);
  nor U14466(n13579,n8896,n8919);
  nor U14467(n13590,n13447,n10961);
  not U14468(n10961,G21468);
  nand U14469(n13447,n10997,n13257);
  nor U14470(n13257,n8896,G21559);
  not U14471(n8896,G21558);
  nor U14472(n13589,n13448,n10987);
  not U14473(n10987,G21500);
  nand U14474(n13448,n10997,n13258);
  nor U14475(n13258,n8919,G21558);
  not U14476(n8919,G21559);
  nor U14477(n13588,n13449,n10977);
  not U14478(n10977,G21532);
  nand U14479(n13449,n10997,n10994);
  nor U14480(n10994,G21558,G21559);
  nor U14481(n10997,n10990,n8916);
  not U14482(n8916,G21561);
  not U14483(n10990,G21560);
  nand U14484(n10143,n8955,n13592);
  nand U14485(n13592,G21390,n8964);
  not U14486(n8964,G21391);
  nand U14487(n8955,G21391,n8980);
  not U14488(n8980,G21390);
  nand U14489(n13259,G21609,n7590);
  not U14490(n9118,G21427);
endmodule

