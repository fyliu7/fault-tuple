
module b22s_1 ( G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, 
        G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, 
        G29, G30, G31, G32, G35973, G35974, G35975, G35976, G35977, G35978, 
        G35979, G35980, G35981, G35982, G35983, G35984, G35985, G35986, G35987, 
        G35988, G35989, G35990, G35991, G35992, G35993, G35994, G35995, G35996, 
        G35997, G35998, G35999, G36000, G36001, G36002, G36003, G36004, G36005, 
        G36006, G36007, G36008, G36009, G36010, G36011, G36012, G36013, G36014, 
        G36015, G36016, G36017, G36018, G36019, G36020, G36021, G36022, G36023, 
        G36024, G36025, G36026, G36027, G36028, G36029, G36030, G36031, G36032, 
        G36033, G36034, G36035, G36036, G36037, G36038, G36039, G36040, G36041, 
        G36042, G36043, G36044, G36045, G36046, G36047, G36048, G36049, G36050, 
        G36051, G36052, G36053, G36054, G36055, G36056, G36057, G36058, G36059, 
        G36060, G36061, G36062, G36063, G36064, G36065, G36066, G36067, G36068, 
        G36069, G36070, G36071, G36072, G36073, G36074, G36075, G36076, G36077, 
        G36078, G36079, G36080, G36081, G36082, G36083, G36084, G36085, G36086, 
        G36087, G36088, G36089, G36090, G36091, G36092, G36093, G36094, G36095, 
        G36096, G36097, G36098, G36099, G36100, G36101, G36102, G36103, G36104, 
        G36105, G36106, G36107, G36108, G36109, G36110, G36111, G36112, G36113, 
        G36114, G36115, G36116, G36117, G36118, G36119, G36120, G36121, G36122, 
        G36123, G36124, G36125, G36126, G36127, G36128, G36129, G36130, G36131, 
        G36132, G36133, G36134, G36135, G36136, G36137, G36138, G36139, G36140, 
        G36141, G36142, G36143, G36144, G36145, G36146, G36147, G36148, G36149, 
        G36150, G36151, G36152, G36153, G36154, G36155, G36156, G36157, G36158, 
        G36159, G36160, G36161, G36162, G36163, G36164, G36165, G36166, G36167, 
        G36168, G36169, G36170, G36171, G36172, G36173, G36174, G36175, G36176, 
        G36177, G36178, G36179, G36180, G36181, G36182, G36183, G36184, G36185, 
        G36186, G36187, G36188, G36189, G36190, G36191, G36192, G36193, G36194, 
        G36195, G36196, G36197, G36198, G36199, G36200, G36201, G36202, G36203, 
        G36204, G36205, G36206, G36207, G36208, G36209, G36210, G36211, G36212, 
        G36213, G36214, G36215, G36216, G36217, G36218, G36219, G36220, G36221, 
        G36222, G36223, G36224, G36225, G36226, G36227, G36228, G36229, G36230, 
        G36231, G36232, G36233, G36234, G36235, G36236, G36237, G36238, G36239, 
        G36240, G36241, G36242, G36243, G36244, G36245, G36246, G36247, G36248, 
        G36249, G36250, G36251, G36252, G36253, G36254, G36255, G36256, G36257, 
        G36258, G36259, G36260, G36261, G36262, G36263, G36264, G36265, G36266, 
        G36267, G36268, G36269, G36270, G36271, G36272, G36273, G36274, G36275, 
        G36276, G36277, G36278, G36279, G36280, G36281, G36282, G36283, G36284, 
        G36285, G36286, G36287, G36288, G36289, G36290, G36291, G36292, G36293, 
        G36294, G36295, G36296, G36297, G36298, G36299, G36300, G36301, G36302, 
        G36303, G36304, G36305, G36306, G36307, G36308, G36309, G36310, G36311, 
        G36312, G36313, G36314, G36315, G36316, G36317, G36318, G36319, G36320, 
        G36321, G36322, G36323, G36324, G36325, G36326, G36327, G36328, G36329, 
        G36330, G36331, G36332, G36333, G36334, G36335, G36336, G36337, G36338, 
        G36339, G36340, G36341, G36342, G36343, G36344, G36345, G36346, G36347, 
        G36348, G36349, G36350, G36351, G36352, G36353, G36354, G36355, G36356, 
        G36357, G36358, G36359, G36360, G36361, G36362, G36363, G36364, G36365, 
        G36366, G36367, G36368, G36369, G36370, G36371, G36372, G36373, G36374, 
        G36375, G36376, G36377, G36378, G36379, G36380, G36381, G36382, G36383, 
        G36384, G36385, G36386, G36387, G36388, G36389, G36390, G36391, G36392, 
        G36393, G36394, G36395, G36396, G36397, G36398, G36399, G36400, G36401, 
        G36402, G36403, G36404, G36405, G36406, G36407, G36408, G36409, G36410, 
        G36411, G36412, G36413, G36414, G36415, G36416, G36417, G36418, G36419, 
        G36420, G36421, G36422, G36423, G36424, G36425, G36426, G36427, G36428, 
        G36429, G36430, G36431, G36432, G36433, G36434, G36435, G36436, G36437, 
        G36438, G36439, G36440, G36441, G36442, G36443, G36444, G36445, G36446, 
        G36447, G36448, G36449, G36450, G36451, G36452, G36453, G36454, G36455, 
        G36456, G36457, G36458, G36459, G36460, G36461, G36462, G36463, G36464, 
        G36465, G36466, G36467, G36468, G36469, G36470, G36471, G36472, G36473, 
        G36474, G36475, G36476, G36477, G36478, G36479, G36480, G36481, G36482, 
        G36483, G36484, G36485, G36486, G36487, G36488, G36489, G36490, G36491, 
        G36492, G36493, G36494, G36495, G36496, G36497, G36498, G36499, G36500, 
        G36501, G36502, G36503, G36504, G36505, G36506, G36507, G36508, G36509, 
        G36510, G36511, G36512, G36513, G36514, G36515, G36516, G36517, G36518, 
        G36519, G36520, G36521, G36522, G36523, G36524, G36525, G36526, G36527, 
        G36528, G36529, G36530, G36531, G36532, G36533, G36534, G36535, G36536, 
        G36537, G36538, G36539, G36540, G36541, G36542, G36543, G36544, G36545, 
        G36546, G36547, G36548, G36549, G36550, G36551, G36552, G36553, G36554, 
        G36555, G36556, G36557, G36558, G36559, G36560, G36561, G36562, G36563, 
        G36564, G36565, G36566, G36567, G36568, G36569, G36570, G36571, G36572, 
        G36573, G36574, G36575, G36576, G36577, G36578, G36579, G36580, G36581, 
        G36582, G36583, G36584, G36585, G36586, G36587, G36588, G36589, G36590, 
        G36591, G36592, G36593, G36594, G36595, G36596, G36597, G36598, G36599, 
        G36600, G36601, G36602, G36603, G36604, G36605, G36606, G36607, G36608, 
        G36609, G36610, G36611, G36612, G36613, G36614, G36615, G36616, G36617, 
        G36618, G36619, G36620, G36621, G36622, G36623, G36624, G36625, G36626, 
        G36627, G36628, G36629, G36630, G36631, G36632, G36633, G36634, G36635, 
        G36636, G36637, G36638, G36639, G36640, G36641, G36642, G36643, G36644, 
        G36645, G36646, G36647, G36648, G36649, G36650, G36651, G36652, G36653, 
        G36654, G36655, G36656, G36657, G36658, G36659, G36660, G36661, G36662, 
        G36663, G36664, G36665, G36666, G36667, G36668, G36669, G36670, G36671, 
        G36672, G36673, G36674, G36675, G36676, G36677, G36678, G36679, G36680, 
        G36681, G36682, G36683, G36684, G36685, G36686, G36687, G36688, G36689, 
        G36690, G36691, G36692, G36693, G36694, G36695, G36696, G36697, G36698, 
        G36699, G36700, G36701, G36702, G36703, G36704, G36705, G36706, G36707, 
        G10148, G10226, G10228, G10230, G10232, G10234, G10236, G10238, G10240, 
        G10242, G10208, G10210, G10212, G10214, G10216, G10218, G10220, G10222, 
        G10188, G10149, G792, G793, G1407, G1408, G1409, G1410, G1411, G1412, 
        G1413, G1414, G1415, G1416, G1417, G1418, G1419, G1420, G1421, G1422, 
        G1423, G1424, G1425, G1426, G1427, G1428, G1429, G1430, G1431, G1432, 
        G1433, G1434, G1435, G1436, G1437, G1438, G1715, G1716, G1439, G1440, 
        G1441, G1442, G1443, G1444, G1445, G1446, G1447, G1448, G1449, G1450, 
        G1451, G1452, G1453, G1454, G1455, G1456, G1457, G1458, G1459, G1460, 
        G1461, G1462, G1463, G1464, G1465, G1466, G1467, G1468, G1727, G1730, 
        G1733, G1736, G1739, G1742, G1745, G1748, G1751, G1754, G1757, G1760, 
        G1763, G1766, G1769, G1772, G1775, G1778, G1781, G1783, G1784, G1785, 
        G1786, G1787, G1788, G1789, G1790, G1791, G1792, G1793, G1794, G1795, 
        G1796, G1797, G1798, G1799, G1800, G1801, G1802, G1803, G1804, G1805, 
        G1806, G1807, G1808, G1809, G1810, G1811, G1812, G1813, G1814, G1815, 
        G1816, G1817, G1818, G1819, G1820, G1821, G1822, G1823, G1824, G1825, 
        G1826, G1827, G1469, G1828, G1470, G1471, G1472, G1473, G1474, G1475, 
        G1476, G1477, G1478, G1479, G1480, G1481, G1482, G1483, G1484, G1485, 
        G1486, G1487, G1488, G1489, G1490, G1491, G1492, G1493, G1494, G1495, 
        G1496, G1497, G1498, G1499, G1500, G1501, G1502, G1503, G1504, G1505, 
        G1506, G1507, G1508, G1509, G1510, G1511, G1512, G1513, G1514, G1515, 
        G1516, G1517, G1518, G1519, G1829, G1830, G1831, G1832, G1833, G1834, 
        G1835, G1836, G1837, G1838, G1839, G1840, G1841, G1842, G1843, G1844, 
        G1845, G1846, G1847, G1848, G1849, G1850, G1851, G1852, G1853, G1854, 
        G1855, G1856, G1857, G1858, G1859, G1860, G1520, G1521, G1522, G1523, 
        G1524, G1525, G1526, G1527, G1528, G1529, G1530, G1531, G1532, G1533, 
        G1534, G1535, G1536, G1537, G1538, G1539, G1540, G1541, G1542, G1543, 
        G1544, G1545, G1546, G1547, G1548, G1549, G1406, G1341, G1625, G4390, 
        G4391, G4392, G4393, G4394, G4395, G4396, G4397, G4398, G4399, G4400, 
        G4401, G4402, G4403, G4404, G4405, G4406, G4407, G4408, G4409, G4410, 
        G4411, G4412, G4413, G4414, G4415, G4416, G4417, G4418, G4419, G4420, 
        G4421, G4692, G4693, G4422, G4423, G4424, G4425, G4426, G4427, G4428, 
        G4429, G4430, G4431, G4432, G4433, G4434, G4435, G4436, G4437, G4438, 
        G4439, G4440, G4441, G4442, G4443, G4444, G4445, G4446, G4447, G4448, 
        G4449, G4450, G4451, G4704, G4707, G4710, G4713, G4716, G4719, G4722, 
        G4725, G4728, G4731, G4734, G4737, G4740, G4743, G4746, G4749, G4752, 
        G4755, G4758, G4760, G4761, G4762, G4763, G4764, G4765, G4766, G4767, 
        G4768, G4769, G4770, G4771, G4772, G4773, G4774, G4775, G4776, G4777, 
        G4778, G4779, G4780, G4781, G4782, G4783, G4784, G4785, G4786, G4787, 
        G4788, G4789, G4790, G4791, G4792, G4793, G4794, G4795, G4796, G4797, 
        G4798, G4799, G4800, G4801, G4802, G4803, G4804, G4452, G4453, G4454, 
        G4455, G4456, G4457, G4458, G4459, G4460, G4461, G4462, G4463, G4464, 
        G4465, G4466, G4467, G4468, G4469, G4470, G4471, G4472, G4473, G4474, 
        G4475, G4476, G4477, G4478, G4479, G4480, G4481, G4482, G4483, G4484, 
        G4485, G4486, G4487, G4488, G4489, G4490, G4491, G4492, G4493, G4494, 
        G4495, G4496, G4497, G4498, G4499, G4500, G4501, G4502, G4503, G4805, 
        G4806, G4807, G4808, G4809, G4810, G4811, G4812, G4813, G4814, G4815, 
        G4816, G4817, G4818, G4819, G4820, G4821, G4822, G4823, G4824, G4825, 
        G4826, G4827, G4828, G4829, G4830, G4831, G4832, G4833, G4834, G4835, 
        G4836, G4504, G4505, G4506, G4507, G4508, G4509, G4510, G4511, G4512, 
        G4513, G4514, G4515, G4516, G4517, G4518, G4519, G4520, G4521, G4522, 
        G4523, G4524, G4525, G4526, G4527, G4528, G4529, G4530, G4531, G4532, 
        G4533, G4389, G4388, G4591, G7318, G7319, G7320, G7321, G7322, G7323, 
        G7324, G7325, G7326, G7327, G7328, G7329, G7330, G7331, G7332, G7333, 
        G7334, G7335, G7336, G7337, G7338, G7339, G7340, G7341, G7342, G7343, 
        G7344, G7345, G7346, G7347, G7348, G7349, G7660, G7661, G7350, G7351, 
        G7352, G7353, G7354, G7355, G7356, G7357, G7358, G7359, G7360, G7361, 
        G7362, G7363, G7364, G7365, G7366, G7367, G7368, G7369, G7370, G7371, 
        G7372, G7373, G7374, G7375, G7376, G7377, G7378, G7379, G7380, G7381, 
        G7382, G7383, G7384, G7385, G7386, G7387, G7388, G7389, G7390, G7391, 
        G7392, G7393, G7394, G7395, G7396, G7397, G7398, G7399, G7400, G7401, 
        G7402, G7403, G7404, G7405, G7406, G7407, G7408, G7409, G7410, G7411, 
        G7412, G7413, G7414, G7415, G7416, G7417, G7418, G7419, G7420, G7421, 
        G7422, G7423, G7424, G7425, G7426, G7427, G7428, G7429, G7430, G7431, 
        G7432, G7433, G7434, G7435, G7436, G7437, G7438, G7439, G7440, G7441, 
        G7442, G7443, G7444, G7445, G7446, G7447, G7448, G7449, G7450, G7451, 
        G7452, G7453, G7454, G7455, G7456, G7457, G7458, G7459, G7460, G7461, 
        G7462, G7463, G7464, G7465, G7466, G7467, G7468, G7469, G7470, G7471, 
        G7472, G7473, G7474, G7475, G7476, G7477, G7478, G7479, G7480, G7481, 
        G7482, G7483, G7484, G7485, G7486, G7487, G7488, G7489, G7490, G7491, 
        G7492, G7493, G7494, G7495, G7689, G7690, G7691, G7692, G7693, G7694, 
        G7695, G7696, G7697, G7698, G7699, G7700, G7701, G7702, G7703, G7704, 
        G7705, G7706, G7707, G7708, G7709, G7710, G7711, G7712, G7713, G7714, 
        G7715, G7716, G7717, G7718, G7719, G7720, G7496, G7497, G7498, G7499, 
        G7500, G7501, G7502, G7503, G7504, G7505, G7506, G7507, G7508, G7509, 
        G7510, G7511, G7512, G7513, G7514, G7515, G7516, G7517, G7518, G7519, 
        G7520, G7521, G7522, G7523, G7524, G7525, G7317, G7316, G7605 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
         G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
         G31, G32, G35973, G35974, G35975, G35976, G35977, G35978, G35979,
         G35980, G35981, G35982, G35983, G35984, G35985, G35986, G35987,
         G35988, G35989, G35990, G35991, G35992, G35993, G35994, G35995,
         G35996, G35997, G35998, G35999, G36000, G36001, G36002, G36003,
         G36004, G36005, G36006, G36007, G36008, G36009, G36010, G36011,
         G36012, G36013, G36014, G36015, G36016, G36017, G36018, G36019,
         G36020, G36021, G36022, G36023, G36024, G36025, G36026, G36027,
         G36028, G36029, G36030, G36031, G36032, G36033, G36034, G36035,
         G36036, G36037, G36038, G36039, G36040, G36041, G36042, G36043,
         G36044, G36045, G36046, G36047, G36048, G36049, G36050, G36051,
         G36052, G36053, G36054, G36055, G36056, G36057, G36058, G36059,
         G36060, G36061, G36062, G36063, G36064, G36065, G36066, G36067,
         G36068, G36069, G36070, G36071, G36072, G36073, G36074, G36075,
         G36076, G36077, G36078, G36079, G36080, G36081, G36082, G36083,
         G36084, G36085, G36086, G36087, G36088, G36089, G36090, G36091,
         G36092, G36093, G36094, G36095, G36096, G36097, G36098, G36099,
         G36100, G36101, G36102, G36103, G36104, G36105, G36106, G36107,
         G36108, G36109, G36110, G36111, G36112, G36113, G36114, G36115,
         G36116, G36117, G36118, G36119, G36120, G36121, G36122, G36123,
         G36124, G36125, G36126, G36127, G36128, G36129, G36130, G36131,
         G36132, G36133, G36134, G36135, G36136, G36137, G36138, G36139,
         G36140, G36141, G36142, G36143, G36144, G36145, G36146, G36147,
         G36148, G36149, G36150, G36151, G36152, G36153, G36154, G36155,
         G36156, G36157, G36158, G36159, G36160, G36161, G36162, G36163,
         G36164, G36165, G36166, G36167, G36168, G36169, G36170, G36171,
         G36172, G36173, G36174, G36175, G36176, G36177, G36178, G36179,
         G36180, G36181, G36182, G36183, G36184, G36185, G36186, G36187,
         G36188, G36189, G36190, G36191, G36192, G36193, G36194, G36195,
         G36196, G36197, G36198, G36199, G36200, G36201, G36202, G36203,
         G36204, G36205, G36206, G36207, G36208, G36209, G36210, G36211,
         G36212, G36213, G36214, G36215, G36216, G36217, G36218, G36219,
         G36220, G36221, G36222, G36223, G36224, G36225, G36226, G36227,
         G36228, G36229, G36230, G36231, G36232, G36233, G36234, G36235,
         G36236, G36237, G36238, G36239, G36240, G36241, G36242, G36243,
         G36244, G36245, G36246, G36247, G36248, G36249, G36250, G36251,
         G36252, G36253, G36254, G36255, G36256, G36257, G36258, G36259,
         G36260, G36261, G36262, G36263, G36264, G36265, G36266, G36267,
         G36268, G36269, G36270, G36271, G36272, G36273, G36274, G36275,
         G36276, G36277, G36278, G36279, G36280, G36281, G36282, G36283,
         G36284, G36285, G36286, G36287, G36288, G36289, G36290, G36291,
         G36292, G36293, G36294, G36295, G36296, G36297, G36298, G36299,
         G36300, G36301, G36302, G36303, G36304, G36305, G36306, G36307,
         G36308, G36309, G36310, G36311, G36312, G36313, G36314, G36315,
         G36316, G36317, G36318, G36319, G36320, G36321, G36322, G36323,
         G36324, G36325, G36326, G36327, G36328, G36329, G36330, G36331,
         G36332, G36333, G36334, G36335, G36336, G36337, G36338, G36339,
         G36340, G36341, G36342, G36343, G36344, G36345, G36346, G36347,
         G36348, G36349, G36350, G36351, G36352, G36353, G36354, G36355,
         G36356, G36357, G36358, G36359, G36360, G36361, G36362, G36363,
         G36364, G36365, G36366, G36367, G36368, G36369, G36370, G36371,
         G36372, G36373, G36374, G36375, G36376, G36377, G36378, G36379,
         G36380, G36381, G36382, G36383, G36384, G36385, G36386, G36387,
         G36388, G36389, G36390, G36391, G36392, G36393, G36394, G36395,
         G36396, G36397, G36398, G36399, G36400, G36401, G36402, G36403,
         G36404, G36405, G36406, G36407, G36408, G36409, G36410, G36411,
         G36412, G36413, G36414, G36415, G36416, G36417, G36418, G36419,
         G36420, G36421, G36422, G36423, G36424, G36425, G36426, G36427,
         G36428, G36429, G36430, G36431, G36432, G36433, G36434, G36435,
         G36436, G36437, G36438, G36439, G36440, G36441, G36442, G36443,
         G36444, G36445, G36446, G36447, G36448, G36449, G36450, G36451,
         G36452, G36453, G36454, G36455, G36456, G36457, G36458, G36459,
         G36460, G36461, G36462, G36463, G36464, G36465, G36466, G36467,
         G36468, G36469, G36470, G36471, G36472, G36473, G36474, G36475,
         G36476, G36477, G36478, G36479, G36480, G36481, G36482, G36483,
         G36484, G36485, G36486, G36487, G36488, G36489, G36490, G36491,
         G36492, G36493, G36494, G36495, G36496, G36497, G36498, G36499,
         G36500, G36501, G36502, G36503, G36504, G36505, G36506, G36507,
         G36508, G36509, G36510, G36511, G36512, G36513, G36514, G36515,
         G36516, G36517, G36518, G36519, G36520, G36521, G36522, G36523,
         G36524, G36525, G36526, G36527, G36528, G36529, G36530, G36531,
         G36532, G36533, G36534, G36535, G36536, G36537, G36538, G36539,
         G36540, G36541, G36542, G36543, G36544, G36545, G36546, G36547,
         G36548, G36549, G36550, G36551, G36552, G36553, G36554, G36555,
         G36556, G36557, G36558, G36559, G36560, G36561, G36562, G36563,
         G36564, G36565, G36566, G36567, G36568, G36569, G36570, G36571,
         G36572, G36573, G36574, G36575, G36576, G36577, G36578, G36579,
         G36580, G36581, G36582, G36583, G36584, G36585, G36586, G36587,
         G36588, G36589, G36590, G36591, G36592, G36593, G36594, G36595,
         G36596, G36597, G36598, G36599, G36600, G36601, G36602, G36603,
         G36604, G36605, G36606, G36607, G36608, G36609, G36610, G36611,
         G36612, G36613, G36614, G36615, G36616, G36617, G36618, G36619,
         G36620, G36621, G36622, G36623, G36624, G36625, G36626, G36627,
         G36628, G36629, G36630, G36631, G36632, G36633, G36634, G36635,
         G36636, G36637, G36638, G36639, G36640, G36641, G36642, G36643,
         G36644, G36645, G36646, G36647, G36648, G36649, G36650, G36651,
         G36652, G36653, G36654, G36655, G36656, G36657, G36658, G36659,
         G36660, G36661, G36662, G36663, G36664, G36665, G36666, G36667,
         G36668, G36669, G36670, G36671, G36672, G36673, G36674, G36675,
         G36676, G36677, G36678, G36679, G36680, G36681, G36682, G36683,
         G36684, G36685, G36686, G36687, G36688, G36689, G36690, G36691,
         G36692, G36693, G36694, G36695, G36696, G36697, G36698, G36699,
         G36700, G36701, G36702, G36703, G36704, G36705, G36706, G36707;
  output G10148, G10226, G10228, G10230, G10232, G10234, G10236, G10238,
         G10240, G10242, G10208, G10210, G10212, G10214, G10216, G10218,
         G10220, G10222, G10188, G10149, G792, G793, G1407, G1408, G1409,
         G1410, G1411, G1412, G1413, G1414, G1415, G1416, G1417, G1418, G1419,
         G1420, G1421, G1422, G1423, G1424, G1425, G1426, G1427, G1428, G1429,
         G1430, G1431, G1432, G1433, G1434, G1435, G1436, G1437, G1438, G1715,
         G1716, G1439, G1440, G1441, G1442, G1443, G1444, G1445, G1446, G1447,
         G1448, G1449, G1450, G1451, G1452, G1453, G1454, G1455, G1456, G1457,
         G1458, G1459, G1460, G1461, G1462, G1463, G1464, G1465, G1466, G1467,
         G1468, G1727, G1730, G1733, G1736, G1739, G1742, G1745, G1748, G1751,
         G1754, G1757, G1760, G1763, G1766, G1769, G1772, G1775, G1778, G1781,
         G1783, G1784, G1785, G1786, G1787, G1788, G1789, G1790, G1791, G1792,
         G1793, G1794, G1795, G1796, G1797, G1798, G1799, G1800, G1801, G1802,
         G1803, G1804, G1805, G1806, G1807, G1808, G1809, G1810, G1811, G1812,
         G1813, G1814, G1815, G1816, G1817, G1818, G1819, G1820, G1821, G1822,
         G1823, G1824, G1825, G1826, G1827, G1469, G1828, G1470, G1471, G1472,
         G1473, G1474, G1475, G1476, G1477, G1478, G1479, G1480, G1481, G1482,
         G1483, G1484, G1485, G1486, G1487, G1488, G1489, G1490, G1491, G1492,
         G1493, G1494, G1495, G1496, G1497, G1498, G1499, G1500, G1501, G1502,
         G1503, G1504, G1505, G1506, G1507, G1508, G1509, G1510, G1511, G1512,
         G1513, G1514, G1515, G1516, G1517, G1518, G1519, G1829, G1830, G1831,
         G1832, G1833, G1834, G1835, G1836, G1837, G1838, G1839, G1840, G1841,
         G1842, G1843, G1844, G1845, G1846, G1847, G1848, G1849, G1850, G1851,
         G1852, G1853, G1854, G1855, G1856, G1857, G1858, G1859, G1860, G1520,
         G1521, G1522, G1523, G1524, G1525, G1526, G1527, G1528, G1529, G1530,
         G1531, G1532, G1533, G1534, G1535, G1536, G1537, G1538, G1539, G1540,
         G1541, G1542, G1543, G1544, G1545, G1546, G1547, G1548, G1549, G1406,
         G1341, G1625, G4390, G4391, G4392, G4393, G4394, G4395, G4396, G4397,
         G4398, G4399, G4400, G4401, G4402, G4403, G4404, G4405, G4406, G4407,
         G4408, G4409, G4410, G4411, G4412, G4413, G4414, G4415, G4416, G4417,
         G4418, G4419, G4420, G4421, G4692, G4693, G4422, G4423, G4424, G4425,
         G4426, G4427, G4428, G4429, G4430, G4431, G4432, G4433, G4434, G4435,
         G4436, G4437, G4438, G4439, G4440, G4441, G4442, G4443, G4444, G4445,
         G4446, G4447, G4448, G4449, G4450, G4451, G4704, G4707, G4710, G4713,
         G4716, G4719, G4722, G4725, G4728, G4731, G4734, G4737, G4740, G4743,
         G4746, G4749, G4752, G4755, G4758, G4760, G4761, G4762, G4763, G4764,
         G4765, G4766, G4767, G4768, G4769, G4770, G4771, G4772, G4773, G4774,
         G4775, G4776, G4777, G4778, G4779, G4780, G4781, G4782, G4783, G4784,
         G4785, G4786, G4787, G4788, G4789, G4790, G4791, G4792, G4793, G4794,
         G4795, G4796, G4797, G4798, G4799, G4800, G4801, G4802, G4803, G4804,
         G4452, G4453, G4454, G4455, G4456, G4457, G4458, G4459, G4460, G4461,
         G4462, G4463, G4464, G4465, G4466, G4467, G4468, G4469, G4470, G4471,
         G4472, G4473, G4474, G4475, G4476, G4477, G4478, G4479, G4480, G4481,
         G4482, G4483, G4484, G4485, G4486, G4487, G4488, G4489, G4490, G4491,
         G4492, G4493, G4494, G4495, G4496, G4497, G4498, G4499, G4500, G4501,
         G4502, G4503, G4805, G4806, G4807, G4808, G4809, G4810, G4811, G4812,
         G4813, G4814, G4815, G4816, G4817, G4818, G4819, G4820, G4821, G4822,
         G4823, G4824, G4825, G4826, G4827, G4828, G4829, G4830, G4831, G4832,
         G4833, G4834, G4835, G4836, G4504, G4505, G4506, G4507, G4508, G4509,
         G4510, G4511, G4512, G4513, G4514, G4515, G4516, G4517, G4518, G4519,
         G4520, G4521, G4522, G4523, G4524, G4525, G4526, G4527, G4528, G4529,
         G4530, G4531, G4532, G4533, G4389, G4388, G4591, G7318, G7319, G7320,
         G7321, G7322, G7323, G7324, G7325, G7326, G7327, G7328, G7329, G7330,
         G7331, G7332, G7333, G7334, G7335, G7336, G7337, G7338, G7339, G7340,
         G7341, G7342, G7343, G7344, G7345, G7346, G7347, G7348, G7349, G7660,
         G7661, G7350, G7351, G7352, G7353, G7354, G7355, G7356, G7357, G7358,
         G7359, G7360, G7361, G7362, G7363, G7364, G7365, G7366, G7367, G7368,
         G7369, G7370, G7371, G7372, G7373, G7374, G7375, G7376, G7377, G7378,
         G7379, G7380, G7381, G7382, G7383, G7384, G7385, G7386, G7387, G7388,
         G7389, G7390, G7391, G7392, G7393, G7394, G7395, G7396, G7397, G7398,
         G7399, G7400, G7401, G7402, G7403, G7404, G7405, G7406, G7407, G7408,
         G7409, G7410, G7411, G7412, G7413, G7414, G7415, G7416, G7417, G7418,
         G7419, G7420, G7421, G7422, G7423, G7424, G7425, G7426, G7427, G7428,
         G7429, G7430, G7431, G7432, G7433, G7434, G7435, G7436, G7437, G7438,
         G7439, G7440, G7441, G7442, G7443, G7444, G7445, G7446, G7447, G7448,
         G7449, G7450, G7451, G7452, G7453, G7454, G7455, G7456, G7457, G7458,
         G7459, G7460, G7461, G7462, G7463, G7464, G7465, G7466, G7467, G7468,
         G7469, G7470, G7471, G7472, G7473, G7474, G7475, G7476, G7477, G7478,
         G7479, G7480, G7481, G7482, G7483, G7484, G7485, G7486, G7487, G7488,
         G7489, G7490, G7491, G7492, G7493, G7494, G7495, G7689, G7690, G7691,
         G7692, G7693, G7694, G7695, G7696, G7697, G7698, G7699, G7700, G7701,
         G7702, G7703, G7704, G7705, G7706, G7707, G7708, G7709, G7710, G7711,
         G7712, G7713, G7714, G7715, G7716, G7717, G7718, G7719, G7720, G7496,
         G7497, G7498, G7499, G7500, G7501, G7502, G7503, G7504, G7505, G7506,
         G7507, G7508, G7509, G7510, G7511, G7512, G7513, G7514, G7515, G7516,
         G7517, G7518, G7519, G7520, G7521, G7522, G7523, G7524, G7525, G7317,
         G7316, G7605;
  wire   n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847;
  nor U13198(n17852,n15634,n17877);
  nor U13199(n21669,n15649,n21691);
  nor U13200(n17851,n15649,n17877);
  nor U13201(n19456,n15634,G36460);
  nor U13202(n19459,n15649,G36460);
  nor U13203(n21670,n15634,n21691);
  nor U13204(n23061,n15649,G36215);
  nor U13205(n23058,n15634,G36215);
  nand U13206(n17109,n17015,n17438);
  not U13207(n15649,n15634);
  nand U13208(n15634,n23544,n23545);
  not U13209(n17937,n17085);
  nand U13210(n17085,n17304,n16674);
  nand U13211(n17882,n19387,n19388);
  nand U13212(n20838,n21229,n21230);
  not U13213(n16290,n16298);
  nand U13214(n16298,n16676,n16286);
  nand U13215(n13339,n13652,n12952,n13653,n13635);
  or U13216(n22110,n22106,n22105);
  and U13217(n20839,n20843,n21231);
  nand U13218(n15281,n14579,n12521);
  nand U13219(n14460,n14319,n12527);
  nand U13220(n16936,n16704,n16533);
  nand U13221(n20539,n20311,n20142);
  nand U13222(n14230,n14042,n12894);
  nand U13223(n21697,n22992,n22993);
  nand U13224(n14527,n15551,n15552);
  nand U13225(n14528,n15556,n15557);
  nand U13226(n17883,n19392,n19393);
  nand U13227(n21698,n22997,n22998);
  nand U13228(n13344,n13654,n13655);
  nand U13229(n22847,n20251,n21788,n22851);
  nand U13230(n22795,n20239,n21788,n22799);
  nand U13231(n22754,n20227,n21788,n22758);
  nand U13232(n22710,n20215,n21788,n22714);
  nand U13233(n22665,n20203,n21788,n22669);
  nand U13234(n19904,n20269,n20270);
  and U13235(n17108,n17424,n17114);
  nand U13236(n20846,n21223,n21248,n21229);
  nand U13237(n17843,n16677,n19401);
  nand U13238(n22944,n22106,G36101);
  nand U13239(n22883,n22106,G36102);
  nand U13240(n22869,n22106,G36103);
  nand U13241(n22824,n22106,G36104);
  nand U13242(n22779,n22106,G36105);
  nand U13243(n22731,n22106,G36106);
  nor U13244(n14514,n13653,n14517);
  not U13245(n19800,n19798);
  nor U13246(n19798,n19894,n19895);
  not U13247(n16093,G4591);
  nor U13248(G4591,n17829,G4389);
  nand U13249(n16935,n16705,n16535);
  nand U13250(n20538,n20312,n20144);
  nand U13251(n14238,n14053,n12524);
  nand U13252(n19087,n17974,n16172);
  nand U13253(n19037,n17974,n16169);
  nand U13254(n14479,n14320,n13133);
  nand U13255(n14473,n14320,n12786);
  nand U13256(n14467,n14320,n12748);
  nand U13257(n15402,n14591,n12533);
  nand U13258(n15366,n14591,n12530);
  nand U13259(n15328,n14591,n12527);
  nand U13260(n15393,n14545,n13133);
  nand U13261(n15357,n14545,n12786);
  nand U13262(n15319,n14545,n12748);
  nand U13263(n15388,n14583,n14246);
  nand U13264(n15352,n14583,n14237);
  nand U13265(n15314,n14583,n14228);
  nand U13266(n15240,n14583,n15241);
  nand U13267(n14529,n15561,n15562);
  nand U13268(n17881,n19397,n19398);
  nand U13269(n21696,n23002,n23003);
  nand U13270(n16294,n16663,n16664);
  not U13271(G4389,G36460);
  not U13272(n16190,n16192);
  nand U13273(n16192,n16286,n16287);
  not U13274(G1625,n19677);
  nand U13275(n19677,n21335,G36215);
  nand U13276(n19783,n20282,n23006);
  not U13277(n13028,n12970);
  nand U13278(n12970,n13325,n13326);
  not U13279(n17976,n17914);
  nand U13280(n13340,n13641,n13642,n13648);
  not U13281(n13648,n13344);
  not U13282(n14023,n14029);
  nand U13283(n20843,n20269,n21197,n21232);
  nand U13284(n17114,n17440,n17426);
  not U13285(n15631,n15823);
  nand U13286(n14516,n13660,n13903);
  not U13287(n13903,n13661);
  nand U13288(n22104,n22105,G36088);
  nand U13289(n22146,n22105,G36087);
  nand U13290(n22189,n22105,G36086);
  nand U13291(n22238,n22105,G36085);
  nand U13292(n22280,n22105,G36084);
  nand U13293(n22325,n22105,G36083);
  nand U13294(n22368,n22105,G36082);
  not U13295(n19458,n19544);
  and U13296(n19778,n19771,n19782);
  nand U13297(n21760,n19782,n19690);
  nand U13298(n21802,n19782,n19693);
  nand U13299(n21839,n19782,n19696);
  nand U13300(n21877,n19782,n19699);
  nand U13301(n21911,n19782,n19702);
  nand U13302(n21946,n19782,n19705);
  nand U13303(n21985,n19782,n19708);
  nand U13304(n22019,n19782,n19711);
  nand U13305(n22057,n19782,n19714);
  nand U13306(n22090,n19782,n19717);
  nand U13307(n22134,n19782,n19720);
  not U13308(n19159,n17929);
  nand U13309(n17885,n17929,n17930);
  nand U13310(n17949,n17929,n16779);
  nand U13311(n17995,n17929,n18034);
  nand U13312(n18036,n17929,n18076);
  nand U13313(n18078,n17929,n16832);
  nand U13314(n18116,n17929,n18153);
  nand U13315(n18155,n17929,n18195);
  nand U13316(n18197,n17929,n16933);
  nand U13317(n18234,n17929,n16810);
  nand U13318(n18274,n17929,n18311);
  nand U13319(n18313,n17929,n18366);
  nand U13320(n17948,n17993,n16106);
  nand U13321(n17994,n17993,n16109);
  nand U13322(n18035,n17993,n16112);
  nand U13323(n18077,n17993,n16115);
  nand U13324(n18115,n17993,n16118);
  nand U13325(n18154,n17993,n16121);
  nand U13326(n18196,n17993,n16124);
  nand U13327(n18233,n17993,n16127);
  nand U13328(n18273,n17993,n16130);
  nand U13329(n18312,n17993,n16133);
  nand U13330(n18367,n17993,n16136);
  nand U13331(n18422,n17993,n16139);
  not U13332(n23060,n23301);
  nor U13333(n14310,n14311,n13653);
  nor U13334(n20844,n21230,n21240);
  not U13335(n19906,n19898);
  nor U13336(n19898,n19895,n20279);
  not U13337(n12448,G7605);
  nor U13338(G7605,n14017,G7317);
  nand U13339(n17973,n17924,n17921,n17923);
  nand U13340(n21787,n21747,n21753,n20625);
  not U13341(n21773,n22948);
  nor U13342(n22948,n21725,n21724);
  nand U13343(n14590,n14556,n14558);
  not U13344(G7317,G36705);
  or U13345(G793,G36707,n12444);
  xnor U13346(n12444,G36462,G36217);
  or U13347(G792,G36706,n12445);
  xnor U13348(n12445,G36216,G36461);
  nand U13349(G7720,n12446,n12447);
  nand U13350(n12447,G36674,n12448);
  nand U13351(n12446,G7605,n12449);
  nand U13352(G7719,n12450,n12451);
  nand U13353(n12451,G36673,n12448);
  nand U13354(n12450,G7605,n12452);
  nand U13355(G7718,n12453,n12454);
  nand U13356(n12454,G36672,n12448);
  nand U13357(n12453,G7605,n12455);
  nand U13358(G7717,n12456,n12457);
  nand U13359(n12457,G36671,n12448);
  nand U13360(n12456,G7605,n12458);
  nand U13361(G7716,n12459,n12460);
  nand U13362(n12460,G36670,n12448);
  nand U13363(n12459,G7605,n12461);
  nand U13364(G7715,n12462,n12463);
  nand U13365(n12463,G36669,n12448);
  nand U13366(n12462,G7605,n12464);
  nand U13367(G7714,n12465,n12466);
  nand U13368(n12466,G36668,n12448);
  nand U13369(n12465,G7605,n12467);
  nand U13370(G7713,n12468,n12469);
  nand U13371(n12469,G36667,n12448);
  nand U13372(n12468,G7605,n12470);
  nand U13373(G7712,n12471,n12472);
  nand U13374(n12472,G36666,n12448);
  nand U13375(n12471,G7605,n12473);
  nand U13376(G7711,n12474,n12475);
  nand U13377(n12475,G36665,n12448);
  nand U13378(n12474,G7605,n12476);
  nand U13379(G7710,n12477,n12478);
  nand U13380(n12478,G36664,n12448);
  nand U13381(n12477,G7605,n12479);
  nand U13382(G7709,n12480,n12481);
  nand U13383(n12481,G36663,n12448);
  nand U13384(n12480,G7605,n12482);
  nand U13385(G7708,n12483,n12484);
  nand U13386(n12484,G36662,n12448);
  nand U13387(n12483,G7605,n12485);
  nand U13388(G7707,n12486,n12487);
  nand U13389(n12487,G36661,n12448);
  nand U13390(n12486,G7605,n12488);
  nand U13391(G7706,n12489,n12490);
  nand U13392(n12490,G36660,n12448);
  nand U13393(n12489,G7605,n12491);
  nand U13394(G7705,n12492,n12493);
  nand U13395(n12493,G36659,n12448);
  nand U13396(n12492,G7605,n12494);
  nand U13397(G7704,n12495,n12496);
  nand U13398(n12496,G36658,n12448);
  nand U13399(n12495,G7605,n12497);
  nand U13400(G7703,n12498,n12499);
  nand U13401(n12499,G36657,n12448);
  nand U13402(n12498,G7605,n12500);
  nand U13403(G7702,n12501,n12502);
  nand U13404(n12502,G36656,n12448);
  nand U13405(n12501,G7605,n12503);
  nand U13406(G7701,n12504,n12505);
  nand U13407(n12505,G36655,n12448);
  nand U13408(n12504,G7605,n12506);
  nand U13409(G7700,n12507,n12508);
  nand U13410(n12508,G36654,n12448);
  nand U13411(n12507,G7605,n12509);
  nand U13412(G7699,n12510,n12511);
  nand U13413(n12511,G36653,n12448);
  nand U13414(n12510,G7605,n12512);
  nand U13415(G7698,n12513,n12514);
  nand U13416(n12514,G36652,n12448);
  nand U13417(n12513,G7605,n12515);
  nand U13418(G7697,n12516,n12517);
  nand U13419(n12517,G36651,n12448);
  nand U13420(n12516,G7605,n12518);
  nand U13421(G7696,n12519,n12520);
  nand U13422(n12520,G36650,n12448);
  nand U13423(n12519,G7605,n12521);
  nand U13424(G7695,n12522,n12523);
  nand U13425(n12523,G36649,n12448);
  nand U13426(n12522,G7605,n12524);
  nand U13427(G7694,n12525,n12526);
  nand U13428(n12526,G36648,n12448);
  nand U13429(n12525,G7605,n12527);
  nand U13430(G7693,n12528,n12529);
  nand U13431(n12529,G36647,n12448);
  nand U13432(n12528,G7605,n12530);
  nand U13433(G7692,n12531,n12532);
  nand U13434(n12532,G36646,n12448);
  nand U13435(n12531,G7605,n12533);
  nand U13436(G7691,n12534,n12535);
  nand U13437(n12535,G36645,n12448);
  nand U13438(n12534,G7605,n12536);
  nand U13439(G7690,n12537,n12538);
  nand U13440(n12538,G36644,n12448);
  nand U13441(n12537,G7605,n12539);
  nand U13442(G7689,n12540,n12541);
  nand U13443(n12541,G36643,n12448);
  nand U13444(n12540,G7605,n12542);
  nand U13445(G7661,n12543,n12544);
  nand U13446(n12544,G36496,n12545);
  nand U13447(n12543,n12546,n12547);
  nand U13448(G7660,n12548,n12549);
  nand U13449(n12549,G36495,n12545);
  nand U13450(n12548,n12546,n12550);
  nand U13451(G7525,n12551,n12552,n12553,n12554);
  nor U13452(n12554,n12555,n12556,n12557,n12558);
  nor U13453(n12558,n12559,n12560);
  nor U13454(n12557,n12561,n12562);
  nor U13455(n12556,n12563,n12564);
  nor U13456(n12555,n12565,n12566);
  nand U13457(n12552,n12567,n12568);
  nand U13458(n12551,n12569,n12570);
  nand U13459(G7524,n12571,n12572,n12573,n12574);
  nor U13460(n12574,n12575,n12576,n12577);
  nor U13461(n12577,n12564,n12578);
  nor U13462(n12576,n12579,n12580);
  nor U13463(n12575,n12581,n12562);
  nand U13464(n12573,G36703,G7317);
  nand U13465(n12572,n12582,n12464);
  nand U13466(n12571,n12583,n12567);
  nand U13467(G7523,n12584,n12585,n12586,n12587);
  nor U13468(n12587,n12588,n12589,n12590,n12591);
  nor U13469(n12591,n12592,n12560);
  nor U13470(n12590,n12593,n12562);
  nor U13471(n12589,n12564,n12594);
  nor U13472(n12588,n12595,n12566);
  nand U13473(n12585,n12596,n12567);
  nand U13474(n12584,n12597,n12569);
  nand U13475(G7522,n12598,n12599,n12600,n12601);
  nor U13476(n12601,n12602,n12603,n12604);
  nor U13477(n12604,n12564,n12605);
  nor U13478(n12603,n12579,n12606);
  nor U13479(n12602,n12607,n12562);
  nand U13480(n12600,G36701,G7317);
  nand U13481(n12599,n12582,n12476);
  nand U13482(n12598,n12608,n12567);
  nand U13483(G7521,n12609,n12610,n12611,n12612);
  nor U13484(n12612,n12613,n12614,n12615,n12616);
  nor U13485(n12616,n12617,n12560);
  nor U13486(n12615,n12618,n12562);
  nor U13487(n12614,n12564,n12619);
  not U13488(n12619,n12620);
  and U13489(n12613,n12621,n12622);
  nand U13490(n12611,G36700,G7317);
  nand U13491(n12610,n12567,n12623);
  nand U13492(n12609,n12624,n12569);
  nand U13493(G7520,n12625,n12626,n12627,n12628);
  nor U13494(n12628,n12629,n12630,n12631,n12632);
  nor U13495(n12632,n12633,n12634);
  nor U13496(n12631,n12635,n12636);
  nor U13497(n12630,G36699,n12564);
  nor U13498(n12629,G36705,n12637);
  nand U13499(n12627,n12582,n12536);
  nand U13500(n12626,n12622,n12638);
  or U13501(n12625,n12562,n12639);
  nand U13502(G7519,n12640,n12641,n12642,n12643);
  nor U13503(n12643,n12644,n12645,n12646,n12647);
  nor U13504(n12647,n12648,n12560);
  nor U13505(n12646,n12649,n12562);
  nor U13506(n12645,n12564,n12650);
  nor U13507(n12644,n12651,n12566);
  nand U13508(n12641,n12652,n12567);
  nand U13509(n12640,n12653,n12569);
  nand U13510(G7518,n12654,n12655,n12656,n12657);
  nor U13511(n12657,n12658,n12659,n12660);
  nor U13512(n12660,n12564,n12661);
  nor U13513(n12659,n12579,n12662);
  nor U13514(n12658,n12663,n12562);
  nand U13515(n12656,G36697,G7317);
  nand U13516(n12655,n12582,n12461);
  nand U13517(n12654,n12664,n12567);
  nand U13518(G7517,n12665,n12666,n12667,n12668);
  nor U13519(n12668,n12669,n12670,n12671,n12672);
  nor U13520(n12672,n12673,n12560);
  nor U13521(n12671,n12617,n12562);
  nor U13522(n12670,n12564,n12674);
  nor U13523(n12669,n12675,n12566);
  nand U13524(n12666,n12676,n12567);
  nand U13525(n12665,n12677,n12569);
  nand U13526(G7516,n12678,n12679,n12680,n12681);
  nor U13527(n12681,n12682,n12683,n12684);
  nor U13528(n12684,n12685,n12566);
  nor U13529(n12683,n12686,n12687);
  nor U13530(n12682,n12688,n12562);
  nand U13531(n12680,n12569,n12689);
  nand U13532(n12679,n12582,n12542);
  nand U13533(n12678,n12690,n12567);
  nand U13534(G7515,n12691,n12692,n12693,n12694);
  nor U13535(n12694,n12695,n12696,n12697);
  nor U13536(n12697,n12564,n12698);
  nor U13537(n12696,n12579,n12699);
  nor U13538(n12695,n12700,n12562);
  nand U13539(n12693,G36694,G7317);
  nand U13540(n12692,n12582,n12482);
  nand U13541(n12691,n12701,n12567);
  nand U13542(G7514,n12702,n12703,n12704,n12705);
  nor U13543(n12705,n12706,n12707,n12708,n12709);
  nor U13544(n12709,n12618,n12560);
  nor U13545(n12708,n12592,n12562);
  nor U13546(n12707,n12564,n12710);
  nor U13547(n12706,n12711,n12566);
  nand U13548(n12703,n12712,n12567);
  nand U13549(n12702,n12713,n12569);
  nand U13550(G7513,n12714,n12715,n12716,n12717);
  nor U13551(n12717,n12718,n12719,n12720);
  nor U13552(n12720,n12564,n12721);
  nor U13553(n12719,n12579,n12722);
  nor U13554(n12718,n12723,n12562);
  nand U13555(n12716,G36692,G7317);
  nand U13556(n12715,n12582,n12470);
  nand U13557(n12714,n12724,n12567);
  nand U13558(G7512,n12725,n12726,n12727,n12728);
  nor U13559(n12728,n12729,n12730,n12731,n12732);
  nor U13560(n12732,n12593,n12560);
  nor U13561(n12731,n12733,n12562);
  nor U13562(n12730,n12564,n12734);
  nor U13563(n12729,n12735,n12566);
  nand U13564(n12726,n12736,n12567);
  nand U13565(n12725,n12737,n12569);
  nand U13566(G7511,n12738,n12739,n12740,n12741);
  nor U13567(n12741,n12742,n12743,n12744,n12745);
  nor U13568(n12745,n12639,n12560);
  nor U13569(n12744,n12559,n12562);
  nor U13570(n12743,n12564,n12746);
  nor U13571(n12742,n12747,n12566);
  nand U13572(n12739,n12748,n12567);
  nand U13573(n12738,n12569,n12749);
  nand U13574(G7510,n12750,n12751,n12752,n12753);
  nor U13575(n12753,n12754,n12755,n12756,n12757);
  nor U13576(n12757,n12758,n12560);
  nor U13577(n12756,n12648,n12562);
  nor U13578(n12755,n12759,n12564);
  nor U13579(n12754,n12760,n12566);
  nand U13580(n12751,n12761,n12567);
  nand U13581(n12750,n12762,n12569);
  nand U13582(G7509,n12763,n12764,n12765,n12766);
  nor U13583(n12766,n12767,n12768,n12769);
  nor U13584(n12769,n12564,n12770);
  nor U13585(n12768,n12579,n12771);
  nor U13586(n12767,n12772,n12562);
  nand U13587(n12765,G36688,G7317);
  nand U13588(n12764,n12582,n12473);
  nand U13589(n12763,n12773,n12567);
  nand U13590(G7508,n12774,n12775,n12776,n12777);
  nor U13591(n12777,n12778,n12779,n12780,n12781);
  nor U13592(n12781,n12782,n12560);
  nor U13593(n12780,n12783,n12562);
  nor U13594(n12779,n12564,n12784);
  nor U13595(n12778,n12785,n12566);
  nand U13596(n12775,n12786,n12567);
  nand U13597(n12774,n12569,n12787);
  nand U13598(G7507,n12788,n12789,n12790,n12791);
  nor U13599(n12791,n12792,n12793,n12794,n12795);
  nor U13600(n12795,n12561,n12560);
  nor U13601(n12794,n12796,n12562);
  nor U13602(n12793,n12564,n12797);
  nor U13603(n12792,n12798,n12566);
  nand U13604(n12789,n12799,n12567);
  nand U13605(n12788,n12800,n12569);
  nand U13606(G7506,n12801,n12802,n12803);
  nor U13607(n12803,n12804,n12805,n12806);
  nor U13608(n12806,n12807,n12566);
  nor U13609(n12805,n12686,n12808);
  nor U13610(n12804,n12809,n12562);
  nand U13611(n12802,n12810,n12567);
  nand U13612(n12801,n12569,n12811);
  nand U13613(G7505,n12812,n12813,n12814,n12815);
  nor U13614(n12815,n12816,n12817,n12818);
  nor U13615(n12818,n12564,n12819);
  nor U13616(n12817,n12579,n12820);
  nor U13617(n12816,n12821,n12562);
  nand U13618(n12814,G36684,G7317);
  nand U13619(n12813,n12582,n12485);
  nand U13620(n12812,n12822,n12567);
  nand U13621(G7504,n12823,n12824,n12825,n12826);
  nor U13622(n12826,n12827,n12828,n12829,n12830);
  nor U13623(n12830,n12831,n12560);
  nor U13624(n12829,n12832,n12562);
  nor U13625(n12828,n12564,n12833);
  nor U13626(n12827,n12834,n12566);
  nand U13627(n12824,n12835,n12567);
  nand U13628(n12823,n12836,n12569);
  nand U13629(G7503,n12837,n12838,n12839,n12840);
  nor U13630(n12840,n12841,n12842,n12843);
  nor U13631(n12843,n12564,n12844);
  nor U13632(n12842,n12579,n12845);
  nor U13633(n12841,n12846,n12562);
  nand U13634(n12839,G36682,G7317);
  nand U13635(n12838,n12582,n12479);
  nand U13636(n12837,n12847,n12567);
  nand U13637(G7502,n12848,n12849,n12850,n12851);
  nor U13638(n12851,n12852,n12853,n12854,n12855);
  nor U13639(n12855,n12796,n12560);
  nor U13640(n12854,n12831,n12562);
  nor U13641(n12853,n12564,n12856);
  nor U13642(n12852,n12857,n12566);
  nand U13643(n12849,n12858,n12567);
  nand U13644(n12848,n12859,n12569);
  nand U13645(G7501,n12860,n12861,n12862,n12863);
  nor U13646(n12863,n12864,n12865,n12866);
  nor U13647(n12866,n12867,n12566);
  nor U13648(n12865,n12686,n12868);
  and U13649(n12686,n12564,G36705);
  nor U13650(n12864,n12782,n12562);
  nand U13651(n12862,n12569,n12869);
  nand U13652(n12861,n12582,n12539);
  nand U13653(n12860,n12870,n12567);
  nand U13654(G7500,n12871,n12872,n12873,n12874);
  nor U13655(n12874,n12875,n12876,n12877,n12878);
  nor U13656(n12878,n12733,n12560);
  nor U13657(n12877,n12879,n12562);
  nor U13658(n12876,n12564,n12880);
  nor U13659(n12875,n12881,n12566);
  nand U13660(n12872,n12882,n12567);
  nand U13661(n12871,n12883,n12569);
  nand U13662(G7499,n12884,n12885,n12886,n12887);
  nor U13663(n12887,n12888,n12889,n12890,n12891);
  nor U13664(n12891,n12783,n12560);
  nor U13665(n12890,n12673,n12562);
  nor U13666(n12889,n12564,n12892);
  nor U13667(n12888,n12893,n12566);
  nand U13668(n12885,n12894,n12567);
  nand U13669(n12884,n12569,n12895);
  nand U13670(G7498,n12896,n12897,n12898,n12899);
  nor U13671(n12899,n12900,n12901,n12902);
  nor U13672(n12902,n12564,n12903);
  nor U13673(n12901,n12579,n12904);
  nor U13674(n12579,n12569,n12622);
  not U13675(n12622,n12566);
  nor U13676(n12900,n12905,n12562);
  nand U13677(n12898,G36677,G7317);
  nand U13678(n12897,n12582,n12467);
  not U13679(n12582,n12560);
  nand U13680(n12896,n12906,n12567);
  nand U13681(G7497,n12907,n12908,n12909,n12910);
  nor U13682(n12910,n12911,n12912,n12913,n12914);
  nor U13683(n12914,n12832,n12560);
  nand U13684(n12560,n12915,n12916,n12917);
  nor U13685(n12913,n12758,n12562);
  nand U13686(n12562,n12915,n12918,n12917);
  nor U13687(n12912,n12564,n12919);
  and U13688(n12564,n12920,n12921,n12922,n12448);
  nand U13689(n12921,n12923,n12924);
  nand U13690(n12924,n12925,n12926,n12927);
  nand U13691(n12927,n12928,n12929);
  nand U13692(n12926,n12930,n12931);
  or U13693(n12930,n12932,n12933);
  nand U13694(n12925,n12934,n12935);
  nand U13695(n12920,n12915,n12929);
  nor U13696(n12911,n12936,n12566);
  nand U13697(n12566,n12923,n12933,n12937);
  nand U13698(n12908,n12938,n12567);
  not U13699(n12567,n12635);
  nand U13700(n12635,n12923,n12939);
  nand U13701(n12939,n12940,n12941);
  nand U13702(n12941,n12917,n12928);
  nand U13703(n12940,n12937,n12932);
  nand U13704(n12932,n12942,n12943,n12944,n12945);
  nand U13705(n12945,n12946,n12947);
  or U13706(n12947,n12948,n12949);
  nand U13707(n12944,n12950,n12951);
  or U13708(n12943,n12952,n12953);
  nand U13709(n12907,n12954,n12569);
  not U13710(n12569,n12634);
  nand U13711(G7496,n12955,n12956);
  nand U13712(n12956,n12957,n12958);
  nand U13713(n12958,n12959,n12960,n12961,n12962);
  nand U13714(n12962,n12928,n12963);
  nor U13715(n12961,n12964,n12965);
  nor U13716(n12965,n12966,n12950);
  nor U13717(n12966,n12967,n12968);
  nor U13718(n12968,n12969,n12970);
  and U13719(n12967,n12963,n12951);
  nor U13720(n12964,n12971,n12972,n12973);
  nor U13721(n12973,n12974,n12975,n12976,n12977);
  nor U13722(n12977,n12950,n12963);
  nand U13723(n12963,n12978,n12979,n12980,n12981);
  nor U13724(n12981,n12982,n12983,n12984,n12985);
  nand U13725(n12985,n12986,n12987,n12988,n12989);
  not U13726(n12989,n12990);
  or U13727(n12984,n12991,n12992,n12993,n12994);
  or U13728(n12983,n12995,n12996,n12997,n12998);
  or U13729(n12982,n12999,n13000,n13001,n13002);
  nor U13730(n12980,n13003,n13004,n13005,n13006);
  xor U13731(n13006,n12542,n12811);
  xor U13732(n13005,n13007,n12452);
  nand U13733(n13004,n13008,n13009,n13010);
  xor U13734(n13010,n12449,n13011);
  nand U13735(n13008,n12663,n13012);
  or U13736(n13003,n13013,n13014,n13015,n13016);
  nor U13737(n12979,n13017,n13018,n13019,n13020);
  nor U13738(n12978,n13021,n13022,n13023,n13024);
  nor U13739(n12976,n13025,n13026,n13027);
  nor U13740(n12975,n13028,n13029);
  nor U13741(n12972,n12953,n13030);
  xor U13742(n13030,n12970,n12950);
  nand U13743(n12960,n13031,n13027);
  nand U13744(n13027,n13032,n13033);
  or U13745(n13033,n13034,n13011);
  nand U13746(n13032,n13035,n13036);
  nand U13747(n13036,n13037,n13038);
  nand U13748(n13038,n13039,n13040,n13041);
  nand U13749(n13041,n13007,n13042);
  nand U13750(n13040,n13043,n13044,n13045);
  nand U13751(n13045,n13046,n13047,n13048);
  nand U13752(n13048,n13049,n13050,n13051);
  nand U13753(n13051,n13052,n13053,n13054);
  nand U13754(n13054,n13055,n13056,n13057);
  nand U13755(n13057,n13058,n13059,n13060);
  nand U13756(n13060,n13061,n13062,n13063);
  nand U13757(n13063,n13064,n13065,n13066);
  nand U13758(n13066,n13067,n13068,n13069);
  nand U13759(n13069,n13070,n13071,n13072);
  nand U13760(n13072,n13073,n13074,n13075);
  nand U13761(n13075,n13076,n13077,n13078);
  nand U13762(n13078,n13079,n13080,n13081);
  nand U13763(n13081,n13082,n13083,n13084);
  nand U13764(n13084,n13085,n13086,n13087);
  nand U13765(n13087,n13088,n13089,n13090);
  nand U13766(n13090,n13091,n13092,n13093);
  nand U13767(n13093,n13094,n13095,n13096);
  nand U13768(n13096,n13097,n13098,n13099);
  nand U13769(n13099,n13100,n13101,n13102);
  nand U13770(n13102,n13103,n13104,n13105);
  nand U13771(n13105,n13106,n13107,n13108);
  nand U13772(n13108,n13109,n13110,n13111);
  nand U13773(n13111,n13112,n13113,n13114);
  nand U13774(n13114,n13115,n13116,n13117,n13118);
  nand U13775(n13118,n13119,n13120,n13121,n12970);
  nand U13776(n13121,n13122,n13123,n13124);
  nand U13777(n13124,n12870,n13125);
  nand U13778(n13123,n13126,n13127,n13128);
  nand U13779(n13128,n13129,n12689);
  nand U13780(n13127,n12811,n13130,n13131);
  not U13781(n13131,n12810);
  nand U13782(n13130,n13132,n12690);
  or U13783(n13126,n13125,n12870);
  nand U13784(n13122,n13133,n12633);
  or U13785(n13120,n13134,n12786);
  nand U13786(n13119,n13135,n12636);
  not U13787(n12636,n13133);
  nand U13788(n13117,n12987,n13136,n13028);
  nand U13789(n13136,n12986,n13137);
  nand U13790(n13137,n12988,n13138);
  nand U13791(n13138,n12811,n13009,n13139);
  nand U13792(n13009,n13132,n12539);
  not U13793(n13132,n12689);
  and U13794(n12988,n13140,n13141);
  nand U13795(n13141,n12688,n12869);
  nand U13796(n13140,n12809,n12689);
  and U13797(n12986,n13142,n13143);
  nand U13798(n13143,n12633,n12533);
  nand U13799(n13142,n13125,n12536);
  and U13800(n12987,n13144,n13145);
  nand U13801(n13145,n12639,n12787);
  nand U13802(n13144,n12782,n13135);
  nand U13803(n13116,n13028,n12990);
  nand U13804(n12990,n13146,n13147);
  nand U13805(n13147,n13148,n12527);
  nand U13806(n13146,n13134,n12530);
  nand U13807(n13115,n13149,n12970);
  nand U13808(n13149,n13150,n13151);
  nand U13809(n13151,n12748,n13148);
  nand U13810(n13150,n12786,n13134);
  nand U13811(n13113,n13028,n12991);
  nand U13812(n12991,n13152,n13153);
  nand U13813(n13153,n12559,n12895);
  nand U13814(n13152,n12783,n12749);
  nand U13815(n13112,n13154,n12970);
  nand U13816(n13154,n13155,n13156);
  or U13817(n13156,n13157,n12894);
  or U13818(n13155,n13148,n12748);
  nand U13819(n13110,n13028,n12992);
  nand U13820(n12992,n13158,n13159);
  nand U13821(n13159,n13160,n12521);
  nand U13822(n13158,n13157,n12524);
  nand U13823(n13109,n13161,n12970);
  nand U13824(n13161,n13162,n13163);
  nand U13825(n13163,n12568,n13160);
  nand U13826(n13162,n12894,n13157);
  nand U13827(n13107,n13028,n12993);
  nand U13828(n12993,n13164,n13165);
  nand U13829(n13165,n12561,n12677);
  nand U13830(n13164,n12673,n12570);
  nand U13831(n13106,n13166,n12970);
  nand U13832(n13166,n13167,n13168);
  or U13833(n13168,n13169,n12676);
  or U13834(n13167,n13160,n12568);
  nand U13835(n13104,n13028,n12994);
  nand U13836(n12994,n13170,n13171);
  nand U13837(n13171,n13172,n12515);
  nand U13838(n13170,n13169,n12518);
  nand U13839(n13103,n13173,n12970);
  nand U13840(n13173,n13174,n13175);
  nand U13841(n13175,n12799,n13172);
  nand U13842(n13174,n12676,n13169);
  nand U13843(n13101,n13028,n12995);
  nand U13844(n12995,n13176,n13177);
  nand U13845(n13177,n12796,n12624);
  nand U13846(n13176,n12617,n12800);
  nand U13847(n13100,n13178,n12970);
  nand U13848(n13178,n13179,n13180);
  nand U13849(n13180,n13181,n12624);
  or U13850(n13179,n13172,n12799);
  nand U13851(n13098,n13028,n12996);
  nand U13852(n12996,n13182,n13183);
  nand U13853(n13183,n13184,n12509);
  nand U13854(n13182,n13185,n12512);
  nand U13855(n13097,n13186,n12970);
  nand U13856(n13186,n13187,n13188);
  nand U13857(n13188,n12858,n13184);
  nand U13858(n13187,n13185,n12623);
  nand U13859(n13095,n13028,n12997);
  nand U13860(n12997,n13189,n13190);
  nand U13861(n13190,n12831,n12713);
  nand U13862(n13189,n12618,n12859);
  nand U13863(n13094,n13191,n12970);
  nand U13864(n13191,n13192,n13193);
  or U13865(n13193,n13194,n12712);
  or U13866(n13192,n13184,n12858);
  nand U13867(n13092,n13028,n12998);
  nand U13868(n12998,n13195,n13196);
  nand U13869(n13196,n13197,n12503);
  nand U13870(n13195,n13194,n12506);
  nand U13871(n13091,n13198,n12970);
  nand U13872(n13198,n13199,n13200);
  nand U13873(n13200,n12835,n13197);
  nand U13874(n13199,n12712,n13194);
  nand U13875(n13089,n13028,n12999);
  nand U13876(n12999,n13201,n13202);
  nand U13877(n13202,n12832,n12597);
  nand U13878(n13201,n12592,n12836);
  nand U13879(n13088,n13203,n12970);
  nand U13880(n13203,n13204,n13205);
  or U13881(n13205,n13206,n12596);
  or U13882(n13204,n13197,n12835);
  nand U13883(n13086,n13028,n13000);
  nand U13884(n13000,n13207,n13208);
  nand U13885(n13208,n13209,n12497);
  nand U13886(n13207,n13206,n12500);
  nand U13887(n13085,n13210,n12970);
  nand U13888(n13210,n13211,n13212);
  nand U13889(n13212,n12938,n13209);
  nand U13890(n13211,n12596,n13206);
  nand U13891(n13083,n13028,n13001);
  nand U13892(n13001,n13213,n13214);
  nand U13893(n13214,n12758,n12737);
  nand U13894(n13213,n12593,n12954);
  nand U13895(n13082,n13215,n12970);
  nand U13896(n13215,n13216,n13217);
  or U13897(n13217,n13218,n12736);
  or U13898(n13216,n13209,n12938);
  nand U13899(n13080,n13028,n13002);
  nand U13900(n13002,n13219,n13220);
  nand U13901(n13220,n13221,n12491);
  nand U13902(n13219,n13218,n12494);
  nand U13903(n13079,n13222,n12970);
  nand U13904(n13222,n13223,n13224);
  nand U13905(n13224,n12761,n13221);
  nand U13906(n13223,n12736,n13218);
  nand U13907(n13077,n13028,n13024);
  nand U13908(n13024,n13225,n13226);
  nand U13909(n13226,n12648,n12883);
  nand U13910(n13225,n12733,n12762);
  nand U13911(n13076,n13227,n12970);
  nand U13912(n13227,n13228,n13229);
  or U13913(n13229,n13230,n12882);
  or U13914(n13228,n13221,n12761);
  nand U13915(n13074,n13028,n13023);
  nand U13916(n13023,n13231,n13232);
  nand U13917(n13232,n13233,n12485);
  nand U13918(n13231,n13230,n12488);
  nand U13919(n13073,n13234,n12970);
  nand U13920(n13234,n13235,n13236);
  nand U13921(n13236,n12652,n13233);
  nand U13922(n13235,n12882,n13230);
  nand U13923(n13071,n13028,n13022);
  nand U13924(n13022,n13237,n13238);
  nand U13925(n13238,n12649,n13239);
  nand U13926(n13237,n12879,n12653);
  nand U13927(n13070,n13240,n12970);
  nand U13928(n13240,n13241,n13242);
  or U13929(n13242,n12820,n12822);
  or U13930(n13241,n13233,n12652);
  nand U13931(n13068,n13028,n13021);
  nand U13932(n13021,n13243,n13244);
  nand U13933(n13244,n12699,n12479);
  nand U13934(n13243,n12820,n12482);
  nand U13935(n13067,n13245,n12970);
  nand U13936(n13245,n13246,n13247);
  nand U13937(n13247,n12701,n12699);
  nand U13938(n13246,n12822,n12820);
  nand U13939(n13065,n13028,n13020);
  nand U13940(n13020,n13248,n13249);
  nand U13941(n13249,n12700,n13250);
  nand U13942(n13248,n12821,n13251);
  nand U13943(n13064,n13252,n12970);
  nand U13944(n13252,n13253,n13254);
  or U13945(n13254,n12845,n12847);
  or U13946(n13253,n12699,n12701);
  nand U13947(n13062,n13028,n13019);
  nand U13948(n13019,n13255,n13256);
  nand U13949(n13256,n12606,n12473);
  nand U13950(n13255,n12845,n12476);
  nand U13951(n13061,n13257,n12970);
  nand U13952(n13257,n13258,n13259);
  nand U13953(n13259,n12608,n12606);
  nand U13954(n13258,n12847,n12845);
  nand U13955(n13059,n13028,n13018);
  nand U13956(n13018,n13260,n13261);
  nand U13957(n13261,n12607,n13262);
  nand U13958(n13260,n12846,n13263);
  nand U13959(n13058,n13264,n12970);
  nand U13960(n13264,n13265,n13266);
  or U13961(n13266,n12771,n12773);
  or U13962(n13265,n12606,n12608);
  nand U13963(n13056,n13028,n13017);
  nand U13964(n13017,n13267,n13268);
  nand U13965(n13268,n12722,n12467);
  nand U13966(n13267,n12771,n12470);
  nand U13967(n13055,n13269,n12970);
  nand U13968(n13269,n13270,n13271);
  nand U13969(n13271,n12724,n12722);
  nand U13970(n13270,n12773,n12771);
  nand U13971(n13053,n13028,n13013);
  nand U13972(n13013,n13272,n13273);
  nand U13973(n13273,n12723,n13274);
  nand U13974(n13272,n12772,n13275);
  nand U13975(n13052,n13276,n12970);
  nand U13976(n13276,n13277,n13278);
  or U13977(n13278,n12904,n12906);
  or U13978(n13277,n12722,n12724);
  nand U13979(n13050,n13028,n13014);
  nand U13980(n13014,n13279,n13280);
  nand U13981(n13280,n12580,n12461);
  nand U13982(n13279,n12904,n12464);
  nand U13983(n13049,n13281,n12970);
  nand U13984(n13281,n13282,n13283);
  nand U13985(n13283,n12583,n12580);
  nand U13986(n13282,n12906,n12904);
  nand U13987(n13047,n13028,n13015);
  nand U13988(n13015,n13284,n13285);
  nand U13989(n13285,n12581,n13286);
  nand U13990(n13284,n12905,n13287);
  nand U13991(n13046,n13288,n12970);
  nand U13992(n13288,n13289,n13290);
  or U13993(n13290,n12662,n12664);
  or U13994(n13289,n12580,n12583);
  nand U13995(n13044,n13028,n13016);
  nand U13996(n13016,n13291,n13292);
  nand U13997(n13292,n13293,n12455);
  nand U13998(n13291,n12662,n12458);
  nand U13999(n13043,n13294,n12970);
  nand U14000(n13294,n13295,n13296);
  nand U14001(n13296,n13297,n13293);
  nand U14002(n13295,n12664,n12662);
  nand U14003(n13039,n13298,n13299,n13012);
  nand U14004(n13299,n13028,n12455);
  nand U14005(n13298,n13297,n12970);
  or U14006(n13037,n13042,n13007);
  nand U14007(n13042,n13300,n13301);
  or U14008(n13301,n12970,n12452);
  nand U14009(n13300,n13302,n12970);
  nand U14010(n13302,n13303,n13304);
  nand U14011(n13304,n13305,n13306,n13307);
  not U14012(n13305,n13308);
  nand U14013(n13035,n13034,n13011);
  nand U14014(n13034,n13309,n13310);
  nand U14015(n13310,n13028,n12449);
  nand U14016(n13309,n13311,n12970);
  xor U14017(n13311,n13312,n13313);
  xor U14018(n13312,n13303,n13314);
  nor U14019(n13314,n13315,n13316);
  nor U14020(n13315,n13317,n13318);
  nand U14021(n13303,n13308,n13319);
  nand U14022(n13319,n13307,n13306);
  nand U14023(n13307,n13320,n13321);
  nand U14024(n13308,n13322,n13323);
  nand U14025(n13323,n13324,n12452);
  nand U14026(n12959,n12948,n12970);
  nand U14027(n13326,n13327,n13328);
  nand U14028(n13325,n13329,n13330,n13331);
  nand U14029(n13331,n13332,n13333);
  nand U14030(n13330,n13334,n13335,n13336);
  or U14031(n13336,n13333,n13332);
  and U14032(n13332,n13337,n13338);
  nand U14033(n13338,n13007,n13339);
  nand U14034(n13337,n13340,n12452);
  nand U14035(n13333,n13341,n13342);
  nand U14036(n13342,n13343,n12452);
  nand U14037(n13341,n13007,n13344);
  nand U14038(n13335,n13345,n13346,n13347);
  not U14039(n13347,n13348);
  nand U14040(n13334,n13349,n13350);
  nand U14041(n13350,n13348,n13351);
  nand U14042(n13351,n13345,n13346);
  nand U14043(n13346,n13352,n13353,n13354);
  nand U14044(n13354,n13355,n13356);
  nand U14045(n13353,n13357,n13358,n13359);
  not U14046(n13359,n13360);
  nand U14047(n13352,n13361,n13362);
  nand U14048(n13362,n13360,n13363);
  nand U14049(n13363,n13357,n13358);
  nand U14050(n13358,n13364,n13365,n13366);
  nand U14051(n13366,n13367,n13368);
  nand U14052(n13365,n13369,n13370,n13371);
  not U14053(n13371,n13372);
  nand U14054(n13364,n13373,n13374);
  nand U14055(n13374,n13372,n13375);
  nand U14056(n13375,n13369,n13370);
  nand U14057(n13370,n13376,n13377,n13378);
  nand U14058(n13378,n13379,n13380);
  nand U14059(n13377,n13381,n13382,n13383);
  not U14060(n13383,n13384);
  nand U14061(n13376,n13385,n13386);
  nand U14062(n13386,n13384,n13387);
  nand U14063(n13387,n13381,n13382);
  nand U14064(n13382,n13388,n13389,n13390);
  nand U14065(n13390,n13391,n13392);
  nand U14066(n13389,n13393,n13394,n13395);
  not U14067(n13395,n13396);
  nand U14068(n13388,n13397,n13398);
  nand U14069(n13398,n13396,n13399);
  nand U14070(n13399,n13393,n13394);
  nand U14071(n13394,n13400,n13401,n13402);
  nand U14072(n13402,n13403,n13404);
  nand U14073(n13401,n13405,n13406,n13407);
  not U14074(n13407,n13408);
  nand U14075(n13400,n13409,n13410);
  nand U14076(n13410,n13408,n13411);
  nand U14077(n13411,n13405,n13406);
  nand U14078(n13406,n13412,n13413,n13414);
  nand U14079(n13414,n13415,n13416);
  nand U14080(n13413,n13417,n13418,n13419);
  not U14081(n13419,n13420);
  nand U14082(n13412,n13421,n13422);
  nand U14083(n13422,n13420,n13423);
  nand U14084(n13423,n13417,n13418);
  nand U14085(n13418,n13424,n13425,n13426);
  nand U14086(n13426,n13427,n13428);
  nand U14087(n13425,n13429,n13430,n13431);
  not U14088(n13431,n13432);
  nand U14089(n13424,n13433,n13434);
  nand U14090(n13434,n13432,n13435);
  nand U14091(n13435,n13429,n13430);
  nand U14092(n13430,n13436,n13437,n13438);
  nand U14093(n13438,n13439,n13440);
  nand U14094(n13437,n13441,n13442,n13443);
  not U14095(n13443,n13444);
  nand U14096(n13436,n13445,n13446);
  nand U14097(n13446,n13444,n13447);
  nand U14098(n13447,n13441,n13442);
  nand U14099(n13442,n13448,n13449,n13450);
  nand U14100(n13450,n13451,n13452);
  nand U14101(n13449,n13453,n13454,n13455);
  not U14102(n13455,n13456);
  nand U14103(n13448,n13457,n13458);
  nand U14104(n13458,n13456,n13459);
  nand U14105(n13459,n13453,n13454);
  nand U14106(n13454,n13460,n13461,n13462);
  nand U14107(n13462,n13463,n13464);
  nand U14108(n13461,n13465,n13466,n13467);
  not U14109(n13467,n13468);
  nand U14110(n13460,n13469,n13470);
  nand U14111(n13470,n13468,n13471);
  nand U14112(n13471,n13465,n13466);
  nand U14113(n13466,n13472,n13473,n13474);
  nand U14114(n13474,n13475,n13476);
  nand U14115(n13473,n13477,n13478,n13479);
  not U14116(n13479,n13480);
  nand U14117(n13472,n13481,n13482);
  nand U14118(n13482,n13480,n13483);
  nand U14119(n13483,n13477,n13478);
  nand U14120(n13478,n13484,n13485,n13486);
  nand U14121(n13486,n13487,n13488);
  nand U14122(n13485,n13489,n13490,n13491);
  not U14123(n13491,n13492);
  nand U14124(n13484,n13493,n13494);
  nand U14125(n13494,n13492,n13495);
  nand U14126(n13495,n13489,n13490);
  nand U14127(n13490,n13496,n13497,n13498);
  nand U14128(n13498,n13499,n13500);
  nand U14129(n13497,n13501,n13502,n13503);
  not U14130(n13503,n13504);
  nand U14131(n13496,n13505,n13506);
  nand U14132(n13506,n13504,n13507);
  nand U14133(n13507,n13501,n13502);
  nand U14134(n13502,n13508,n13509,n13510);
  nand U14135(n13510,n13511,n13512);
  nand U14136(n13509,n13513,n13514,n13515,n13516);
  nor U14137(n13516,n13517,n13518);
  and U14138(n13518,n13344,n12811);
  and U14139(n13517,n12542,n13519);
  or U14140(n13515,n13512,n13511);
  and U14141(n13511,n13520,n13514,n13521);
  nand U14142(n13521,n12689,n13344);
  nand U14143(n13520,n13522,n12539);
  nand U14144(n13512,n13523,n13524);
  nand U14145(n13524,n12689,n13339);
  nand U14146(n13523,n13340,n12539);
  nand U14147(n13513,n13525,n13526);
  nand U14148(n13526,n12811,n13339);
  nand U14149(n13525,n12542,n13340);
  nand U14150(n13508,n13527,n13528);
  or U14151(n13501,n13528,n13527);
  and U14152(n13527,n13529,n13514,n13530);
  nand U14153(n13530,n12869,n13344);
  nand U14154(n13529,n13519,n12536);
  nand U14155(n13528,n13531,n13532);
  nand U14156(n13532,n12869,n13339);
  nand U14157(n13531,n13340,n12536);
  nand U14158(n13504,n13533,n13514,n13534);
  nand U14159(n13534,n13135,n13344);
  nand U14160(n13533,n13522,n12533);
  nand U14161(n13505,n13535,n13536);
  nand U14162(n13536,n13135,n13339);
  nand U14163(n13535,n13340,n12533);
  or U14164(n13489,n13500,n13499);
  and U14165(n13499,n13537,n13514,n13538);
  nand U14166(n13538,n12787,n13344);
  nand U14167(n13537,n13519,n12530);
  nand U14168(n13500,n13539,n13540);
  nand U14169(n13540,n12787,n13339);
  nand U14170(n13539,n13340,n12530);
  nand U14171(n13492,n13541,n13514,n13542);
  nand U14172(n13542,n12749,n13344);
  nand U14173(n13541,n13522,n12527);
  nand U14174(n13493,n13543,n13544);
  nand U14175(n13544,n12749,n13339);
  nand U14176(n13543,n13340,n12527);
  or U14177(n13477,n13488,n13487);
  and U14178(n13487,n13545,n13514,n13546);
  nand U14179(n13546,n12895,n13344);
  nand U14180(n13545,n13519,n12524);
  nand U14181(n13488,n13547,n13548);
  nand U14182(n13548,n12895,n13339);
  nand U14183(n13547,n13340,n12524);
  nand U14184(n13480,n13549,n13514,n13550);
  nand U14185(n13550,n12570,n13344);
  nand U14186(n13549,n13522,n12521);
  nand U14187(n13481,n13551,n13552);
  nand U14188(n13552,n12570,n13339);
  nand U14189(n13551,n13340,n12521);
  or U14190(n13465,n13476,n13475);
  and U14191(n13475,n13553,n13514,n13554);
  nand U14192(n13554,n12677,n13344);
  nand U14193(n13553,n13519,n12518);
  nand U14194(n13476,n13555,n13556);
  nand U14195(n13556,n12677,n13339);
  nand U14196(n13555,n13340,n12518);
  nand U14197(n13468,n13557,n13514,n13558);
  nand U14198(n13558,n12800,n13344);
  nand U14199(n13557,n13522,n12515);
  nand U14200(n13469,n13559,n13560);
  nand U14201(n13560,n12800,n13339);
  nand U14202(n13559,n13340,n12515);
  or U14203(n13453,n13464,n13463);
  and U14204(n13463,n13561,n13514,n13562);
  nand U14205(n13562,n12624,n13344);
  nand U14206(n13561,n13519,n12512);
  nand U14207(n13464,n13563,n13564);
  nand U14208(n13564,n12624,n13339);
  nand U14209(n13563,n13340,n12512);
  nand U14210(n13456,n13565,n13514,n13566);
  nand U14211(n13566,n12859,n13344);
  nand U14212(n13565,n13522,n12509);
  nand U14213(n13457,n13567,n13568);
  nand U14214(n13568,n12859,n13339);
  nand U14215(n13567,n13340,n12509);
  or U14216(n13441,n13452,n13451);
  and U14217(n13451,n13569,n13514,n13570);
  nand U14218(n13570,n12713,n13344);
  nand U14219(n13569,n13519,n12506);
  nand U14220(n13452,n13571,n13572);
  nand U14221(n13572,n12713,n13339);
  nand U14222(n13571,n13340,n12506);
  nand U14223(n13444,n13573,n13514,n13574);
  nand U14224(n13574,n12836,n13344);
  nand U14225(n13573,n13522,n12503);
  nand U14226(n13445,n13575,n13576);
  nand U14227(n13576,n12836,n13339);
  nand U14228(n13575,n13340,n12503);
  or U14229(n13429,n13440,n13439);
  and U14230(n13439,n13577,n13514,n13578);
  nand U14231(n13578,n12597,n13344);
  nand U14232(n13577,n13519,n12500);
  nand U14233(n13440,n13579,n13580);
  nand U14234(n13580,n12597,n13339);
  nand U14235(n13579,n13340,n12500);
  nand U14236(n13432,n13581,n13514,n13582);
  nand U14237(n13582,n12954,n13344);
  nand U14238(n13581,n13522,n12497);
  nand U14239(n13433,n13583,n13584);
  nand U14240(n13584,n12954,n13339);
  nand U14241(n13583,n13340,n12497);
  or U14242(n13417,n13428,n13427);
  and U14243(n13427,n13585,n13514,n13586);
  nand U14244(n13586,n12737,n13344);
  nand U14245(n13585,n13519,n12494);
  nand U14246(n13428,n13587,n13588);
  nand U14247(n13588,n12737,n13339);
  nand U14248(n13587,n13340,n12494);
  nand U14249(n13420,n13589,n13514,n13590);
  nand U14250(n13590,n12762,n13344);
  nand U14251(n13589,n13522,n12491);
  nand U14252(n13421,n13591,n13592);
  nand U14253(n13592,n12762,n13339);
  nand U14254(n13591,n13340,n12491);
  or U14255(n13405,n13416,n13415);
  and U14256(n13415,n13593,n13514,n13594);
  nand U14257(n13594,n12883,n13344);
  nand U14258(n13593,n13519,n12488);
  nand U14259(n13416,n13595,n13596);
  nand U14260(n13596,n12883,n13339);
  nand U14261(n13595,n13340,n12488);
  nand U14262(n13408,n13597,n13514,n13598);
  nand U14263(n13598,n12653,n13344);
  nand U14264(n13597,n13522,n12485);
  nand U14265(n13409,n13599,n13600);
  nand U14266(n13600,n12653,n13339);
  nand U14267(n13599,n13340,n12485);
  or U14268(n13393,n13404,n13403);
  and U14269(n13403,n13601,n13514,n13602);
  nand U14270(n13602,n13239,n13344);
  nand U14271(n13601,n13519,n12482);
  nand U14272(n13404,n13603,n13604);
  nand U14273(n13604,n13239,n13339);
  nand U14274(n13603,n13340,n12482);
  nand U14275(n13396,n13605,n13514,n13606);
  nand U14276(n13606,n13251,n13344);
  nand U14277(n13605,n13522,n12479);
  nand U14278(n13397,n13607,n13608);
  nand U14279(n13608,n13251,n13339);
  nand U14280(n13607,n13340,n12479);
  or U14281(n13381,n13392,n13391);
  and U14282(n13391,n13609,n13514,n13610);
  nand U14283(n13610,n13250,n13344);
  nand U14284(n13609,n13519,n12476);
  nand U14285(n13392,n13611,n13612);
  nand U14286(n13612,n13250,n13339);
  nand U14287(n13611,n13340,n12476);
  nand U14288(n13384,n13613,n13514,n13614);
  nand U14289(n13614,n13263,n13344);
  nand U14290(n13613,n13522,n12473);
  nand U14291(n13385,n13615,n13616);
  nand U14292(n13616,n13263,n13339);
  nand U14293(n13615,n13340,n12473);
  or U14294(n13369,n13380,n13379);
  and U14295(n13379,n13617,n13514,n13618);
  nand U14296(n13618,n13262,n13344);
  nand U14297(n13617,n13519,n12470);
  nand U14298(n13380,n13619,n13620);
  nand U14299(n13620,n13262,n13339);
  nand U14300(n13619,n13340,n12470);
  nand U14301(n13372,n13621,n13514,n13622);
  nand U14302(n13622,n13275,n13344);
  nand U14303(n13621,n13522,n12467);
  nand U14304(n13373,n13623,n13624);
  nand U14305(n13624,n13275,n13339);
  nand U14306(n13623,n13340,n12467);
  or U14307(n13357,n13368,n13367);
  and U14308(n13367,n13625,n13514,n13626);
  nand U14309(n13626,n13274,n13344);
  nand U14310(n13625,n13519,n12464);
  nand U14311(n13368,n13627,n13628);
  nand U14312(n13628,n13274,n13339);
  nand U14313(n13627,n13340,n12464);
  nand U14314(n13360,n13629,n13514,n13630);
  nand U14315(n13630,n13287,n13344);
  nand U14316(n13629,n13522,n12461);
  nand U14317(n13361,n13631,n13632);
  nand U14318(n13632,n13287,n13339);
  nand U14319(n13631,n13340,n12461);
  or U14320(n13345,n13356,n13355);
  and U14321(n13355,n13633,n13514,n13634);
  nand U14322(n13634,n13286,n13344);
  nand U14323(n13633,n13519,n12458);
  nand U14324(n13519,n13514,n13635,n13636);
  nand U14325(n13356,n13637,n13638);
  nand U14326(n13638,n13286,n13339);
  nand U14327(n13637,n13340,n12458);
  nand U14328(n13348,n13639,n13514,n13640);
  nand U14329(n13640,n13012,n13344);
  and U14330(n13514,n13641,n13642,n13324);
  nand U14331(n13639,n13522,n12455);
  nand U14332(n13522,n13636,n13635);
  nand U14333(n13349,n13643,n13644);
  nand U14334(n13644,n13012,n13339);
  nand U14335(n13643,n13340,n12455);
  or U14336(n13329,n13328,n13327);
  and U14337(n13327,n13645,n13646);
  nand U14338(n13646,n13647,n13339);
  nand U14339(n13645,n13340,n12449);
  nand U14340(n13641,n12953,n12946);
  nand U14341(n13328,n13649,n13650);
  nand U14342(n13650,n13343,n12449);
  not U14343(n13343,n13636);
  nand U14344(n13636,n13339,n13651);
  nand U14345(n13651,n13317,n13652,n12952,n13653);
  not U14346(n13317,n12449);
  nand U14347(n13649,n13647,n13344);
  nand U14348(n13655,n13656,n13657);
  nand U14349(n13657,n13026,n13318);
  nand U14350(n12955,n13658,n13659,G36675);
  nand U14351(n13659,n12915,n13660,n13661);
  nand U14352(n13658,n12957,n12946);
  not U14353(n12957,n12922);
  nand U14354(G7495,n13662,n13663,n13664);
  nor U14355(n13664,n13665,n13666,n13667);
  nor U14356(n13667,n13668,n13669);
  nor U14357(n13666,n13670,n13671);
  nor U14358(n13670,n13672,n13673);
  nor U14359(n13672,n13674,n13668);
  nor U14360(n13665,n13675,n13676);
  nand U14361(n13663,n13677,n12810);
  nand U14362(n13662,G36685,G7317);
  nand U14363(G7494,n13678,n13679,n13680,n13681);
  nor U14364(n13681,n13682,n13683);
  nor U14365(n13683,G36705,n12687);
  nor U14366(n13682,n13129,n13684);
  not U14367(n13129,n12690);
  nand U14368(n13680,G36641,n13685);
  nand U14369(n13679,n13686,n13687);
  xor U14370(n13687,n13688,n13689);
  xor U14371(n13688,n13669,n13690);
  nand U14372(n13678,n13689,n13673);
  nand U14373(G7493,n13691,n13692,n13693,n13694);
  nand U14374(n13694,G36640,n13685);
  nor U14375(n13693,n13695,n13696);
  nor U14376(n13696,n13697,n13698);
  nor U14377(n13695,n13699,n13668);
  xor U14378(n13699,n13700,n13701);
  xnor U14379(n13701,n13702,n13703);
  nand U14380(n13692,n13677,n12870);
  nand U14381(n13691,G36680,G7317);
  nand U14382(G7492,n13704,n13705,n13706);
  nor U14383(n13706,n13707,n13708,n13709);
  nor U14384(n13709,n13697,n13710);
  nor U14385(n13708,n13711,n13668);
  xnor U14386(n13711,n13712,n13713);
  xor U14387(n13712,n13714,n13715);
  nor U14388(n13707,n13675,n13716);
  nand U14389(n13705,n13677,n13133);
  nand U14390(n13704,G36699,G7317);
  nand U14391(G7491,n12776,n13717,n13718);
  nor U14392(n13718,n13719,n13720,n13721);
  nor U14393(n13721,n13697,n13722);
  nor U14394(n13720,n13668,n13723);
  xor U14395(n13723,n13724,n13725);
  xnor U14396(n13724,n13726,n13727);
  nor U14397(n13719,n13675,n13728);
  nand U14398(n13717,n13677,n12786);
  nand U14399(n12776,G36687,G7317);
  nand U14400(G7490,n12740,n13729,n13730);
  nor U14401(n13730,n13731,n13732,n13733);
  nor U14402(n13733,n13697,n13734);
  nor U14403(n13732,n13735,n13668);
  xnor U14404(n13735,n13736,n13737);
  xor U14405(n13736,n13738,n13739);
  and U14406(n13731,n13685,G36637);
  nand U14407(n13729,n13677,n12748);
  nand U14408(n12740,G36690,G7317);
  nand U14409(G7489,n12886,n13740,n13741);
  nor U14410(n13741,n13742,n13743,n13744);
  nor U14411(n13744,n13697,n13745);
  nor U14412(n13743,n13668,n13746);
  xor U14413(n13746,n13747,n13748);
  xnor U14414(n13747,n13749,n13750);
  and U14415(n13742,n13685,G36636);
  nand U14416(n13740,n13677,n12894);
  nand U14417(n12886,G36678,G7317);
  nand U14418(G7488,n12553,n13751,n13752);
  nor U14419(n13752,n13753,n13754,n13755);
  nor U14420(n13755,n13697,n13756);
  nor U14421(n13754,n13757,n13668);
  xnor U14422(n13757,n13758,n13759);
  xor U14423(n13758,n13760,n13761);
  and U14424(n13753,n13685,G36635);
  nand U14425(n13751,n13677,n12568);
  nand U14426(n12553,G36704,G7317);
  nand U14427(G7487,n12667,n13762,n13763);
  nor U14428(n13763,n13764,n13765,n13766);
  nor U14429(n13766,n13697,n13767);
  nor U14430(n13765,n13668,n13768);
  xor U14431(n13768,n13769,n13770);
  xnor U14432(n13769,n13771,n13772);
  nor U14433(n13764,n13675,n13773);
  nand U14434(n13762,n13677,n12676);
  nand U14435(n12667,G36696,G7317);
  nand U14436(G7486,n12790,n13774,n13775);
  nor U14437(n13775,n13776,n13777,n13778);
  nor U14438(n13778,n13697,n13779);
  nor U14439(n13777,n13780,n13668);
  xnor U14440(n13780,n13781,n13782);
  xor U14441(n13781,n13783,n13784);
  nor U14442(n13776,n13675,n13785);
  nand U14443(n13774,n13677,n12799);
  nand U14444(n12790,G36686,G7317);
  nand U14445(G7485,n13786,n13787,n13788,n13789);
  nor U14446(n13789,n13790,n13791);
  nor U14447(n13791,G36705,n13792);
  nor U14448(n13790,n13181,n13684);
  nand U14449(n13788,G36632,n13685);
  nand U14450(n13787,n13686,n13793);
  xor U14451(n13793,n13794,n13795);
  nand U14452(n13795,n13796,n13797);
  not U14453(n13686,n13668);
  nand U14454(n13786,n13798,n13673);
  nand U14455(G7484,n12850,n13799,n13800);
  nor U14456(n13800,n13801,n13802,n13803);
  nor U14457(n13803,n13697,n13804);
  nor U14458(n13802,n13805,n13668);
  xnor U14459(n13805,n13806,n13807);
  xor U14460(n13806,n13808,n13809);
  and U14461(n13801,n13685,G36631);
  nand U14462(n13799,n13677,n12858);
  nand U14463(n12850,G36681,G7317);
  nand U14464(G7483,n12704,n13810,n13811);
  nor U14465(n13811,n13812,n13813,n13814);
  nor U14466(n13814,n13697,n13815);
  nor U14467(n13813,n13668,n13816);
  xor U14468(n13816,n13817,n13818);
  xnor U14469(n13817,n13819,n13820);
  and U14470(n13812,n13685,G36630);
  nand U14471(n13810,n13677,n12712);
  nand U14472(n12704,G36693,G7317);
  nand U14473(G7482,n12825,n13821,n13822);
  nor U14474(n13822,n13823,n13824,n13825);
  nor U14475(n13825,n13697,n13826);
  nor U14476(n13824,n13827,n13668);
  xnor U14477(n13827,n13828,n13829);
  xor U14478(n13828,n13830,n13831);
  nor U14479(n13823,n13675,n13832);
  nand U14480(n13821,n13677,n12835);
  nand U14481(n12825,G36683,G7317);
  nand U14482(G7481,n12586,n13833,n13834);
  nor U14483(n13834,n13835,n13836,n13837);
  nor U14484(n13837,n13697,n13838);
  nor U14485(n13836,n13668,n13839);
  xor U14486(n13839,n13840,n13841);
  xnor U14487(n13840,n13842,n13843);
  nor U14488(n13835,n13675,n13844);
  nand U14489(n13833,n13677,n12596);
  nand U14490(n12586,G36702,G7317);
  nand U14491(G7480,n12909,n13845,n13846);
  nor U14492(n13846,n13847,n13848,n13849);
  nor U14493(n13849,n13697,n13850);
  nor U14494(n13848,n13851,n13668);
  xnor U14495(n13851,n13852,n13853);
  xor U14496(n13852,n13854,n13855);
  and U14497(n13847,n13685,G36627);
  nand U14498(n13845,n13677,n12938);
  nand U14499(n12909,G36676,G7317);
  nand U14500(G7479,n12727,n13856,n13857);
  nor U14501(n13857,n13858,n13859,n13860);
  nor U14502(n13860,n13697,n13861);
  nor U14503(n13859,n13668,n13862);
  xor U14504(n13862,n13863,n13864);
  xnor U14505(n13863,n13865,n13866);
  nor U14506(n13858,n13675,n13867);
  nand U14507(n13856,n13677,n12736);
  nand U14508(n12727,G36691,G7317);
  nand U14509(G7478,n12752,n13868,n13869);
  nor U14510(n13869,n13870,n13871,n13872);
  nor U14511(n13872,n13697,n13873);
  nor U14512(n13871,n13874,n13668);
  xnor U14513(n13874,n13875,n13876);
  xor U14514(n13875,n13877,n13878);
  nor U14515(n13870,n13675,n13879);
  nand U14516(n13868,n13677,n12761);
  nand U14517(n12752,G36689,G7317);
  nand U14518(G7477,n12873,n13880,n13881);
  nor U14519(n13881,n13882,n13883,n13884);
  nor U14520(n13884,n13697,n13885);
  nor U14521(n13883,n13668,n13886,n13887);
  nor U14522(n13887,n13885,n13888,n13889);
  nor U14523(n13886,n13890,n13891);
  xor U14524(n13890,n13892,n13893);
  and U14525(n13882,n13685,G36624);
  not U14526(n13685,n13675);
  nand U14527(n13880,n13677,n12882);
  nand U14528(n12873,G36679,G7317);
  nand U14529(G7476,n12642,n13894,n13895);
  nor U14530(n13895,n13896,n13897,n13898);
  nor U14531(n13898,n13697,n13899);
  not U14532(n13697,n13673);
  nand U14533(n13673,n13900,n13901);
  nand U14534(n13901,n13902,n13675,n13903);
  nand U14535(n13902,n12922,n13904);
  nand U14536(n13904,n12923,n13905);
  nand U14537(n13900,n13661,G7605);
  nor U14538(n13897,n13668,n13906,n13907);
  nor U14539(n13907,n13908,n13889,n13909);
  nor U14540(n13909,n13888,n13891);
  nor U14541(n13906,n13910,n13888,n13911);
  nor U14542(n13911,n13889,n13885);
  and U14543(n13889,n13892,n13893);
  nor U14544(n13888,n13892,n13893);
  nand U14545(n13893,n13912,n13913);
  nand U14546(n13913,n13914,G36577);
  nand U14547(n13912,n13915,G36609);
  nand U14548(n13892,n13916,n13917);
  nand U14549(n13917,n13918,n13873);
  or U14550(n13918,n13876,n13877);
  nand U14551(n13916,n13876,n13877);
  nand U14552(n13877,n13919,n13920);
  nand U14553(n13920,n13861,n13921);
  or U14554(n13921,n13866,n13865);
  nand U14555(n13919,n13866,n13865);
  nand U14556(n13865,n13922,n13923);
  nand U14557(n13923,n13924,n13850);
  or U14558(n13924,n13853,n13854);
  nand U14559(n13922,n13853,n13854);
  nand U14560(n13854,n13925,n13926);
  nand U14561(n13926,n13838,n13927);
  or U14562(n13927,n13843,n13842);
  nand U14563(n13925,n13843,n13842);
  nand U14564(n13842,n13928,n13929);
  nand U14565(n13929,n13930,n13826);
  or U14566(n13930,n13829,n13830);
  nand U14567(n13928,n13829,n13830);
  nand U14568(n13830,n13931,n13932);
  nand U14569(n13932,n13815,n13933);
  or U14570(n13933,n13820,n13819);
  nand U14571(n13931,n13820,n13819);
  nand U14572(n13819,n13934,n13935);
  nand U14573(n13935,n13936,n13804);
  or U14574(n13936,n13807,n13808);
  nand U14575(n13934,n13807,n13808);
  nand U14576(n13808,n13937,n13796);
  nand U14577(n13796,n13938,n13939);
  nand U14578(n13937,n13794,n13797);
  nand U14579(n13797,n13940,n13798);
  not U14580(n13940,n13939);
  nand U14581(n13939,n13941,n13942);
  nand U14582(n13942,n13914,G36569);
  nand U14583(n13941,n13915,G36601);
  nand U14584(n13794,n13943,n13944);
  nand U14585(n13944,n13945,n13779);
  or U14586(n13945,n13782,n13783);
  nand U14587(n13943,n13782,n13783);
  nand U14588(n13783,n13946,n13947);
  nand U14589(n13947,n13767,n13948);
  or U14590(n13948,n13772,n13771);
  nand U14591(n13946,n13772,n13771);
  nand U14592(n13771,n13949,n13950);
  nand U14593(n13950,n13951,n13756);
  or U14594(n13951,n13759,n13760);
  nand U14595(n13949,n13759,n13760);
  nand U14596(n13760,n13952,n13953);
  nand U14597(n13953,n13745,n13954);
  or U14598(n13954,n13750,n13749);
  nand U14599(n13952,n13750,n13749);
  nand U14600(n13749,n13955,n13956);
  nand U14601(n13956,n13957,n13734);
  or U14602(n13957,n13737,n13738);
  nand U14603(n13955,n13737,n13738);
  nand U14604(n13738,n13958,n13959);
  nand U14605(n13959,n13722,n13960);
  or U14606(n13960,n13727,n13726);
  nand U14607(n13958,n13727,n13726);
  nand U14608(n13726,n13961,n13962);
  nand U14609(n13962,n13963,n13710);
  or U14610(n13963,n13713,n13714);
  nand U14611(n13961,n13713,n13714);
  nand U14612(n13714,n13964,n13965);
  nand U14613(n13965,n13698,n13966);
  or U14614(n13966,n13703,n13702);
  nand U14615(n13964,n13702,n13703);
  nand U14616(n13703,n13967,n13968);
  nand U14617(n13968,n13914,G36561);
  nand U14618(n13967,n13915,G36593);
  and U14619(n13702,n13969,n13970);
  nand U14620(n13970,n13689,n13971);
  or U14621(n13971,n13669,n13690);
  nand U14622(n13969,n13690,n13669);
  nand U14623(n13669,n13671,n13674);
  nand U14624(n13674,n13972,n13973);
  nand U14625(n13973,n13914,G36559);
  nand U14626(n13972,n13915,G36591);
  and U14627(n13690,n13974,n13975);
  nand U14628(n13975,n13914,G36560);
  nand U14629(n13974,n13915,G36592);
  nand U14630(n13713,n13976,n13977);
  nand U14631(n13977,n13914,G36562);
  nand U14632(n13976,n13915,G36594);
  nand U14633(n13727,n13978,n13979);
  nand U14634(n13979,n13914,G36563);
  nand U14635(n13978,n13915,G36595);
  nand U14636(n13737,n13980,n13981);
  nand U14637(n13981,n13914,G36564);
  nand U14638(n13980,n13915,G36596);
  nand U14639(n13750,n13982,n13983);
  nand U14640(n13983,n13914,G36565);
  nand U14641(n13982,n13915,G36597);
  nand U14642(n13759,n13984,n13985);
  nand U14643(n13985,n13914,G36566);
  nand U14644(n13984,n13915,G36598);
  nand U14645(n13772,n13986,n13987);
  nand U14646(n13987,n13914,G36567);
  nand U14647(n13986,n13915,G36599);
  nand U14648(n13782,n13988,n13989);
  nand U14649(n13989,n13914,G36568);
  nand U14650(n13988,n13915,G36600);
  nand U14651(n13807,n13990,n13991);
  nand U14652(n13991,n13914,G36570);
  nand U14653(n13990,n13915,G36602);
  nand U14654(n13820,n13992,n13993);
  nand U14655(n13993,n13914,G36571);
  nand U14656(n13992,n13915,G36603);
  nand U14657(n13829,n13994,n13995);
  nand U14658(n13995,n13914,G36572);
  nand U14659(n13994,n13915,G36604);
  nand U14660(n13843,n13996,n13997);
  nand U14661(n13997,n13914,G36573);
  nand U14662(n13996,n13915,G36605);
  nand U14663(n13853,n13998,n13999);
  nand U14664(n13999,n13914,G36574);
  nand U14665(n13998,n13915,G36606);
  nand U14666(n13866,n14000,n14001);
  nand U14667(n14001,n13914,G36575);
  nand U14668(n14000,n13915,G36607);
  nand U14669(n13876,n14002,n14003);
  nand U14670(n14003,n13914,G36576);
  nand U14671(n14002,n13915,G36608);
  not U14672(n13910,n13908);
  xor U14673(n13908,n14004,n12971);
  nand U14674(n14004,n14005,n14006);
  nand U14675(n14006,n13914,G36578);
  and U14676(n13914,n13660,n14007);
  nand U14677(n14005,n13915,G36610);
  and U14678(n13915,n14007,n14008);
  or U14679(n14007,n13905,n13324);
  nand U14680(n13668,n13661,n14009);
  nand U14681(n14009,n12922,n14010);
  nand U14682(n14010,n13905,n13675,n12923);
  nand U14683(n13905,n14011,n14012,n14013,n14014);
  not U14684(n14014,n12933);
  nor U14685(n14013,n14015,n13026);
  nand U14686(n12922,n13324,G36705);
  nor U14687(n13896,n14016,n13675);
  nand U14688(n13675,n14017,n14018);
  nand U14689(n13894,n13677,n12652);
  not U14690(n13677,n13684);
  nand U14691(n13684,G7605,n13903);
  nand U14692(n12642,G36698,G7317);
  nand U14693(G7475,n14019,n14020,n14021);
  nand U14694(n14020,n14022,n13647);
  nand U14695(n14019,n14023,G36622);
  nand U14696(G7474,n14024,n14025,n14021);
  and U14697(n14021,n14026,n14027);
  nand U14698(n14027,n14028,n14029);
  nand U14699(n14025,n14022,n13007);
  nand U14700(n14024,n14023,G36621);
  nand U14701(G7473,n14030,n14031,n14032,n14033);
  nor U14702(n14033,n14034,n14035,n14036);
  nor U14703(n14036,n12581,n14037);
  not U14704(n14035,n14026);
  nand U14705(n14026,n14038,n14039,n14040);
  nor U14706(n14034,n13293,n14041);
  nand U14707(n14032,n14042,n13297);
  or U14708(n14031,n14043,n14023);
  nand U14709(n14030,n14023,G36620);
  nand U14710(G7472,n14044,n14045,n14046,n14047);
  nor U14711(n14047,n14048,n14049,n14050);
  nor U14712(n14050,n12662,n14041);
  nor U14713(n14049,n12905,n14037);
  nor U14714(n14048,n12661,n14051);
  not U14715(n12661,n14052);
  nand U14716(n14046,n14023,G36619);
  nand U14717(n14045,n14042,n12664);
  nand U14718(n14044,n14053,n12455);
  nand U14719(G7471,n14054,n14055,n14056,n14057);
  nor U14720(n14057,n14058,n14059,n14060);
  nor U14721(n14060,n12580,n14041);
  nor U14722(n14059,n12723,n14037);
  nor U14723(n14058,n12578,n14051);
  nand U14724(n14056,n14023,G36618);
  nand U14725(n14055,n14042,n12583);
  nand U14726(n14054,n14053,n12458);
  nand U14727(G7470,n14061,n14062,n14063,n14064);
  nor U14728(n14064,n14065,n14066,n14067);
  nor U14729(n14067,n12904,n14041);
  nor U14730(n14066,n12772,n14037);
  nor U14731(n14065,n12903,n14051);
  not U14732(n12903,n14068);
  nand U14733(n14063,n14023,G36617);
  nand U14734(n14062,n14042,n12906);
  nand U14735(n14061,n14053,n12461);
  nand U14736(G7469,n14069,n14070,n14071,n14072);
  nor U14737(n14072,n14073,n14074,n14075);
  nor U14738(n14075,n12722,n14041);
  nor U14739(n14074,n12607,n14037);
  nor U14740(n14073,n12721,n14051);
  not U14741(n12721,n14076);
  nand U14742(n14071,n14023,G36616);
  nand U14743(n14070,n14042,n12724);
  nand U14744(n14069,n14053,n12464);
  nand U14745(G7468,n14077,n14078,n14079,n14080);
  nor U14746(n14080,n14081,n14082,n14083);
  nor U14747(n14083,n12771,n14041);
  nor U14748(n14082,n12846,n14037);
  nor U14749(n14081,n12770,n14051);
  not U14750(n12770,n14084);
  nand U14751(n14079,n14023,G36615);
  nand U14752(n14078,n14042,n12773);
  nand U14753(n14077,n14053,n12467);
  nand U14754(G7467,n14085,n14086,n14087,n14088);
  nor U14755(n14088,n14089,n14090,n14091);
  nor U14756(n14091,n12606,n14041);
  nor U14757(n14090,n12700,n14037);
  nor U14758(n14089,n12605,n14051);
  not U14759(n12605,n14092);
  nand U14760(n14087,n14023,G36614);
  nand U14761(n14086,n14042,n12608);
  nand U14762(n14085,n14053,n12470);
  nand U14763(G7466,n14093,n14094,n14095,n14096);
  nor U14764(n14096,n14097,n14098,n14099);
  nor U14765(n14099,n12845,n14041);
  nor U14766(n14098,n12821,n14037);
  nor U14767(n14097,n12844,n14051);
  not U14768(n12844,n14100);
  nand U14769(n14095,n14023,G36613);
  nand U14770(n14094,n14042,n12847);
  nand U14771(n14093,n14053,n12473);
  nand U14772(G7465,n14101,n14102,n14103,n14104);
  nor U14773(n14104,n14105,n14106,n14107);
  nor U14774(n14107,n12699,n14041);
  nor U14775(n14106,n12649,n14037);
  nor U14776(n14105,n12698,n14051);
  not U14777(n12698,n14108);
  nand U14778(n14103,n14023,G36612);
  nand U14779(n14102,n14042,n12701);
  nand U14780(n14101,n14053,n12476);
  nand U14781(G7464,n14109,n14110,n14111,n14112);
  nor U14782(n14112,n14113,n14114,n14115);
  nor U14783(n14115,n12820,n14041);
  nor U14784(n14114,n12879,n14037);
  nor U14785(n14113,n12819,n14051);
  not U14786(n12819,n14116);
  nand U14787(n14111,n14023,G36611);
  nand U14788(n14110,n14042,n12822);
  nand U14789(n14109,n14053,n12479);
  nand U14790(G7463,n14117,n14118,n14119,n14120);
  nor U14791(n14120,n14121,n14122,n14123);
  nor U14792(n14123,n12651,n14041);
  not U14793(n12651,n14124);
  nor U14794(n14122,n12648,n14037);
  nor U14795(n14121,n12650,n14051);
  not U14796(n12650,n14125);
  nand U14797(n14119,n14023,G36610);
  nand U14798(n14118,n14042,n12652);
  nand U14799(n14117,n14053,n12482);
  nand U14800(G7462,n14126,n14127,n14128,n14129);
  nor U14801(n14129,n14130,n14131,n14132);
  nor U14802(n14132,n12881,n14041);
  not U14803(n12881,n14133);
  nor U14804(n14131,n12733,n14037);
  nor U14805(n14130,n12880,n14051);
  nand U14806(n14128,n14023,G36609);
  nand U14807(n14127,n14042,n12882);
  nand U14808(n14126,n14053,n12485);
  nand U14809(G7461,n14134,n14135,n14136,n14137);
  nor U14810(n14137,n14138,n14139,n14140);
  nor U14811(n14140,n12760,n14041);
  not U14812(n12760,n14141);
  nor U14813(n14139,n12758,n14037);
  nor U14814(n14138,n12759,n14051);
  not U14815(n12759,n14142);
  nand U14816(n14136,n14023,G36608);
  nand U14817(n14135,n14042,n12761);
  nand U14818(n14134,n14053,n12488);
  nand U14819(G7460,n14143,n14144,n14145,n14146);
  nor U14820(n14146,n14147,n14148,n14149);
  nor U14821(n14149,n12735,n14041);
  not U14822(n12735,n14150);
  nor U14823(n14148,n12593,n14037);
  nor U14824(n14147,n12734,n14051);
  not U14825(n12734,n14151);
  nand U14826(n14145,n14023,G36607);
  nand U14827(n14144,n14042,n12736);
  nand U14828(n14143,n14053,n12491);
  nand U14829(G7459,n14152,n14153,n14154,n14155);
  nor U14830(n14155,n14156,n14157,n14158);
  nor U14831(n14158,n12936,n14041);
  not U14832(n12936,n14159);
  nor U14833(n14157,n12832,n14037);
  nor U14834(n14156,n12919,n14051);
  not U14835(n12919,n14160);
  nand U14836(n14154,n14023,G36606);
  nand U14837(n14153,n14042,n12938);
  nand U14838(n14152,n14053,n12494);
  nand U14839(G7458,n14161,n14162,n14163,n14164);
  nor U14840(n14164,n14165,n14166,n14167);
  nor U14841(n14167,n12595,n14041);
  not U14842(n12595,n14168);
  nor U14843(n14166,n12592,n14037);
  nor U14844(n14165,n12594,n14051);
  nand U14845(n14163,n14023,G36605);
  nand U14846(n14162,n14042,n12596);
  nand U14847(n14161,n14053,n12497);
  nand U14848(G7457,n14169,n14170,n14171,n14172);
  nor U14849(n14172,n14173,n14174,n14175);
  nor U14850(n14175,n12834,n14041);
  not U14851(n12834,n14176);
  nor U14852(n14174,n12831,n14037);
  nor U14853(n14173,n12833,n14051);
  not U14854(n12833,n14177);
  nand U14855(n14171,n14023,G36604);
  nand U14856(n14170,n14042,n12835);
  nand U14857(n14169,n14053,n12500);
  nand U14858(G7456,n14178,n14179,n14180,n14181);
  nor U14859(n14181,n14182,n14183,n14184);
  nor U14860(n14184,n12711,n14041);
  not U14861(n12711,n14185);
  nor U14862(n14183,n12618,n14037);
  nor U14863(n14182,n12710,n14051);
  nand U14864(n14180,n14023,G36603);
  nand U14865(n14179,n14042,n12712);
  nand U14866(n14178,n14053,n12503);
  nand U14867(G7455,n14186,n14187,n14188,n14189);
  nor U14868(n14189,n14190,n14191,n14192);
  nor U14869(n14192,n12857,n14041);
  not U14870(n12857,n14193);
  nor U14871(n14191,n12796,n14037);
  nor U14872(n14190,n12856,n14051);
  not U14873(n12856,n14194);
  nand U14874(n14188,n14023,G36602);
  nand U14875(n14187,n14042,n12858);
  nand U14876(n14186,n14053,n12506);
  nand U14877(G7454,n14195,n14196,n14197,n14198);
  nor U14878(n14198,n14199,n14200,n14201);
  nor U14879(n14201,n12618,n14202);
  nor U14880(n14200,n13181,n14203);
  and U14881(n14199,G36601,n14023);
  nand U14882(n14197,n14040,n12620);
  not U14883(n14040,n14051);
  or U14884(n14196,n14037,n12617);
  nand U14885(n14195,n14022,n12621);
  nand U14886(G7453,n14204,n14205,n14206,n14207);
  nor U14887(n14207,n14208,n14209,n14210);
  nor U14888(n14210,n12798,n14041);
  not U14889(n12798,n14211);
  nor U14890(n14209,n12561,n14037);
  nor U14891(n14208,n12797,n14051);
  nand U14892(n14206,n14023,G36600);
  nand U14893(n14205,n14042,n12799);
  nand U14894(n14204,n14053,n12512);
  nand U14895(G7452,n14212,n14213,n14214,n14215);
  nor U14896(n14215,n14216,n14217,n14218);
  nor U14897(n14218,n12675,n14041);
  not U14898(n12675,n14219);
  nor U14899(n14217,n12673,n14037);
  nor U14900(n14216,n12674,n14051);
  nand U14901(n14214,n14023,G36599);
  nand U14902(n14213,n14042,n12676);
  nand U14903(n14212,n14053,n12515);
  nand U14904(G7451,n14220,n14221,n14222,n14223);
  nor U14905(n14223,n14224,n14225,n14226);
  nor U14906(n14226,n12565,n14041);
  not U14907(n12565,n14227);
  nor U14908(n14225,n12559,n14037);
  nor U14909(n14224,n12563,n14051);
  not U14910(n12563,n14228);
  nand U14911(n14222,n14023,G36598);
  nand U14912(n14221,n14042,n12568);
  nand U14913(n14220,n14053,n12518);
  nand U14914(G7450,n14229,n14230,n14231,n14232);
  nor U14915(n14232,n14233,n14234,n14235);
  nor U14916(n14235,n12893,n14041);
  not U14917(n12893,n14236);
  nor U14918(n14234,n12783,n14037);
  nor U14919(n14233,n12892,n14051);
  not U14920(n12892,n14237);
  nand U14921(n14231,n14023,G36597);
  nand U14922(n14229,n14053,n12521);
  nand U14923(G7449,n14238,n14239,n14240,n14241);
  nor U14924(n14241,n14242,n14243,n14244);
  nor U14925(n14244,n12747,n14041);
  not U14926(n12747,n14245);
  nor U14927(n14243,n12639,n14037);
  nor U14928(n14242,n12746,n14051);
  not U14929(n12746,n14246);
  nand U14930(n14240,n14023,G36596);
  nand U14931(n14239,n14042,n12748);
  nand U14932(G7448,n14247,n14248,n14249,n14250);
  nor U14933(n14250,n14251,n14252,n14253);
  nor U14934(n14253,n12785,n14041);
  not U14935(n12785,n14254);
  nor U14936(n14252,n12782,n14037);
  nor U14937(n14251,n12784,n14051);
  nand U14938(n14249,n14023,G36595);
  nand U14939(n14248,n14042,n12786);
  nand U14940(n14247,n14053,n12527);
  nand U14941(G7447,n14255,n14256,n14257,n14258);
  nor U14942(n14258,n14259,n14260,n14261);
  and U14943(n14261,n12638,n14022);
  not U14944(n14022,n14041);
  nor U14945(n14260,n12688,n14037);
  nor U14946(n14259,G36699,n14051);
  nand U14947(n14257,n14023,G36594);
  nand U14948(n14256,n14042,n13133);
  nand U14949(n14255,n14053,n12530);
  nand U14950(G7446,n14262,n14263,n14264,n14265);
  nor U14951(n14265,n14266,n14267,n14268);
  nor U14952(n14268,n12867,n14041);
  not U14953(n12867,n14269);
  nor U14954(n14267,n12809,n14037);
  nor U14955(n14266,n12868,n14051);
  not U14956(n12868,G36680);
  nand U14957(n14264,n14023,G36593);
  nand U14958(n14263,n14042,n12870);
  nand U14959(n14262,n14053,n12533);
  nand U14960(G7445,n14270,n14271,n14272,n14273);
  nor U14961(n14273,n14274,n14275,n14276);
  nor U14962(n14276,n12685,n14041);
  not U14963(n12685,n14277);
  nor U14964(n14275,n13139,n14037);
  nand U14965(n14037,n14278,n14029);
  not U14966(n13139,n12542);
  nor U14967(n14274,n12687,n14051);
  not U14968(n12687,G36695);
  nand U14969(n14272,n14053,n12536);
  nand U14970(n14271,n12690,n14279,n14029);
  nand U14971(n14279,n13642,n13654,n14280,n14281);
  nor U14972(n14281,n14282,n14283);
  nand U14973(n14280,n14284,n13026);
  nand U14974(n14270,n14023,G36592);
  nand U14975(G7444,n14285,n14286,n14287,n14288);
  nand U14976(n14288,n14042,n12810);
  not U14977(n14042,n14203);
  nand U14978(n14203,n14029,n14289);
  nand U14979(n14289,n12942,n14290);
  nand U14980(n14290,n13653,n12935);
  nor U14981(n14287,n14291,n14292);
  nor U14982(n14292,n12808,n14051);
  nand U14983(n14051,n14015,n14029);
  not U14984(n12808,G36685);
  nor U14985(n14291,n12807,n14041);
  nand U14986(n14041,n14029,n12933);
  nand U14987(n12933,n14293,n14294);
  nand U14988(n14294,n12951,n13025);
  nor U14989(n12951,n12974,n13026,n13899);
  nand U14990(n14293,n14295,n13899);
  not U14991(n12807,n14296);
  nand U14992(n14286,n14053,n12539);
  not U14993(n14053,n14202);
  nand U14994(n14202,n14297,n14029);
  nand U14995(n14285,n14023,G36591);
  nand U14996(n14029,n12634,n14298);
  nand U14997(n14298,n14299,n14300,n14301);
  nand U14998(n14300,n14302,n14303);
  nand U14999(n14299,n14304,n14305);
  nand U15000(n14305,n13635,n13029);
  nand U15001(n12634,n14015,n12923);
  not U15002(n14015,n14306);
  nand U15003(G7443,n14307,n14308,n14309);
  nand U15004(n14309,n14310,n13647);
  nand U15005(n14308,G36590,n14311);
  nand U15006(G7442,n14307,n14312,n14313);
  nand U15007(n14313,n14310,n13007);
  nand U15008(n14312,G36589,n14311);
  nand U15009(n14307,n14314,n14028);
  nand U15010(G7441,n14315,n14316,n14317,n14318);
  nand U15011(n14318,n14319,n12458);
  nand U15012(n14317,n14310,n13012);
  nand U15013(n14316,n14320,n13297);
  nor U15014(n14315,n14321,n14322);
  nor U15015(n14322,n14311,n14043);
  and U15016(n14321,n14311,G36588);
  nand U15017(G7440,n14323,n14324,n14325,n14326);
  nor U15018(n14326,n14327,n14328);
  and U15019(n14328,n14311,G36587);
  nor U15020(n14327,n12663,n14329);
  nand U15021(n14325,n14320,n12664);
  nand U15022(n14324,n14319,n12461);
  nand U15023(n14323,n14310,n13286);
  nand U15024(G7439,n14330,n14331,n14332,n14333);
  nor U15025(n14333,n14334,n14335);
  and U15026(n14335,n14311,G36586);
  nor U15027(n14334,n12581,n14329);
  nand U15028(n14332,n14320,n12583);
  nand U15029(n14331,n14319,n12464);
  nand U15030(n14330,n14310,n13287);
  nand U15031(G7438,n14336,n14337,n14338,n14339);
  nor U15032(n14339,n14340,n14341);
  and U15033(n14341,n14311,G36585);
  nor U15034(n14340,n12905,n14329);
  nand U15035(n14338,n14320,n12906);
  nand U15036(n14337,n14319,n12467);
  nand U15037(n14336,n14310,n13274);
  nand U15038(G7437,n14342,n14343,n14344,n14345);
  nor U15039(n14345,n14346,n14347);
  and U15040(n14347,n14311,G36584);
  nor U15041(n14346,n12723,n14329);
  nand U15042(n14344,n14320,n12724);
  nand U15043(n14343,n14319,n12470);
  nand U15044(n14342,n14310,n13275);
  nand U15045(G7436,n14348,n14349,n14350,n14351);
  nor U15046(n14351,n14352,n14353);
  and U15047(n14353,n14311,G36583);
  nor U15048(n14352,n12772,n14329);
  nand U15049(n14350,n14320,n12773);
  nand U15050(n14349,n14319,n12473);
  nand U15051(n14348,n14310,n13262);
  nand U15052(G7435,n14354,n14355,n14356,n14357);
  nor U15053(n14357,n14358,n14359);
  and U15054(n14359,n14311,G36582);
  nor U15055(n14358,n12607,n14329);
  nand U15056(n14356,n14320,n12608);
  nand U15057(n14355,n14319,n12476);
  nand U15058(n14354,n14310,n13263);
  nand U15059(G7434,n14360,n14361,n14362,n14363);
  nor U15060(n14363,n14364,n14365);
  and U15061(n14365,n14311,G36581);
  nor U15062(n14364,n12846,n14329);
  nand U15063(n14362,n14320,n12847);
  nand U15064(n14361,n14319,n12479);
  nand U15065(n14360,n14310,n13250);
  nand U15066(G7433,n14366,n14367,n14368,n14369);
  nor U15067(n14369,n14370,n14371);
  and U15068(n14371,n14311,G36580);
  nor U15069(n14370,n12700,n14329);
  nand U15070(n14368,n14320,n12701);
  nand U15071(n14367,n14319,n12482);
  nand U15072(n14366,n14310,n13251);
  nand U15073(G7432,n14372,n14373,n14374,n14375);
  nor U15074(n14375,n14376,n14377);
  and U15075(n14377,n14311,G36579);
  nor U15076(n14376,n12821,n14329);
  nand U15077(n14374,n14320,n12822);
  nand U15078(n14373,n14319,n12485);
  nand U15079(n14372,n14310,n13239);
  nand U15080(G7431,n14378,n14379,n14380,n14381);
  nor U15081(n14381,n14382,n14383);
  and U15082(n14383,n14311,G36578);
  nor U15083(n14382,n12649,n14329);
  nand U15084(n14380,n14320,n12652);
  nand U15085(n14379,n14319,n12488);
  nand U15086(n14378,n14310,n14124);
  nand U15087(G7430,n14384,n14385,n14386,n14387);
  nor U15088(n14387,n14388,n14389);
  and U15089(n14389,n14311,G36577);
  nor U15090(n14388,n12879,n14329);
  nand U15091(n14386,n14320,n12882);
  nand U15092(n14385,n14319,n12491);
  nand U15093(n14384,n14310,n14133);
  nand U15094(G7429,n14390,n14391,n14392,n14393);
  nor U15095(n14393,n14394,n14395);
  and U15096(n14395,n14311,G36576);
  nor U15097(n14394,n12648,n14329);
  nand U15098(n14392,n14320,n12761);
  nand U15099(n14391,n14319,n12494);
  nand U15100(n14390,n14310,n14141);
  nand U15101(G7428,n14396,n14397,n14398,n14399);
  nor U15102(n14399,n14400,n14401);
  and U15103(n14401,n14311,G36575);
  nor U15104(n14400,n12733,n14329);
  nand U15105(n14398,n14320,n12736);
  nand U15106(n14397,n14319,n12497);
  nand U15107(n14396,n14310,n14150);
  nand U15108(G7427,n14402,n14403,n14404,n14405);
  nor U15109(n14405,n14406,n14407);
  and U15110(n14407,n14311,G36574);
  nor U15111(n14406,n12758,n14329);
  nand U15112(n14404,n14320,n12938);
  nand U15113(n14403,n14319,n12500);
  nand U15114(n14402,n14310,n14159);
  nand U15115(G7426,n14408,n14409,n14410,n14411);
  nor U15116(n14411,n14412,n14413);
  and U15117(n14413,n14311,G36573);
  nor U15118(n14412,n12593,n14329);
  nand U15119(n14410,n14320,n12596);
  nand U15120(n14409,n14319,n12503);
  nand U15121(n14408,n14310,n14168);
  nand U15122(G7425,n14414,n14415,n14416,n14417);
  nor U15123(n14417,n14418,n14419);
  and U15124(n14419,n14311,G36572);
  nor U15125(n14418,n12832,n14329);
  nand U15126(n14416,n14320,n12835);
  nand U15127(n14415,n14319,n12506);
  nand U15128(n14414,n14310,n14176);
  nand U15129(G7424,n14420,n14421,n14422,n14423);
  nor U15130(n14423,n14424,n14425);
  and U15131(n14425,n14311,G36571);
  nor U15132(n14424,n12592,n14329);
  nand U15133(n14422,n14320,n12712);
  nand U15134(n14421,n14319,n12509);
  nand U15135(n14420,n14310,n14185);
  nand U15136(G7423,n14426,n14427,n14428,n14429);
  nor U15137(n14429,n14430,n14431);
  and U15138(n14431,n14311,G36570);
  nor U15139(n14430,n12831,n14329);
  nand U15140(n14428,n14320,n12858);
  nand U15141(n14427,n14319,n12512);
  nand U15142(n14426,n14310,n14193);
  nand U15143(G7422,n14432,n14433,n14434);
  nor U15144(n14434,n14435,n14436,n14437);
  and U15145(n14437,n12621,n14310);
  nor U15146(n14436,n12617,n14438);
  nor U15147(n14435,n13181,n14439);
  nand U15148(n14433,n14440,n12509);
  nand U15149(n14432,G36569,n14311);
  nand U15150(G7421,n14441,n14442,n14443,n14444);
  nor U15151(n14444,n14445,n14446);
  and U15152(n14446,n14311,G36568);
  nor U15153(n14445,n12796,n14329);
  nand U15154(n14443,n14320,n12799);
  nand U15155(n14442,n14319,n12518);
  nand U15156(n14441,n14310,n14211);
  nand U15157(G7420,n14447,n14448,n14449,n14450);
  nor U15158(n14450,n14451,n14452);
  and U15159(n14452,n14311,G36567);
  nor U15160(n14451,n12617,n14329);
  not U15161(n12617,n12515);
  nand U15162(n14449,n14320,n12676);
  nand U15163(n14448,n14319,n12521);
  nand U15164(n14447,n14310,n14219);
  nand U15165(G7419,n14453,n14454,n14455,n14456);
  nor U15166(n14456,n14457,n14458);
  and U15167(n14458,n14311,G36566);
  nor U15168(n14457,n12561,n14329);
  nand U15169(n14455,n14320,n12568);
  nand U15170(n14454,n14319,n12524);
  nand U15171(n14453,n14310,n14227);
  nand U15172(G7418,n14459,n14460,n14461,n14462);
  nor U15173(n14462,n14463,n14464);
  and U15174(n14464,n14311,G36565);
  nor U15175(n14463,n12673,n14329);
  nand U15176(n14461,n14320,n12894);
  nand U15177(n14459,n14310,n14236);
  nand U15178(G7417,n14465,n14466,n14467,n14468);
  nor U15179(n14468,n14469,n14470);
  and U15180(n14470,n14311,G36564);
  nor U15181(n14469,n12559,n14329);
  nand U15182(n14466,n14319,n12530);
  nand U15183(n14465,n14310,n14245);
  nand U15184(G7416,n14471,n14472,n14473,n14474);
  nor U15185(n14474,n14475,n14476);
  and U15186(n14476,n14311,G36563);
  nor U15187(n14475,n12783,n14329);
  nand U15188(n14472,n14319,n12533);
  nand U15189(n14471,n14310,n14254);
  nand U15190(G7415,n14477,n14478,n14479,n14480);
  nor U15191(n14480,n14481,n14482);
  and U15192(n14482,n14311,G36562);
  nor U15193(n14481,n12639,n14329);
  nand U15194(n14478,n14319,n12536);
  nand U15195(n14477,n14310,n12638);
  nand U15196(G7414,n14483,n14484,n14485,n14486);
  nor U15197(n14486,n14487,n14488);
  and U15198(n14488,n14311,G36561);
  nor U15199(n14487,n12782,n14329);
  nand U15200(n14485,n14320,n12870);
  nand U15201(n14484,n14319,n12539);
  nand U15202(n14483,n14310,n14269);
  nand U15203(G7413,n14489,n14490,n14491,n14492);
  nor U15204(n14492,n14493,n14494);
  and U15205(n14494,n14311,G36560);
  nor U15206(n14493,n12688,n14329);
  nand U15207(n14491,n14320,n12690);
  nand U15208(n14490,n14319,n12542);
  not U15209(n14319,n14438);
  nand U15210(n14438,n14314,n14278);
  nand U15211(n14489,n14310,n14277);
  nand U15212(G7412,n14495,n14496,n14497,n14498);
  nand U15213(n14498,n14310,n14296);
  nand U15214(n14497,n14320,n12810);
  not U15215(n14320,n14439);
  nand U15216(n14439,n14314,n14499);
  nand U15217(n14496,n14440,n12539);
  not U15218(n14440,n14329);
  nand U15219(n14329,n14314,n14297);
  not U15220(n14314,n14311);
  nand U15221(n14495,G36559,n14311);
  nand U15222(n14311,n14500,n14501,n14301);
  and U15223(n14301,n12923,n14502,n14503,n14504);
  nand U15224(n14501,n14505,n12952,n14303);
  nand U15225(n14505,n14506,n13029,n14507);
  nand U15226(n14507,n14284,n13025);
  nand U15227(n14500,n14302,n14304);
  not U15228(n14304,n14303);
  and U15229(n14302,n14508,n14509);
  or U15230(n14509,n13635,n12950);
  nand U15231(n13635,n14510,n13899);
  nand U15232(n14508,n13656,n13026);
  nand U15233(G7411,n14511,n14512,n14513);
  nand U15234(n14513,n14514,n13647);
  not U15235(n13647,n13011);
  nand U15236(n13011,n14515,n14516);
  nand U15237(n14511,n14517,G36558);
  nand U15238(G7410,n14518,n14512,n14519);
  nand U15239(n14519,n14514,n13007);
  and U15240(n13007,n14520,n14516);
  nand U15241(n14512,n14028,n14521);
  and U15242(n14028,n14522,n12449,n12934);
  nand U15243(n12449,n14523,n14524,n14525,n14526);
  nand U15244(n14525,G36622,n14527);
  nand U15245(n14524,G36590,n14528);
  nand U15246(n14523,G36558,n14529);
  nand U15247(n14522,n14530,n14531);
  nand U15248(n14531,n14532,n14533);
  nand U15249(n14518,n14517,G36557);
  nand U15250(G7409,n14534,n14535,n14536);
  nor U15251(n14536,n14537,n14538,n14539);
  and U15252(n14539,G36556,n14517);
  nor U15253(n14538,n14517,n14043);
  nand U15254(n14043,n14540,n12452,n14297);
  nand U15255(n12452,n14541,n14542,n14543,n14526);
  nand U15256(n14543,G36621,n14527);
  nand U15257(n14542,G36589,n14528);
  nand U15258(n14541,G36557,n14529);
  nand U15259(n14540,n14530,G36675);
  nor U15260(n14537,n12581,n14544);
  nand U15261(n14535,n14545,n13297);
  xor U15262(n13297,n13321,n14546);
  and U15263(n14546,n13320,n13306);
  nand U15264(n13306,n14547,n13313,n14548);
  nand U15265(n14548,n13322,n12663);
  nand U15266(n14547,n13322,n13318);
  not U15267(n13322,n13316);
  or U15268(n13320,n13316,n14549,n13313);
  xnor U15269(n13313,n14550,n14551);
  nor U15270(n14551,n14552,n14553,n14554,n14555);
  nor U15271(n14555,n14556,n12581);
  nor U15272(n14554,n12662,n14557);
  nor U15273(n14553,n12663,n14558);
  nor U15274(n14552,n13293,n14559);
  nor U15275(n14549,n13318,n12663);
  nand U15276(n13316,n14560,n14561,n14562,n14563);
  nor U15277(n14563,n14564,n14565);
  nor U15278(n14564,n12581,n14557);
  not U15279(n12581,n12458);
  nand U15280(n14562,n13286,n14566);
  nand U15281(n14561,n13012,n14567);
  or U15282(n14560,n14559,n12663);
  not U15283(n12663,n12455);
  nand U15284(n13321,n14568,n14569);
  nand U15285(n14569,n14570,n14571);
  nand U15286(n14534,n14514,n13012);
  not U15287(n13012,n13293);
  nand U15288(n13293,n14572,n14516);
  nand U15289(G7408,n14573,n14574,n14575,n14576);
  nor U15290(n14576,n14577,n14578);
  and U15291(n14578,G36555,n14517);
  nor U15292(n14577,n12905,n14544);
  not U15293(n12905,n12461);
  nand U15294(n14575,n14514,n13286);
  nand U15295(n14574,n14579,n12455);
  nand U15296(n12455,n14580,n14581,n14582,n14526);
  nand U15297(n14526,n14583,n14039,n14038);
  not U15298(n14039,G36697);
  nand U15299(n14582,G36620,n14527);
  nand U15300(n14581,G36588,n14528);
  nand U15301(n14580,G36556,n14529);
  nand U15302(n14573,n14545,n12664);
  xor U15303(n12664,n14571,n14584);
  and U15304(n14584,n14570,n14568);
  nand U15305(n14568,n14585,n14586);
  or U15306(n14570,n14585,n14586);
  nand U15307(n14586,n14587,n14588,n14589);
  nand U15308(n14588,n13286,n14590);
  nand U15309(n14587,n14591,n12458);
  xor U15310(n14585,n14592,n14593);
  and U15311(n14593,n14594,n14595);
  nand U15312(n14595,n13286,n14596);
  not U15313(n13286,n12662);
  nand U15314(n12662,n14597,n14516);
  nand U15315(n14594,n14590,n12458);
  nand U15316(n14571,n14598,n14599);
  nand U15317(n14599,n14600,n14601);
  nand U15318(G7407,n14602,n14603,n14604,n14605);
  nor U15319(n14605,n14606,n14607);
  and U15320(n14607,G36554,n14517);
  nor U15321(n14606,n12723,n14544);
  not U15322(n12723,n12464);
  nand U15323(n14604,n14514,n13287);
  nand U15324(n14603,n14579,n12458);
  nand U15325(n12458,n14608,n14609,n14610,n14611);
  nand U15326(n14611,n14052,n14583);
  xor U15327(n14052,n14038,G36697);
  nand U15328(n14610,G36619,n14527);
  nand U15329(n14609,G36587,n14528);
  nand U15330(n14608,G36555,n14529);
  nand U15331(n14602,n14545,n12583);
  xor U15332(n12583,n14601,n14612);
  and U15333(n14612,n14600,n14598);
  nand U15334(n14598,n14613,n14614);
  or U15335(n14600,n14613,n14614);
  nand U15336(n14614,n14615,n14616,n14589);
  nand U15337(n14616,n13287,n14590);
  nand U15338(n14615,n14591,n12461);
  xor U15339(n14613,n14592,n14617);
  and U15340(n14617,n14618,n14619);
  nand U15341(n14619,n13287,n14596);
  not U15342(n13287,n12580);
  nand U15343(n12580,n14620,n14516);
  nand U15344(n14618,n14590,n12461);
  nand U15345(n14601,n14621,n14622);
  nand U15346(n14622,n14623,n14624);
  nand U15347(G7406,n14625,n14626,n14627,n14628);
  nor U15348(n14628,n14629,n14630);
  and U15349(n14630,G36553,n14517);
  nor U15350(n14629,n12772,n14544);
  not U15351(n12772,n12467);
  nand U15352(n14627,n14514,n13274);
  nand U15353(n14626,n14579,n12461);
  nand U15354(n12461,n14631,n14632,n14633,n14634);
  nand U15355(n14634,n14583,n14635);
  not U15356(n14635,n12578);
  nor U15357(n12578,n14038,n14636);
  and U15358(n14636,G36703,n14637);
  nor U15359(n14038,n14637,G36703);
  nand U15360(n14633,G36618,n14527);
  nand U15361(n14632,G36586,n14528);
  nand U15362(n14631,G36554,n14529);
  nand U15363(n14625,n14545,n12906);
  xor U15364(n12906,n14624,n14638);
  and U15365(n14638,n14623,n14621);
  nand U15366(n14621,n14639,n14640);
  or U15367(n14623,n14639,n14640);
  nand U15368(n14640,n14641,n14642,n14589);
  nand U15369(n14642,n13274,n14590);
  nand U15370(n14641,n14591,n12464);
  xor U15371(n14639,n14592,n14643);
  and U15372(n14643,n14644,n14645);
  nand U15373(n14645,n13274,n14596);
  not U15374(n13274,n12904);
  nand U15375(n12904,n14646,n14516);
  nand U15376(n14644,n14590,n12464);
  nand U15377(n14624,n14647,n14648);
  nand U15378(n14648,n14649,n14650);
  nand U15379(G7405,n14651,n14652,n14653,n14654);
  nor U15380(n14654,n14655,n14656);
  and U15381(n14656,G36552,n14517);
  nor U15382(n14655,n12607,n14544);
  not U15383(n12607,n12470);
  nand U15384(n14653,n14514,n13275);
  nand U15385(n14652,n14579,n12464);
  nand U15386(n12464,n14657,n14658,n14659,n14660);
  nand U15387(n14660,n14583,n14068);
  nand U15388(n14068,n14637,n14661);
  nand U15389(n14661,G36677,n14662);
  or U15390(n14637,n14662,G36677);
  nand U15391(n14659,G36617,n14527);
  nand U15392(n14658,G36585,n14528);
  nand U15393(n14657,G36553,n14529);
  nand U15394(n14651,n14545,n12724);
  xor U15395(n12724,n14650,n14663);
  and U15396(n14663,n14649,n14647);
  nand U15397(n14647,n14664,n14665);
  or U15398(n14649,n14664,n14665);
  nand U15399(n14665,n14666,n14667,n14589);
  nand U15400(n14667,n13275,n14590);
  nand U15401(n14666,n14591,n12467);
  xor U15402(n14664,n14592,n14668);
  and U15403(n14668,n14669,n14670);
  nand U15404(n14670,n13275,n14596);
  not U15405(n13275,n12722);
  nand U15406(n12722,n14671,n14516);
  nand U15407(n14669,n14590,n12467);
  nand U15408(n14650,n14672,n14673);
  nand U15409(n14673,n14674,n14675);
  nand U15410(G7404,n14676,n14677,n14678,n14679);
  nor U15411(n14679,n14680,n14681);
  and U15412(n14681,G36551,n14517);
  nor U15413(n14680,n12846,n14544);
  not U15414(n12846,n12473);
  nand U15415(n14678,n14514,n13262);
  nand U15416(n14677,n14579,n12467);
  nand U15417(n12467,n14682,n14683,n14684,n14685);
  nand U15418(n14685,n14583,n14076);
  nand U15419(n14076,n14662,n14686);
  nand U15420(n14686,G36692,n14687);
  or U15421(n14662,n14687,G36692);
  nand U15422(n14684,G36616,n14527);
  nand U15423(n14683,G36584,n14528);
  nand U15424(n14682,G36552,n14529);
  nand U15425(n14676,n14545,n12773);
  xor U15426(n12773,n14675,n14688);
  and U15427(n14688,n14674,n14672);
  nand U15428(n14672,n14689,n14690);
  or U15429(n14674,n14689,n14690);
  nand U15430(n14690,n14691,n14692,n14589);
  nand U15431(n14692,n13262,n14590);
  nand U15432(n14691,n14591,n12470);
  xor U15433(n14689,n14592,n14693);
  and U15434(n14693,n14694,n14695);
  nand U15435(n14695,n13262,n14596);
  not U15436(n13262,n12771);
  nand U15437(n12771,n14696,n14516);
  nand U15438(n14694,n14590,n12470);
  nand U15439(n14675,n14697,n14698);
  nand U15440(n14698,n14699,n14700);
  nand U15441(G7403,n14701,n14702,n14703,n14704);
  nor U15442(n14704,n14705,n14706);
  and U15443(n14706,G36550,n14517);
  nor U15444(n14705,n12700,n14544);
  not U15445(n12700,n12476);
  nand U15446(n14703,n14514,n13263);
  nand U15447(n14702,n14579,n12470);
  nand U15448(n12470,n14707,n14708,n14709,n14710);
  nand U15449(n14710,n14583,n14084);
  nand U15450(n14084,n14687,n14711);
  nand U15451(n14711,G36688,n14712);
  or U15452(n14687,n14712,G36688);
  nand U15453(n14709,G36615,n14527);
  nand U15454(n14708,G36583,n14528);
  nand U15455(n14707,G36551,n14529);
  nand U15456(n14701,n14545,n12608);
  xor U15457(n12608,n14700,n14713);
  and U15458(n14713,n14699,n14697);
  nand U15459(n14697,n14714,n14715);
  or U15460(n14699,n14714,n14715);
  nand U15461(n14715,n14716,n14717,n14589);
  nand U15462(n14717,n13263,n14590);
  nand U15463(n14716,n14591,n12473);
  xor U15464(n14714,n14592,n14718);
  and U15465(n14718,n14719,n14720);
  nand U15466(n14720,n13263,n14596);
  not U15467(n13263,n12606);
  nand U15468(n12606,n14721,n14516);
  nand U15469(n14719,n14590,n12473);
  nand U15470(n14700,n14722,n14723);
  nand U15471(n14723,n14724,n14725);
  nand U15472(G7402,n14726,n14727,n14728,n14729);
  nor U15473(n14729,n14730,n14731);
  and U15474(n14731,G36549,n14517);
  nor U15475(n14730,n12821,n14544);
  not U15476(n12821,n12479);
  nand U15477(n14728,n14514,n13250);
  nand U15478(n14727,n14579,n12473);
  nand U15479(n12473,n14732,n14733,n14734,n14735);
  nand U15480(n14735,n14583,n14092);
  nand U15481(n14092,n14712,n14736);
  nand U15482(n14736,G36701,n14737);
  or U15483(n14712,n14737,G36701);
  nand U15484(n14734,G36614,n14527);
  nand U15485(n14733,G36582,n14528);
  nand U15486(n14732,G36550,n14529);
  nand U15487(n14726,n14545,n12847);
  xor U15488(n12847,n14725,n14738);
  and U15489(n14738,n14724,n14722);
  nand U15490(n14722,n14739,n14740);
  or U15491(n14724,n14739,n14740);
  nand U15492(n14740,n14741,n14742,n14589);
  nand U15493(n14742,n13250,n14590);
  nand U15494(n14741,n14591,n12476);
  xor U15495(n14739,n14592,n14743);
  and U15496(n14743,n14744,n14745);
  nand U15497(n14745,n13250,n14596);
  not U15498(n13250,n12845);
  nand U15499(n12845,n14746,n14516);
  nand U15500(n14744,n14590,n12476);
  nand U15501(n14725,n14747,n14748);
  nand U15502(n14748,n14749,n14750);
  nand U15503(G7401,n14751,n14752,n14753,n14754);
  nor U15504(n14754,n14755,n14756);
  and U15505(n14756,G36548,n14517);
  nor U15506(n14755,n12649,n14544);
  not U15507(n12649,n12482);
  nand U15508(n14753,n14514,n13251);
  nand U15509(n14752,n14579,n12476);
  nand U15510(n12476,n14757,n14758,n14759,n14760);
  nand U15511(n14760,n14583,n14100);
  nand U15512(n14100,n14737,n14761);
  nand U15513(n14761,G36682,n14762);
  or U15514(n14737,n14762,G36682);
  nand U15515(n14759,G36613,n14527);
  nand U15516(n14758,G36581,n14528);
  nand U15517(n14757,G36549,n14529);
  nand U15518(n14751,n14545,n12701);
  xor U15519(n12701,n14750,n14763);
  and U15520(n14763,n14749,n14747);
  nand U15521(n14747,n14764,n14765);
  or U15522(n14749,n14764,n14765);
  nand U15523(n14765,n14766,n14767,n14589);
  nand U15524(n14767,n13251,n14590);
  nand U15525(n14766,n14591,n12479);
  xor U15526(n14764,n14592,n14768);
  and U15527(n14768,n14769,n14770);
  nand U15528(n14770,n13251,n14596);
  not U15529(n13251,n12699);
  nand U15530(n12699,n14771,n14516);
  nand U15531(n14769,n14590,n12479);
  nand U15532(n14750,n14772,n14773);
  nand U15533(n14773,n14774,n14775);
  nand U15534(G7400,n14776,n14777,n14778,n14779);
  nor U15535(n14779,n14780,n14781);
  and U15536(n14781,G36547,n14517);
  nor U15537(n14780,n12879,n14544);
  not U15538(n12879,n12485);
  nand U15539(n14778,n14514,n13239);
  nand U15540(n14777,n14579,n12479);
  nand U15541(n12479,n14782,n14783,n14784,n14785);
  nand U15542(n14785,n14583,n14108);
  nand U15543(n14108,n14762,n14786);
  nand U15544(n14786,G36694,n14787);
  or U15545(n14762,n14787,G36694);
  nand U15546(n14784,G36612,n14527);
  nand U15547(n14783,G36580,n14528);
  nand U15548(n14782,G36548,n14529);
  nand U15549(n14776,n14545,n12822);
  xor U15550(n12822,n14775,n14788);
  and U15551(n14788,n14774,n14772);
  nand U15552(n14772,n14789,n14790);
  or U15553(n14774,n14789,n14790);
  nand U15554(n14790,n14791,n14792,n14589);
  nand U15555(n14792,n13239,n14590);
  nand U15556(n14791,n14591,n12482);
  xor U15557(n14789,n14793,n14550);
  nand U15558(n14793,n14794,n14795);
  nand U15559(n14795,n13239,n14596);
  not U15560(n13239,n12820);
  nand U15561(n12820,n14796,n14516);
  nand U15562(n14794,n14590,n12482);
  nand U15563(n14775,n14797,n14798);
  nand U15564(n14798,n14799,n14800);
  nand U15565(G7399,n14801,n14802,n14803,n14804);
  nor U15566(n14804,n14805,n14806);
  and U15567(n14806,G36546,n14517);
  nor U15568(n14805,n12648,n14544);
  not U15569(n12648,n12488);
  nand U15570(n14803,n14545,n12652);
  xor U15571(n12652,n14800,n14807);
  and U15572(n14807,n14799,n14797);
  nand U15573(n14797,n14808,n14809);
  or U15574(n14799,n14808,n14809);
  nand U15575(n14809,n14810,n14811,n14589);
  not U15576(n14589,n14565);
  nand U15577(n14565,n14812,n14813);
  nand U15578(n14813,n14814,G36578);
  nand U15579(n14812,n14815,G36610);
  nand U15580(n14811,n12653,n14590);
  nand U15581(n14810,n14591,n12485);
  xor U15582(n14808,n14816,n14550);
  nand U15583(n14816,n14817,n14818,n14819);
  nand U15584(n14819,n14590,n12485);
  nand U15585(n14818,n12971,n14820);
  nand U15586(n14817,n12653,n14596);
  not U15587(n12653,n13233);
  nand U15588(n13233,n14821,n14822);
  nand U15589(n14822,n14823,n13899);
  or U15590(n14821,n14824,n14823);
  nand U15591(n14800,n14825,n14826);
  nand U15592(n14826,n14827,n14828);
  nand U15593(n14802,n14514,n14124);
  nand U15594(n14124,n14829,n14830);
  nand U15595(n14830,n12971,n14831);
  nand U15596(n14829,n14824,n14516);
  nand U15597(n14801,n14579,n12482);
  nand U15598(n12482,n14832,n14833,n14834,n14835);
  nand U15599(n14835,n14583,n14116);
  nand U15600(n14116,n14787,n14836);
  nand U15601(n14836,G36684,n14837);
  or U15602(n14787,n14837,G36684);
  nand U15603(n14834,G36611,n14527);
  nand U15604(n14833,G36579,n14528);
  nand U15605(n14832,G36547,n14529);
  nand U15606(G7398,n14838,n14839,n14840,n14841);
  nor U15607(n14841,n14842,n14843);
  and U15608(n14843,G36545,n14517);
  nor U15609(n14842,n12733,n14544);
  not U15610(n12733,n12491);
  nand U15611(n14840,n14545,n12882);
  xor U15612(n12882,n14828,n14844);
  and U15613(n14844,n14827,n14825);
  nand U15614(n14825,n14845,n14846);
  or U15615(n14827,n14845,n14846);
  nand U15616(n14846,n14847,n14848,n14849,n14850);
  nand U15617(n14850,n12883,n14590);
  nand U15618(n14849,n14591,n12488);
  nand U15619(n14848,n14814,G36577);
  nand U15620(n14847,n14815,G36609);
  xor U15621(n14845,n14851,n14550);
  nand U15622(n14851,n14852,n14853,n14854);
  nand U15623(n14854,n14590,n12488);
  nand U15624(n14853,n12883,n14596);
  not U15625(n12883,n13230);
  nand U15626(n13230,n14855,n14856);
  or U15627(n14856,n14857,n14823);
  nand U15628(n14855,n13885,n14823);
  nand U15629(n14852,n13891,n14820);
  nand U15630(n14828,n14858,n14859);
  nand U15631(n14859,n14860,n14861);
  nand U15632(n14839,n14514,n14133);
  nand U15633(n14133,n14862,n14863);
  nand U15634(n14863,n13891,n14831);
  not U15635(n13891,n13885);
  nand U15636(n13885,n14864,n14865);
  or U15637(n14865,G36481,G36494);
  nand U15638(n14864,G36494,n14866);
  nand U15639(n14862,n14857,n14516);
  nand U15640(n14838,n14579,n12485);
  nand U15641(n12485,n14867,n14868,n14869,n14870);
  nand U15642(n14870,n14583,n14125);
  nand U15643(n14125,n14837,n14871);
  nand U15644(n14871,G36698,n14872);
  or U15645(n14837,n14872,G36698);
  or U15646(n14872,n14873,G36679);
  nand U15647(n14869,G36610,n14527);
  nand U15648(n14868,G36578,n14528);
  nand U15649(n14867,G36546,n14529);
  nand U15650(G7397,n14874,n14875,n14876,n14877);
  nor U15651(n14877,n14878,n14879);
  and U15652(n14879,G36544,n14517);
  nor U15653(n14878,n12758,n14544);
  not U15654(n12758,n12494);
  nand U15655(n14876,n14545,n12761);
  xor U15656(n12761,n14861,n14880);
  and U15657(n14880,n14860,n14858);
  nand U15658(n14858,n14881,n14882);
  or U15659(n14860,n14881,n14882);
  nand U15660(n14882,n14883,n14884,n14885,n14886);
  nand U15661(n14886,n12762,n14590);
  nand U15662(n14885,n14591,n12491);
  nand U15663(n14884,n14814,G36576);
  nand U15664(n14883,n14815,G36608);
  xor U15665(n14881,n14887,n14550);
  nand U15666(n14887,n14888,n14889,n14890);
  nand U15667(n14890,n14590,n12491);
  nand U15668(n14889,n12762,n14596);
  not U15669(n12762,n13221);
  nand U15670(n13221,n14891,n14892);
  nand U15671(n14892,n14823,n13873);
  or U15672(n14891,n14893,n14823);
  nand U15673(n14888,n13878,n14820);
  nand U15674(n14861,n14894,n14895);
  nand U15675(n14895,n14896,n14897);
  nand U15676(n14875,n14514,n14141);
  nand U15677(n14141,n14898,n14899);
  nand U15678(n14899,n13878,n14831);
  not U15679(n13878,n13873);
  nand U15680(n13873,n14900,n14901,n14902);
  nand U15681(n14901,n14903,n14904);
  nand U15682(n14900,G36480,n14905,G36494);
  nand U15683(n14898,n14893,n14516);
  nand U15684(n14874,n14579,n12488);
  nand U15685(n12488,n14906,n14907,n14908,n14909);
  nand U15686(n14909,n14910,n14583);
  not U15687(n14910,n12880);
  xor U15688(n12880,n14873,G36679);
  nand U15689(n14908,G36609,n14527);
  nand U15690(n14907,G36577,n14528);
  nand U15691(n14906,G36545,n14529);
  nand U15692(G7396,n14911,n14912,n14913,n14914);
  nor U15693(n14914,n14915,n14916);
  and U15694(n14916,G36543,n14517);
  nor U15695(n14915,n12593,n14544);
  not U15696(n12593,n12497);
  nand U15697(n14913,n14545,n12736);
  xor U15698(n12736,n14897,n14917);
  and U15699(n14917,n14896,n14894);
  nand U15700(n14894,n14918,n14919);
  or U15701(n14896,n14918,n14919);
  nand U15702(n14919,n14920,n14921,n14922,n14923);
  nand U15703(n14923,n12737,n14590);
  nand U15704(n14922,n14591,n12494);
  nand U15705(n14921,n14814,G36575);
  nand U15706(n14920,n14815,G36607);
  xor U15707(n14918,n14924,n14550);
  nand U15708(n14924,n14925,n14926,n14927);
  nand U15709(n14927,n14590,n12494);
  nand U15710(n14926,n12737,n14596);
  not U15711(n12737,n13218);
  nand U15712(n13218,n14928,n14929);
  or U15713(n14929,n14930,n14823);
  nand U15714(n14928,n13861,n14823);
  nand U15715(n14925,n13864,n14820);
  nand U15716(n14897,n14931,n14932);
  nand U15717(n14932,n14933,n14934);
  nand U15718(n14912,n14514,n14150);
  nand U15719(n14150,n14935,n14936);
  nand U15720(n14936,n13864,n14831);
  not U15721(n13864,n13861);
  nand U15722(n13861,n14937,n14938);
  or U15723(n14938,G36479,G36494);
  nand U15724(n14937,G36494,n14939);
  nand U15725(n14935,n14930,n14516);
  nand U15726(n14911,n14579,n12491);
  nand U15727(n12491,n14940,n14941,n14942,n14943);
  nand U15728(n14943,n14583,n14142);
  nand U15729(n14142,n14944,n14873);
  or U15730(n14873,n14945,G36689);
  nand U15731(n14944,G36689,n14945);
  nand U15732(n14942,G36608,n14527);
  nand U15733(n14941,G36576,n14528);
  nand U15734(n14940,G36544,n14529);
  nand U15735(G7395,n14946,n14947,n14948,n14949);
  nor U15736(n14949,n14950,n14951);
  and U15737(n14951,G36542,n14517);
  nor U15738(n14950,n12832,n14544);
  not U15739(n12832,n12500);
  nand U15740(n14948,n14545,n12938);
  xor U15741(n12938,n14934,n14952);
  and U15742(n14952,n14933,n14931);
  nand U15743(n14931,n14953,n14954);
  or U15744(n14933,n14953,n14954);
  nand U15745(n14954,n14955,n14956,n14957,n14958);
  nand U15746(n14958,n12954,n14590);
  nand U15747(n14957,n14591,n12497);
  nand U15748(n14956,n14814,G36574);
  nand U15749(n14955,n14815,G36606);
  xor U15750(n14953,n14959,n14550);
  nand U15751(n14959,n14960,n14961,n14962);
  nand U15752(n14962,n14590,n12497);
  nand U15753(n14961,n12954,n14596);
  not U15754(n12954,n13209);
  nand U15755(n13209,n14963,n14964);
  nand U15756(n14964,n14823,n13850);
  or U15757(n14963,n14965,n14823);
  nand U15758(n14960,n13855,n14820);
  nand U15759(n14934,n14966,n14967);
  nand U15760(n14967,n14968,n14969);
  nand U15761(n14947,n14514,n14159);
  nand U15762(n14159,n14970,n14971);
  nand U15763(n14971,n13855,n14831);
  not U15764(n13855,n13850);
  nand U15765(n13850,n14972,n14973,n14974);
  nand U15766(n14973,n14975,n14904);
  nand U15767(n14972,G36478,n14976,G36494);
  nand U15768(n14970,n14965,n14516);
  nand U15769(n14946,n14579,n12494);
  nand U15770(n12494,n14977,n14978,n14979,n14980);
  nand U15771(n14980,n14583,n14151);
  nand U15772(n14151,n14945,n14981);
  nand U15773(n14981,G36691,n14982);
  or U15774(n14945,n14982,G36691);
  nand U15775(n14979,G36607,n14527);
  nand U15776(n14978,G36575,n14528);
  nand U15777(n14977,G36543,n14529);
  nand U15778(G7394,n14983,n14984,n14985,n14986);
  nor U15779(n14986,n14987,n14988);
  and U15780(n14988,G36541,n14517);
  nor U15781(n14987,n12592,n14544);
  not U15782(n12592,n12503);
  nand U15783(n14985,n14545,n12596);
  xor U15784(n12596,n14969,n14989);
  and U15785(n14989,n14966,n14968);
  or U15786(n14968,n14990,n14991);
  nand U15787(n14966,n14990,n14991);
  nand U15788(n14991,n14992,n14993,n14994,n14995);
  nand U15789(n14995,n12597,n14590);
  nand U15790(n14994,n14591,n12500);
  nand U15791(n14993,n14814,G36573);
  nand U15792(n14992,n14815,G36605);
  xor U15793(n14990,n14996,n14550);
  nand U15794(n14996,n14997,n14998,n14999);
  nand U15795(n14999,n14590,n12500);
  nand U15796(n14998,n12597,n14596);
  not U15797(n12597,n13206);
  nand U15798(n13206,n15000,n15001);
  nand U15799(n15001,n15002,n14516);
  nand U15800(n15000,n13838,n14823);
  nand U15801(n14997,n13841,n14820);
  nand U15802(n14969,n15003,n15004);
  nand U15803(n15004,n15005,n15006);
  nand U15804(n14984,n14514,n14168);
  nand U15805(n14168,n15007,n15008);
  nand U15806(n15008,n13841,n14831);
  not U15807(n13841,n13838);
  nand U15808(n13838,n15009,n15010);
  or U15809(n15010,G36477,G36494);
  nand U15810(n15009,G36494,n15011);
  nand U15811(n15007,n15012,n14516);
  nand U15812(n14983,n14579,n12497);
  nand U15813(n12497,n15013,n15014,n15015,n15016);
  nand U15814(n15016,n14583,n14160);
  nand U15815(n14160,n14982,n15017);
  nand U15816(n15017,G36676,n15018);
  or U15817(n15018,n15019,G36702);
  or U15818(n14982,G36676,G36702,n15019);
  nand U15819(n15015,G36606,n14527);
  nand U15820(n15014,G36574,n14528);
  nand U15821(n15013,G36542,n14529);
  nand U15822(G7393,n15020,n15021,n15022,n15023);
  nor U15823(n15023,n15024,n15025);
  and U15824(n15025,G36540,n14517);
  nor U15825(n15024,n12831,n14544);
  not U15826(n12831,n12506);
  nand U15827(n15022,n14545,n12835);
  xor U15828(n12835,n15006,n15026);
  and U15829(n15026,n15005,n15003);
  nand U15830(n15003,n15027,n15028);
  or U15831(n15005,n15027,n15028);
  nand U15832(n15028,n15029,n15030,n15031,n15032);
  nand U15833(n15032,n12836,n14590);
  nand U15834(n15031,n14591,n12503);
  nand U15835(n15030,n14814,G36572);
  nand U15836(n15029,n14815,G36604);
  xor U15837(n15027,n15033,n14550);
  nand U15838(n15033,n15034,n15035,n15036);
  nand U15839(n15036,n14590,n12503);
  nand U15840(n15035,n12836,n14596);
  not U15841(n12836,n13197);
  nand U15842(n13197,n15037,n15038);
  nand U15843(n15038,n14823,n13826);
  or U15844(n15037,n15039,n14823);
  nand U15845(n15034,n13831,n14820);
  nand U15846(n15006,n15040,n15041);
  nand U15847(n15041,n15042,n15043);
  nand U15848(n15021,n14514,n14176);
  nand U15849(n14176,n15044,n15045);
  nand U15850(n15045,n13831,n14831);
  not U15851(n13831,n13826);
  nand U15852(n13826,n15046,n15047,n15048);
  nand U15853(n15047,n15049,n14904);
  nand U15854(n15046,G36476,n15050,G36494);
  nand U15855(n15044,n15039,n14516);
  nand U15856(n15020,n14579,n12500);
  nand U15857(n12500,n15051,n15052,n15053,n15054);
  nand U15858(n15054,n15055,n14583);
  not U15859(n15055,n12594);
  xor U15860(n12594,n15019,G36702);
  nand U15861(n15053,G36605,n14527);
  nand U15862(n15052,G36573,n14528);
  nand U15863(n15051,G36541,n14529);
  nand U15864(G7392,n15056,n15057,n15058,n15059);
  nor U15865(n15059,n15060,n15061);
  and U15866(n15061,G36539,n14517);
  nor U15867(n15060,n12618,n14544);
  not U15868(n12618,n12509);
  nand U15869(n15058,n14545,n12712);
  xor U15870(n12712,n15043,n15062);
  and U15871(n15062,n15042,n15040);
  nand U15872(n15040,n15063,n15064);
  or U15873(n15042,n15063,n15064);
  nand U15874(n15064,n15065,n15066,n15067,n15068);
  nand U15875(n15068,n12713,n14590);
  nand U15876(n15067,n14591,n12506);
  nand U15877(n15066,n14814,G36571);
  nand U15878(n15065,n14815,G36603);
  xor U15879(n15063,n15069,n14550);
  nand U15880(n15069,n15070,n15071,n15072);
  nand U15881(n15072,n14590,n12506);
  nand U15882(n15071,n12713,n14596);
  not U15883(n12713,n13194);
  nand U15884(n13194,n15073,n15074);
  or U15885(n15074,n15075,n14823);
  nand U15886(n15073,n13815,n14823);
  nand U15887(n15070,n13818,n14820);
  nand U15888(n15043,n15076,n15077);
  or U15889(n15077,n15078,n15079);
  nand U15890(n15057,n14514,n14185);
  nand U15891(n14185,n15080,n15081);
  nand U15892(n15081,n13818,n14831);
  not U15893(n13818,n13815);
  nand U15894(n13815,n15082,n15083);
  or U15895(n15083,G36475,G36494);
  nand U15896(n15082,G36494,n15084);
  nand U15897(n15080,n15075,n14516);
  nand U15898(n15056,n14579,n12503);
  nand U15899(n12503,n15085,n15086,n15087,n15088);
  nand U15900(n15088,n14583,n14177);
  nand U15901(n14177,n15019,n15089);
  nand U15902(n15089,G36683,n15090);
  or U15903(n15090,n15091,G36693);
  or U15904(n15019,G36683,G36693,n15091);
  nand U15905(n15087,G36604,n14527);
  nand U15906(n15086,G36572,n14528);
  nand U15907(n15085,G36540,n14529);
  nand U15908(G7391,n15092,n15093,n15094,n15095);
  nor U15909(n15095,n15096,n15097);
  and U15910(n15097,G36538,n14517);
  nor U15911(n15096,n12796,n14544);
  not U15912(n12796,n12512);
  nand U15913(n15094,n14545,n12858);
  xnor U15914(n12858,n15079,n15098);
  nor U15915(n15098,n15078,n15099);
  not U15916(n15099,n15076);
  nand U15917(n15076,n15100,n15101);
  nor U15918(n15078,n15100,n15101);
  nand U15919(n15101,n15102,n15103,n15104,n15105);
  nand U15920(n15105,n12859,n14590);
  nand U15921(n15104,n14591,n12509);
  nand U15922(n15103,n14814,G36570);
  nand U15923(n15102,n14815,G36602);
  xor U15924(n15100,n15106,n14550);
  nand U15925(n15106,n15107,n15108,n15109);
  nand U15926(n15109,n14590,n12509);
  nand U15927(n15108,n12859,n14596);
  not U15928(n12859,n13184);
  nand U15929(n13184,n15110,n15111);
  nand U15930(n15111,n14823,n13804);
  or U15931(n15110,n15112,n14823);
  nand U15932(n15107,n13809,n14820);
  nand U15933(n15093,n14514,n14193);
  nand U15934(n14193,n15113,n15114);
  nand U15935(n15114,n13809,n14831);
  not U15936(n13809,n13804);
  nand U15937(n13804,n15115,n15116,n15117);
  nand U15938(n15116,n15118,n14904);
  nand U15939(n15115,G36474,n15119,G36494);
  nand U15940(n15113,n15112,n14516);
  nand U15941(n15092,n14579,n12506);
  nand U15942(n12506,n15120,n15121,n15122,n15123);
  nand U15943(n15123,n15124,n14583);
  not U15944(n15124,n12710);
  xor U15945(n12710,n15091,G36693);
  nand U15946(n15122,G36603,n14527);
  nand U15947(n15121,G36571,n14528);
  nand U15948(n15120,G36539,n14529);
  nand U15949(G7390,n15125,n15126,n15127,n15128);
  nand U15950(n15128,n14579,n12509);
  nand U15951(n12509,n15129,n15130,n15131,n15132);
  nand U15952(n15132,n14583,n14194);
  nand U15953(n14194,n15091,n15133);
  nand U15954(n15133,G36681,n15134);
  nand U15955(n15134,n15135,n13792);
  nand U15956(n15091,n15136,n13792,n15135);
  not U15957(n13792,G36700);
  not U15958(n15136,G36681);
  nand U15959(n15131,G36602,n14527);
  nand U15960(n15130,G36570,n14528);
  nand U15961(n15129,G36538,n14529);
  nor U15962(n15127,n15137,n15138);
  nor U15963(n15138,n13181,n15139);
  not U15964(n13181,n12623);
  nand U15965(n12623,n15140,n15141);
  nand U15966(n15141,n15142,n15143);
  nand U15967(n15142,n15144,n15145);
  nand U15968(n15140,n15079,n15144);
  and U15969(n15079,n15145,n15146);
  nand U15970(n15146,n15143,n15144);
  nand U15971(n15144,n15147,n15148);
  not U15972(n15148,n15149);
  xor U15973(n15147,n15150,n14592);
  nand U15974(n15143,n15151,n15152);
  nand U15975(n15152,n15153,n15154);
  nand U15976(n15145,n15155,n15149);
  nand U15977(n15149,n15156,n15157,n15158,n15159);
  nand U15978(n15159,n12624,n14590);
  nand U15979(n15158,n14591,n12512);
  nand U15980(n15157,n14814,G36569);
  nand U15981(n15156,n14815,G36601);
  xor U15982(n15155,n14550,n15150);
  nand U15983(n15150,n15160,n15161,n15162);
  nand U15984(n15162,n14590,n12512);
  nand U15985(n15161,n12624,n14596);
  not U15986(n12624,n13185);
  nand U15987(n13185,n15163,n15164);
  nand U15988(n15164,n15165,n14516);
  nand U15989(n15163,n13938,n14823);
  nand U15990(n15160,n13798,n14820);
  and U15991(n15137,n12621,n14514);
  nand U15992(n12621,n15166,n15167);
  nand U15993(n15167,n13798,n14831);
  not U15994(n13798,n13938);
  nand U15995(n13938,n15168,n15169);
  or U15996(n15169,G36473,G36494);
  nand U15997(n15168,G36494,n15170);
  nand U15998(n15166,n15171,n14516);
  nand U15999(n15126,n15172,n12515);
  nand U16000(n15125,n14517,G36537);
  nand U16001(G7389,n15173,n15174,n15175,n15176);
  nor U16002(n15176,n15177,n15178);
  and U16003(n15178,G36536,n14517);
  nor U16004(n15177,n12561,n14544);
  not U16005(n12561,n12518);
  nand U16006(n15175,n14545,n12799);
  xor U16007(n12799,n15154,n15179);
  and U16008(n15179,n15153,n15151);
  nand U16009(n15151,n15180,n15181);
  or U16010(n15153,n15180,n15181);
  nand U16011(n15181,n15182,n15183,n15184,n15185);
  nand U16012(n15185,n12800,n14590);
  nand U16013(n15184,n14591,n12515);
  nand U16014(n15183,n14814,G36568);
  nand U16015(n15182,n14815,G36600);
  xor U16016(n15180,n15186,n14550);
  nand U16017(n15186,n15187,n15188,n15189);
  nand U16018(n15189,n14590,n12515);
  nand U16019(n15188,n12800,n14596);
  not U16020(n12800,n13172);
  nand U16021(n13172,n15190,n15191);
  nand U16022(n15191,n14823,n13779);
  or U16023(n15190,n15192,n14823);
  nand U16024(n15187,n13784,n14820);
  nand U16025(n15154,n15193,n15194);
  nand U16026(n15194,n15195,n15196);
  nand U16027(n15174,n14514,n14211);
  nand U16028(n14211,n15197,n15198);
  nand U16029(n15198,n13784,n14831);
  not U16030(n13784,n13779);
  nand U16031(n13779,n15199,n15200,n15201);
  nand U16032(n15200,n15202,n14904);
  nand U16033(n15199,G36472,n15203,G36494);
  nand U16034(n15197,n15192,n14516);
  nand U16035(n15173,n14579,n12512);
  nand U16036(n12512,n15204,n15205,n15206,n15207);
  nand U16037(n15207,n12620,n14583);
  xor U16038(n12620,n15135,G36700);
  nand U16039(n15206,G36601,n14527);
  nand U16040(n15205,G36569,n14528);
  nand U16041(n15204,G36537,n14529);
  nand U16042(G7388,n15208,n15209,n15210,n15211);
  nor U16043(n15211,n15212,n15213);
  and U16044(n15213,G36535,n14517);
  nor U16045(n15212,n12673,n14544);
  not U16046(n12673,n12521);
  nand U16047(n15210,n14545,n12676);
  xor U16048(n12676,n15196,n15214);
  and U16049(n15214,n15195,n15193);
  nand U16050(n15193,n15215,n15216);
  or U16051(n15195,n15215,n15216);
  nand U16052(n15216,n15217,n15218,n15219,n15220);
  nand U16053(n15220,n12677,n14590);
  nand U16054(n15219,n14591,n12518);
  nand U16055(n15218,n14814,G36567);
  nand U16056(n15217,n14815,G36599);
  xor U16057(n15215,n15221,n14550);
  nand U16058(n15221,n15222,n15223,n15224);
  nand U16059(n15224,n14590,n12518);
  nand U16060(n15223,n12677,n14596);
  not U16061(n12677,n13169);
  nand U16062(n13169,n15225,n15226);
  or U16063(n15226,n15227,n14823);
  nand U16064(n15225,n13767,n14823);
  nand U16065(n15222,n13770,n14820);
  nand U16066(n15196,n15228,n15229);
  nand U16067(n15229,n15230,n15231);
  nand U16068(n15209,n14514,n14219);
  nand U16069(n14219,n15232,n15233);
  nand U16070(n15233,n13770,n14831);
  not U16071(n13770,n13767);
  nand U16072(n13767,n15234,n15235);
  or U16073(n15235,G36471,G36494);
  nand U16074(n15234,G36494,n15236);
  nand U16075(n15232,n15227,n14516);
  nand U16076(n15208,n14579,n12515);
  nand U16077(n12515,n15237,n15238,n15239,n15240);
  not U16078(n15241,n12797);
  nor U16079(n12797,n15135,n15242);
  and U16080(n15242,G36686,n15243);
  nor U16081(n15135,n15243,G36686);
  or U16082(n15243,n15244,G36696);
  nand U16083(n15239,G36600,n14527);
  nand U16084(n15238,G36568,n14528);
  nand U16085(n15237,G36536,n14529);
  nand U16086(G7387,n15245,n15246,n15247,n15248);
  nor U16087(n15248,n15249,n15250);
  and U16088(n15250,G36534,n14517);
  nor U16089(n15249,n12559,n14544);
  not U16090(n12559,n12524);
  nand U16091(n15247,n14545,n12568);
  xor U16092(n12568,n15231,n15251);
  and U16093(n15251,n15230,n15228);
  nand U16094(n15228,n15252,n15253);
  or U16095(n15230,n15252,n15253);
  nand U16096(n15253,n15254,n15255,n15256,n15257);
  nand U16097(n15257,n12570,n14590);
  nand U16098(n15256,n14591,n12521);
  nand U16099(n15255,n14814,G36566);
  nand U16100(n15254,n14815,G36598);
  xor U16101(n15252,n14550,n15258);
  nand U16102(n15258,n15259,n15260,n15261);
  nand U16103(n15261,n14590,n12521);
  nand U16104(n15260,n12570,n14596);
  not U16105(n12570,n13160);
  nand U16106(n13160,n15262,n15263);
  nand U16107(n15263,n14823,n13756);
  or U16108(n15262,n15264,n14823);
  nand U16109(n15259,n13761,n14820);
  nand U16110(n15231,n15265,n15266);
  nand U16111(n15266,n15267,n15268);
  nand U16112(n15246,n14514,n14227);
  nand U16113(n14227,n15269,n15270);
  nand U16114(n15270,n13761,n14831);
  not U16115(n13761,n13756);
  nand U16116(n13756,n15271,n15272,n15273);
  nand U16117(n15272,n15274,n14904);
  nand U16118(n15271,G36470,n15275,G36494);
  nand U16119(n15269,n15264,n14516);
  nand U16120(n15245,n14579,n12518);
  nand U16121(n12518,n15276,n15277,n15278,n15279);
  nand U16122(n15279,n15280,n14583);
  not U16123(n15280,n12674);
  xor U16124(n12674,G36696,n15244);
  nand U16125(n15278,G36599,n14527);
  nand U16126(n15277,G36567,n14528);
  nand U16127(n15276,G36535,n14529);
  nand U16128(G7386,n15281,n15282,n15283,n15284);
  nor U16129(n15284,n15285,n15286);
  and U16130(n15286,G36533,n14517);
  nor U16131(n15285,n12783,n14544);
  not U16132(n12783,n12527);
  nand U16133(n15283,n14545,n12894);
  xor U16134(n12894,n15267,n15287);
  and U16135(n15287,n15265,n15268);
  or U16136(n15268,n15288,n15289);
  nand U16137(n15265,n15288,n15289);
  nand U16138(n15289,n15290,n15291,n15292,n15293);
  nand U16139(n15293,n12895,n14590);
  nand U16140(n15292,n14591,n12524);
  nand U16141(n15291,n14814,G36565);
  nand U16142(n15290,n14815,G36597);
  xor U16143(n15288,n15294,n14550);
  nand U16144(n15294,n15295,n15296,n15297);
  nand U16145(n15297,n14590,n12524);
  nand U16146(n15296,n12895,n14596);
  not U16147(n12895,n13157);
  nand U16148(n13157,n15298,n15299);
  nand U16149(n15299,n15300,n14516);
  nand U16150(n15298,n14823,n13745);
  nand U16151(n15295,n13748,n14820);
  nand U16152(n15267,n15301,n15302);
  nand U16153(n15302,n15303,n15304);
  nand U16154(n15282,n14514,n14236);
  nand U16155(n14236,n15305,n15306);
  nand U16156(n15306,n13748,n14831);
  not U16157(n13748,n13745);
  nand U16158(n13745,n15307,n15308);
  or U16159(n15308,G36469,G36494);
  nand U16160(n15307,G36494,n15309);
  nand U16161(n15305,n15310,n14516);
  nand U16162(n12521,n15311,n15312,n15313,n15314);
  nand U16163(n14228,n15315,n15244);
  or U16164(n15244,n15316,G36704);
  nand U16165(n15315,G36704,n15316);
  nand U16166(n15313,G36598,n14527);
  nand U16167(n15312,G36566,n14528);
  nand U16168(n15311,G36534,n14529);
  nand U16169(G7385,n15317,n15318,n15319,n15320);
  nor U16170(n15320,n15321,n15322);
  and U16171(n15322,G36532,n14517);
  nor U16172(n15321,n12639,n14544);
  not U16173(n12639,n12530);
  xor U16174(n12748,n15304,n15323);
  and U16175(n15323,n15303,n15301);
  nand U16176(n15301,n15324,n15325);
  or U16177(n15303,n15324,n15325);
  nand U16178(n15325,n15326,n15327,n15328,n15329);
  nand U16179(n15329,n12749,n14590);
  nand U16180(n15327,n14814,G36564);
  nand U16181(n15326,n14815,G36596);
  xor U16182(n15324,n15330,n14550);
  nand U16183(n15330,n15331,n15332,n15333);
  nand U16184(n15333,n14590,n12527);
  nand U16185(n15332,n12749,n14596);
  not U16186(n12749,n13148);
  nand U16187(n13148,n15334,n15335);
  nand U16188(n15335,n15336,n14516);
  nand U16189(n15334,n14823,n13734);
  nand U16190(n15331,n13739,n14820);
  nand U16191(n15304,n15337,n15338);
  nand U16192(n15338,n15339,n15340);
  nand U16193(n15318,n14514,n14245);
  nand U16194(n14245,n15341,n15342);
  nand U16195(n15342,n13739,n14831);
  not U16196(n13739,n13734);
  nand U16197(n13734,n15343,n15344,n15345);
  nand U16198(n15344,n15346,n14904);
  nand U16199(n15343,G36468,n15347,G36494);
  nand U16200(n15341,n15348,n14516);
  nand U16201(n15317,n14579,n12524);
  nand U16202(n12524,n15349,n15350,n15351,n15352);
  nand U16203(n14237,n15316,n15353);
  nand U16204(n15353,G36678,n15354);
  or U16205(n15316,n15354,G36678);
  nand U16206(n15351,G36597,n14527);
  nand U16207(n15350,G36565,n14528);
  nand U16208(n15349,G36533,n14529);
  nand U16209(G7384,n15355,n15356,n15357,n15358);
  nor U16210(n15358,n15359,n15360);
  and U16211(n15360,G36531,n14517);
  nor U16212(n15359,n12782,n14544);
  not U16213(n12782,n12533);
  xor U16214(n12786,n15340,n15361);
  and U16215(n15361,n15339,n15337);
  nand U16216(n15337,n15362,n15363);
  or U16217(n15339,n15362,n15363);
  nand U16218(n15363,n15364,n15365,n15366,n15367);
  nand U16219(n15367,n12787,n14590);
  nand U16220(n15365,n14814,G36563);
  nand U16221(n15364,n14815,G36595);
  xor U16222(n15362,n15368,n14550);
  nand U16223(n15368,n15369,n15370,n15371);
  nand U16224(n15371,n14590,n12530);
  nand U16225(n15370,n12787,n14596);
  not U16226(n12787,n13134);
  nand U16227(n13134,n15372,n15373);
  nand U16228(n15373,n15374,n14516);
  nand U16229(n15372,n13722,n14823);
  nand U16230(n15369,n13725,n14820);
  nand U16231(n15340,n15375,n15376);
  nand U16232(n15376,n15377,n15378);
  nand U16233(n15356,n14514,n14254);
  nand U16234(n14254,n15379,n15380);
  nand U16235(n15380,n13725,n14831);
  not U16236(n13725,n13722);
  nand U16237(n13722,n15381,n15382);
  or U16238(n15382,G36467,G36494);
  nand U16239(n15381,G36494,n15383);
  nand U16240(n15379,n15384,n14516);
  nand U16241(n15355,n14579,n12527);
  nand U16242(n12527,n15385,n15386,n15387,n15388);
  nand U16243(n14246,n15354,n15389);
  nand U16244(n15389,G36690,n15390);
  or U16245(n15390,G36699,G36687);
  or U16246(n15354,G36690,G36699,G36687);
  nand U16247(n15387,G36596,n14527);
  nand U16248(n15386,G36564,n14528);
  nand U16249(n15385,G36532,n14529);
  nand U16250(G7383,n15391,n15392,n15393,n15394);
  nor U16251(n15394,n15395,n15396);
  and U16252(n15396,G36530,n14517);
  nor U16253(n15395,n12688,n14544);
  xor U16254(n13133,n15378,n15397);
  and U16255(n15397,n15377,n15375);
  nand U16256(n15375,n15398,n15399);
  or U16257(n15377,n15398,n15399);
  nand U16258(n15399,n15400,n15401,n15402,n15403);
  nand U16259(n15403,n13135,n14590);
  nand U16260(n15401,n14814,G36562);
  nand U16261(n15400,n14815,G36594);
  xor U16262(n15398,n15404,n14550);
  nand U16263(n15404,n15405,n15406,n15407);
  nand U16264(n15407,n14590,n12533);
  nand U16265(n15406,n13135,n14596);
  not U16266(n13135,n12633);
  nand U16267(n12633,n15408,n15409);
  nand U16268(n15409,n14823,n13710);
  or U16269(n15408,n15410,n14823);
  nand U16270(n15405,n13715,n14820);
  nand U16271(n15378,n15411,n15412);
  nand U16272(n15412,n15413,n15414);
  nand U16273(n15392,n14514,n12638);
  nand U16274(n12638,n15415,n15416);
  nand U16275(n15416,n13715,n14831);
  not U16276(n13715,n13710);
  nand U16277(n13710,n15417,n15418,n15419);
  nand U16278(n15418,n15420,n14904);
  nand U16279(n15417,G36466,n15421,G36494);
  nand U16280(n15415,n15410,n14516);
  nand U16281(n15391,n14579,n12530);
  nand U16282(n12530,n15422,n15423,n15424,n15425);
  nand U16283(n15425,n15426,n14583);
  not U16284(n15426,n12784);
  xor U16285(n12784,G36687,G36699);
  nand U16286(n15424,G36595,n14527);
  nand U16287(n15423,G36563,n14528);
  nand U16288(n15422,G36531,n14529);
  nand U16289(G7382,n15427,n15428,n15429,n15430);
  nor U16290(n15430,n15431,n15432);
  and U16291(n15432,G36529,n14517);
  nor U16292(n15431,n12809,n14544);
  not U16293(n12809,n12539);
  nand U16294(n15429,n14545,n12870);
  xor U16295(n12870,n15413,n15433);
  and U16296(n15433,n15411,n15414);
  or U16297(n15414,n15434,n15435);
  nand U16298(n15411,n15434,n15435);
  nand U16299(n15435,n15436,n15437,n15438,n15439);
  nand U16300(n15439,n12869,n14590);
  nand U16301(n15438,n14591,n12536);
  nand U16302(n15437,n14814,G36561);
  nand U16303(n15436,n14815,G36593);
  xor U16304(n15434,n15440,n14550);
  nand U16305(n15440,n15441,n15442,n15443);
  nand U16306(n15443,n14590,n12536);
  nand U16307(n15442,n12869,n14596);
  not U16308(n12869,n13125);
  nand U16309(n13125,n15444,n15445);
  or U16310(n15445,n15446,n14823);
  nand U16311(n15444,n13698,n14823);
  nand U16312(n15441,n13700,n14820);
  nand U16313(n15413,n15447,n15448);
  nand U16314(n15448,n15449,n15450);
  nand U16315(n15428,n14514,n14269);
  nand U16316(n14269,n15451,n15452);
  nand U16317(n15452,n13700,n14831);
  not U16318(n13700,n13698);
  nand U16319(n13698,n15453,n15454);
  or U16320(n15454,G36465,G36494);
  nand U16321(n15453,G36494,n15455);
  nand U16322(n15451,n15446,n14516);
  nand U16323(n15427,n14579,n12533);
  nand U16324(n12533,n15456,n15457,n15458,n15459);
  nand U16325(n15459,G36594,n14527);
  nand U16326(n15458,G36562,n14528);
  nand U16327(n15457,G36530,n14529);
  nand U16328(n15456,n14583,n12637);
  not U16329(n12637,G36699);
  nand U16330(G7381,n15460,n15461,n15462,n15463);
  nor U16331(n15463,n15464,n15465);
  and U16332(n15465,G36528,n14517);
  nor U16333(n15464,n12688,n15466);
  not U16334(n12688,n12536);
  nand U16335(n12536,n15467,n15468,n15469,n15470);
  nand U16336(n15470,G36593,n14527);
  nand U16337(n15469,G36561,n14528);
  nand U16338(n15468,G36529,n14529);
  nand U16339(n15467,G36680,n14583);
  nand U16340(n15462,n15172,n12542);
  not U16341(n15172,n14544);
  nand U16342(n14544,n14278,n14521);
  and U16343(n14278,n12934,n12916);
  nand U16344(n12916,n15471,n15472);
  nand U16345(n15472,n15473,n15474);
  nand U16346(n15471,G36491,n15475);
  nand U16347(n15461,n14514,n14277);
  nand U16348(n14277,n15476,n15477);
  nand U16349(n15477,n13689,n14831);
  nand U16350(n15460,n14545,n12690);
  xor U16351(n12690,n15450,n15478);
  and U16352(n15478,n15449,n15447);
  nand U16353(n15447,n15479,n15480);
  or U16354(n15449,n15479,n15480);
  nand U16355(n15480,n15481,n15482,n15483,n15484);
  nand U16356(n15484,n12689,n14590);
  nand U16357(n15483,n14591,n12539);
  nand U16358(n15482,n14814,G36560);
  nand U16359(n15481,n14815,G36592);
  xor U16360(n15479,n15485,n14550);
  nand U16361(n15485,n15486,n15487,n15488);
  nand U16362(n15488,n14590,n12539);
  nand U16363(n15487,n12689,n14596);
  nand U16364(n12689,n15489,n15476);
  nand U16365(n15476,n15490,n14516);
  nand U16366(n15489,n14823,n13689);
  nand U16367(n15486,n13689,n14820);
  and U16368(n13689,n15491,n15492);
  nand U16369(n15492,n15493,n14904);
  or U16370(n15491,n15494,n14904);
  nand U16371(n15450,n15495,n15496);
  nand U16372(n15496,n15497,n14550);
  nand U16373(G7380,n15498,n15499,n15500,n15501);
  nand U16374(n15501,n14514,n14296);
  nand U16375(n14296,n15502,n15503);
  nand U16376(n15503,G36463,n14831);
  not U16377(n14831,n14530);
  nand U16378(n15500,n14545,n12810);
  xor U16379(n12810,n15504,n14592);
  nand U16380(n15504,n15495,n15497);
  nand U16381(n15497,n15505,n15506);
  not U16382(n15506,n15507);
  xor U16383(n15505,n15508,n14592);
  not U16384(n14592,n14550);
  nand U16385(n15495,n15509,n15507);
  nand U16386(n15507,n15510,n15511,n15512,n15513);
  nand U16387(n15513,n14591,n12542);
  or U16388(n14591,n14596,n13324);
  nand U16389(n15512,n12811,n14590);
  nand U16390(n15511,n14814,G36559);
  nand U16391(n15510,n14815,G36591);
  xor U16392(n15509,n14550,n15508);
  nand U16393(n15508,n15514,n15515,n15516);
  nand U16394(n15516,n12811,n14596);
  nand U16395(n14596,n14559,n14557);
  nand U16396(n14557,n15517,n15518);
  nand U16397(n14559,n15518,n14504);
  nand U16398(n15518,n15519,n15520,n15521);
  nand U16399(n15521,n15522,n13899);
  nand U16400(n15520,n15523,n15524);
  not U16401(n15524,n12935);
  or U16402(n15519,n14011,n15525);
  nor U16403(n14011,n13656,n12948);
  not U16404(n12948,n13654);
  nand U16405(n13654,n14284,n12950);
  nand U16406(n12811,n15526,n15502);
  nand U16407(n15502,n15527,n14516);
  nand U16408(n15526,n14823,G36463);
  not U16409(n14823,n14516);
  nand U16410(n15515,n14590,n12542);
  nand U16411(n12542,n15528,n15529,n15530,n15531);
  nand U16412(n15531,G36591,n14527);
  nand U16413(n15530,G36559,n14528);
  nand U16414(n15529,G36527,n14529);
  nand U16415(n15528,G36685,n14583);
  not U16416(n14558,n14567);
  nand U16417(n14567,n15532,n15533);
  nand U16418(n15533,n12971,n14502,n15522);
  nand U16419(n14502,n15534,n14303);
  nand U16420(n15532,n15535,n14504);
  not U16421(n14504,n15517);
  nand U16422(n15535,n15536,n15537);
  nand U16423(n15537,n15523,n14284);
  nand U16424(n15536,n15538,n14283);
  not U16425(n14283,n14012);
  nor U16426(n14012,n12949,n13031);
  not U16427(n14556,n14566);
  nand U16428(n14566,n15539,n15540,n15541,n15542);
  nand U16429(n15542,n15522,n12971,n15534,n14303);
  and U16430(n15522,n15523,n12953);
  nand U16431(n15541,n15517,n15538,n13031);
  nor U16432(n13031,n13899,n12974,n13025);
  nand U16433(n15540,n14284,n15517,n15523);
  nor U16434(n15523,n12950,n15525);
  nand U16435(n15539,n15517,n15538,n12949);
  nor U16436(n12949,n12974,n12971,n13025);
  nand U16437(n15514,G36463,n14820);
  or U16438(n14820,n14815,n14814);
  nor U16439(n14814,n14008,n14017);
  not U16440(n14008,n13660);
  nor U16441(n14815,n14017,n13660);
  nand U16442(n14550,n15543,n15544,n15538);
  nand U16443(n15544,n13025,n13899);
  nand U16444(n15543,n12950,n12974);
  not U16445(n14545,n15139);
  nand U16446(n15139,n14521,n14499);
  nand U16447(n14499,n15545,n12969,n12942);
  not U16448(n12942,n14282);
  nand U16449(n14282,n15546,n13652);
  nand U16450(n13652,n13025,n13899,n13026);
  nand U16451(n15546,n13656,n12946);
  nand U16452(n15545,n12953,n13653);
  nand U16453(n15499,n14579,n12539);
  nand U16454(n12539,n15547,n15548,n15549,n15550);
  nand U16455(n15550,G36592,n14527);
  nand U16456(n15552,G36493,n15553,n14904);
  nand U16457(n15551,n15554,n15555,G36494);
  nand U16458(n15549,G36560,n14528);
  nand U16459(n15557,G36492,n15558,n14904);
  nand U16460(n15556,n15559,n15560,G36494);
  nand U16461(n15548,G36528,n14529);
  nand U16462(n15562,n15553,n15558,n14904);
  not U16463(n15553,G36492);
  nand U16464(n15561,n15560,n15555,G36494);
  not U16465(n15555,n15559);
  nand U16466(n15547,G36695,n14583);
  nand U16467(n14583,n15563,n15564);
  nand U16468(n15564,G36493,G36492,n14904);
  nand U16469(n15563,n15559,n15554,G36494);
  not U16470(n14579,n15466);
  nand U16471(n15466,n14297,n14521);
  and U16472(n14297,n12934,n12918);
  nand U16473(n12918,n14530,n15565);
  not U16474(n15565,n14532);
  nand U16475(n14532,n15566,n15567);
  nand U16476(n15567,n15568,G36494,n15473);
  nand U16477(n15566,n15569,G36491);
  nor U16478(n14530,n15570,n15571);
  nor U16479(n15571,G36491,G36494,G36490);
  and U16480(n15570,n15572,n15474);
  nand U16481(n15498,n14517,G36527);
  not U16482(n14517,n14521);
  nand U16483(n14521,n15573,n15574);
  nand U16484(n15574,n12923,n15575);
  nand U16485(n15575,n15576,n15577);
  nand U16486(n15577,n12917,n14306,n13642,n13029);
  nand U16487(n13642,n14510,n12971);
  not U16488(n14510,n14506);
  nand U16489(n14506,n13026,n12953);
  not U16490(n12953,n12974);
  nand U16491(n14306,n14284,n14295);
  not U16492(n14295,n13653);
  nand U16493(n13653,n13025,n12946);
  not U16494(n14284,n12969);
  nand U16495(n12969,n12971,n12974);
  not U16496(n12917,n12929);
  nand U16497(n12929,n14503,n14303,n15534);
  nand U16498(n15576,n12928,n12937);
  nor U16499(n12928,n12952,n12974);
  nand U16500(n12952,n12971,n13025,n13026);
  not U16501(n12971,n13899);
  nand U16502(n15573,n12915,n12937);
  not U16503(n12937,n12931);
  nand U16504(n12931,n15517,n14503);
  nand U16505(n14503,n15578,n15579);
  nand U16506(n15579,n15580,n15581,n15582,n15583);
  nor U16507(n15583,n15584,n15585,n15586,n15587);
  nand U16508(n15587,n15588,n15589,n15590);
  nand U16509(n15586,n15591,n15592,n15593,n15594);
  nand U16510(n15585,n15595,n15596,n15597,n15598);
  nand U16511(n15584,n15599,n15600,n15601,n15602);
  nor U16512(n15582,n15603,G36497,G36499,G36498);
  nand U16513(n15603,n15604,n15605,n15606,n15607);
  nor U16514(n15581,G36511,G36510,G36509,G36508);
  nor U16515(n15580,G36507,G36506,G36505,G36504);
  nor U16516(n15517,n14303,n15534);
  and U16517(n15534,n15608,n15609);
  nand U16518(n15609,G36495,n15578);
  not U16519(n15578,n15610);
  nand U16520(n15608,n12550,n15610);
  nand U16521(n12550,n15611,n15612);
  nand U16522(n14303,n12547,n15613);
  or U16523(n15613,n15610,G36496);
  nand U16524(n12547,n15612,n15614);
  and U16525(n12915,n13026,n12923,n13656);
  nor U16526(n13656,n12935,n13025);
  nand U16527(n12935,n12974,n13899);
  nand U16528(n13899,n15615,n15616,n15617);
  nand U16529(n15616,n15618,n14904);
  nand U16530(n15615,G36482,n15619,G36494);
  nand U16531(n12974,n15620,n15621,n15622);
  nand U16532(n15621,n15623,n14904);
  nand U16533(n15620,G36483,n15617,G36494);
  nor U16534(G7379,n12546,n15602);
  not U16535(n15602,G36526);
  nor U16536(G7378,n12546,n15601);
  not U16537(n15601,G36525);
  nor U16538(G7377,n12546,n15600);
  not U16539(n15600,G36524);
  nor U16540(G7376,n12546,n15599);
  not U16541(n15599,G36523);
  nor U16542(G7375,n12546,n15598);
  not U16543(n15598,G36522);
  nor U16544(G7374,n12546,n15597);
  not U16545(n15597,G36521);
  nor U16546(G7373,n12546,n15596);
  not U16547(n15596,G36520);
  nor U16548(G7372,n12546,n15595);
  not U16549(n15595,G36519);
  nor U16550(G7371,n12546,n15594);
  not U16551(n15594,G36518);
  nor U16552(G7370,n12546,n15593);
  not U16553(n15593,G36517);
  nor U16554(G7369,n12546,n15592);
  not U16555(n15592,G36516);
  nor U16556(G7368,n12546,n15591);
  not U16557(n15591,G36515);
  nor U16558(G7367,n12546,n15589);
  not U16559(n15589,G36514);
  nor U16560(G7366,n12546,n15588);
  not U16561(n15588,G36513);
  nor U16562(G7365,n12546,n15590);
  not U16563(n15590,G36512);
  and U16564(G7364,n12545,G36511);
  and U16565(G7363,n12545,G36510);
  and U16566(G7362,n12545,G36509);
  and U16567(G7361,n12545,G36508);
  and U16568(G7360,n12545,G36507);
  and U16569(G7359,n12545,G36506);
  and U16570(G7358,n12545,G36505);
  and U16571(G7357,n12545,G36504);
  nor U16572(G7356,n12546,n15607);
  not U16573(n15607,G36503);
  nor U16574(G7355,n12546,n15606);
  not U16575(n15606,G36502);
  nor U16576(G7354,n12546,n15605);
  not U16577(n15605,G36501);
  nor U16578(G7353,n12546,n15604);
  not U16579(n15604,G36500);
  not U16580(n12546,n12545);
  and U16581(G7352,n12545,G36499);
  and U16582(G7351,n12545,G36498);
  and U16583(G7350,n12545,G36497);
  nand U16584(n12545,n12923,n15610);
  nand U16585(n15610,n15624,n15625,n15626);
  not U16586(n15626,n15612);
  nand U16587(n15625,n15627,n14533);
  not U16588(n14533,G36675);
  nand U16589(n15624,n15611,n15614,G36675);
  and U16590(n12923,n15538,G36705);
  nor U16591(n15538,n13324,n15525);
  not U16592(n13324,n13318);
  nand U16593(G7349,n15628,n15629);
  nand U16594(n15629,n15630,n15558,n15631);
  not U16595(n15558,G36493);
  nand U16596(n15628,n14515,G7317);
  nand U16597(n14515,n15632,n15633);
  nand U16598(n15633,n15634,n15635);
  nand U16599(n15635,n15636,n15637);
  nand U16600(n15637,n15638,n15639,n15640);
  xor U16601(n15640,G36429,G36184);
  nand U16602(n15639,G36428,n15641);
  nand U16603(n15636,n15641,n15642,n15643);
  xor U16604(n15643,G36184,n15644);
  nand U16605(n15642,n15638,n15645);
  nand U16606(n15638,n15646,n15647);
  nand U16607(n15641,G36183,n15648);
  not U16608(n15648,n15646);
  nand U16609(n15632,G1,n15649);
  nand U16610(G7348,n15650,n15651,n15652);
  nand U16611(n15652,n15653,G36493);
  nand U16612(n15651,n15631,n15554);
  not U16613(n15554,n15560);
  xor U16614(n15560,n15630,G36493);
  nand U16615(n15650,n14520,G7317);
  nand U16616(n14520,n15654,n15655);
  nand U16617(n15655,n15634,n15656);
  xor U16618(n15656,n15646,n15657);
  xor U16619(n15657,G36428,G36183);
  nand U16620(n15646,n15658,n15659);
  nand U16621(n15659,G36427,n15660);
  or U16622(n15660,n15661,n15662);
  nand U16623(n15658,n15662,n15661);
  nand U16624(n15654,n15649,G2);
  nand U16625(G7347,n15663,n15664,n15665);
  nand U16626(n15665,n15653,G36492);
  nand U16627(n15664,n15631,n15559);
  nor U16628(n15559,n15630,n15666);
  and U16629(n15666,G36492,n15667);
  nor U16630(n15630,n15667,G36492);
  nand U16631(n15663,n14572,G7317);
  nand U16632(n14572,n15668,n15669);
  nand U16633(n15669,n15634,n15670);
  xor U16634(n15670,n15662,n15671);
  xor U16635(n15671,G36427,G36182);
  nand U16636(n15662,n15672,n15673);
  nand U16637(n15673,G36426,n15674);
  or U16638(n15674,n15675,n15676);
  nand U16639(n15672,n15675,n15676);
  nand U16640(n15668,n15649,G3);
  nand U16641(G7346,n15677,n15678,n15679);
  nand U16642(n15679,n15653,G36491);
  nand U16643(n15678,n14597,G7317);
  nand U16644(n14597,n15680,n15681);
  nand U16645(n15681,n15634,n15682);
  xor U16646(n15682,n15675,n15683);
  xor U16647(n15683,G36426,G36181);
  nand U16648(n15675,n15684,n15685);
  nand U16649(n15685,G36425,n15686);
  or U16650(n15686,n15687,n15688);
  nand U16651(n15684,n15687,n15688);
  nand U16652(n15680,n15649,G4);
  nand U16653(n15677,n15631,n15473);
  nand U16654(G7345,n15689,n15690,n15691);
  nand U16655(n15691,n15653,G36490);
  nand U16656(n15690,n14620,G7317);
  nand U16657(n14620,n15692,n15693);
  nand U16658(n15693,n15634,n15694);
  xor U16659(n15694,n15687,n15695);
  xor U16660(n15695,G36425,G36180);
  nand U16661(n15687,n15696,n15697);
  nand U16662(n15697,G36424,n15698);
  or U16663(n15698,n15699,n15700);
  nand U16664(n15696,n15700,n15699);
  nand U16665(n15692,n15649,G5);
  nand U16666(n15689,n15631,n15568);
  not U16667(n15568,n15474);
  nand U16668(G7344,n15701,n15702,n15703);
  nand U16669(n15703,n15653,G36489);
  nand U16670(n15702,n15704,n15705,n15631);
  nand U16671(n15701,n14646,G7317);
  nand U16672(n14646,n15706,n15707);
  nand U16673(n15707,n15634,n15708);
  xor U16674(n15708,n15700,n15709);
  xor U16675(n15709,G36424,G36179);
  nand U16676(n15700,n15710,n15711);
  nand U16677(n15711,G36423,n15712);
  or U16678(n15712,n15713,n15714);
  nand U16679(n15710,n15714,n15713);
  nand U16680(n15706,G6,n15649);
  nand U16681(G7343,n15715,n15716,n15717);
  nand U16682(n15717,n14671,G7317);
  nand U16683(n14671,n15718,n15719);
  nand U16684(n15719,n15634,n15720);
  xor U16685(n15720,n15714,n15721);
  xor U16686(n15721,G36423,G36178);
  nand U16687(n15714,n15722,n15723);
  nand U16688(n15723,G36422,n15724);
  or U16689(n15724,n15725,n15726);
  nand U16690(n15722,n15726,n15725);
  nand U16691(n15718,G7,n15649);
  nand U16692(n15716,G36488,n15727);
  nand U16693(n15727,n15728,n15729);
  nand U16694(n15729,n15631,n15730);
  nand U16695(n15715,n15631,n15731,n15732);
  nand U16696(G7342,n15733,n15734,n15735);
  nand U16697(n15735,n15653,G36487);
  nand U16698(n15734,n15736,n15731,n15631);
  nand U16699(n15733,n14696,G7317);
  nand U16700(n14696,n15737,n15738);
  nand U16701(n15738,n15634,n15739);
  xor U16702(n15739,n15726,n15740);
  xor U16703(n15740,G36422,G36177);
  nand U16704(n15726,n15741,n15742);
  nand U16705(n15742,G36421,n15743);
  or U16706(n15743,n15744,n15745);
  nand U16707(n15741,n15745,n15744);
  nand U16708(n15737,G8,n15649);
  nand U16709(G7341,n15746,n15747,n15748);
  nand U16710(n15748,n14721,G7317);
  nand U16711(n14721,n15749,n15750);
  nand U16712(n15750,n15634,n15751);
  xor U16713(n15751,n15745,n15752);
  xor U16714(n15752,G36421,G36176);
  nand U16715(n15745,n15753,n15754);
  nand U16716(n15754,G36420,n15755);
  or U16717(n15755,n15756,n15757);
  nand U16718(n15753,n15757,n15756);
  nand U16719(n15749,G9,n15649);
  nand U16720(n15747,G36486,n15758);
  nand U16721(n15758,n15728,n15759);
  nand U16722(n15759,n15631,n15760);
  nand U16723(n15746,n15631,n15761,n15762);
  nand U16724(G7340,n15763,n15764,n15765);
  nand U16725(n15765,n15653,G36485);
  nand U16726(n15764,n15766,n15761,n15631);
  nand U16727(n15763,n14746,G7317);
  nand U16728(n14746,n15767,n15768);
  nand U16729(n15768,n15634,n15769);
  xor U16730(n15769,n15757,n15770);
  xor U16731(n15770,G36420,G36175);
  nand U16732(n15757,n15771,n15772);
  nand U16733(n15772,G36419,n15773);
  or U16734(n15773,n15774,n15775);
  nand U16735(n15771,n15775,n15774);
  nand U16736(n15767,G10,n15649);
  nand U16737(G7339,n15776,n15777,n15778);
  nand U16738(n15778,n15653,G36484);
  nand U16739(n15777,n15779,n15780,n15631);
  nand U16740(n15776,n14771,G7317);
  nand U16741(n14771,n15781,n15782);
  nand U16742(n15782,n15634,n15783);
  xor U16743(n15783,n15775,n15784);
  xor U16744(n15784,G36419,G36174);
  nand U16745(n15775,n15785,n15786);
  nand U16746(n15786,G36418,n15787);
  or U16747(n15787,n15788,n15789);
  nand U16748(n15785,n15789,n15788);
  nand U16749(n15781,G11,n15649);
  nand U16750(G7338,n15790,n15791,n15792);
  nand U16751(n15792,n14796,G7317);
  nand U16752(n14796,n15793,n15794);
  nand U16753(n15794,n15634,n15795);
  xor U16754(n15795,n15789,n15796);
  xor U16755(n15796,G36418,G36173);
  nand U16756(n15789,n15797,n15798);
  nand U16757(n15798,G36417,n15799);
  or U16758(n15799,n15800,n15801);
  nand U16759(n15797,n15801,n15800);
  nand U16760(n15793,G12,n15649);
  nand U16761(n15791,G36483,n15802);
  nand U16762(n15802,n15728,n15803);
  nand U16763(n15803,n15631,n15804);
  nand U16764(n15790,n15631,n15617,n15623);
  nand U16765(G7337,n15805,n15806,n15807);
  nand U16766(n15807,n14824,G7317);
  nand U16767(n14824,n15808,n15809);
  nand U16768(n15809,n15634,n15810);
  xor U16769(n15810,n15801,n15811);
  xor U16770(n15811,G36417,G36172);
  nand U16771(n15801,n15812,n15813);
  nand U16772(n15813,G36416,n15814);
  or U16773(n15814,n15815,n15816);
  nand U16774(n15812,n15816,n15815);
  nand U16775(n15808,G13,n15649);
  nand U16776(n15806,G36482,n15817);
  nand U16777(n15817,n15728,n15818);
  nand U16778(n15818,n15631,n15819);
  nand U16779(n15805,n15631,n15619,n15618);
  nand U16780(G7336,n15820,n15821,n15822);
  nand U16781(n15822,n15653,G36481);
  or U16782(n15821,n14866,n15823);
  nand U16783(n14866,n15619,n15824);
  nand U16784(n15824,G36481,n14902);
  not U16785(n15619,n15819);
  nand U16786(n15820,n14857,G7317);
  nand U16787(n14857,n15825,n15826);
  nand U16788(n15826,n15634,n15827);
  xor U16789(n15827,n15816,n15828);
  xor U16790(n15828,G36416,G36171);
  nand U16791(n15816,n15829,n15830);
  nand U16792(n15830,G36415,n15831);
  or U16793(n15831,n15832,n15833);
  nand U16794(n15829,n15833,n15832);
  nand U16795(n15825,G14,n15649);
  nand U16796(G7335,n15834,n15835,n15836);
  nand U16797(n15836,n14893,G7317);
  nand U16798(n14893,n15837,n15838);
  nand U16799(n15838,n15634,n15839);
  xor U16800(n15839,n15833,n15840);
  xor U16801(n15840,G36415,G36170);
  nand U16802(n15833,n15841,n15842);
  nand U16803(n15842,G36414,n15843);
  nand U16804(n15843,G36169,n15844);
  or U16805(n15841,n15844,G36169);
  nand U16806(n15837,G15,n15649);
  nand U16807(n15835,G36480,n15845);
  nand U16808(n15845,n15728,n15846);
  nand U16809(n15846,n15631,n15847);
  nand U16810(n15834,n15631,n14905,n14903);
  nand U16811(G7334,n15848,n15849,n15850);
  nand U16812(n15850,n15653,G36479);
  or U16813(n15849,n14939,n15823);
  nand U16814(n14939,n14905,n15851);
  nand U16815(n15851,G36479,n14974);
  not U16816(n14905,n15847);
  nand U16817(n15848,n14930,G7317);
  nand U16818(n14930,n15852,n15853);
  nand U16819(n15853,n15634,n15854);
  xnor U16820(n15854,n15844,n15855);
  xor U16821(n15855,G36414,G36169);
  and U16822(n15844,n15856,n15857);
  nand U16823(n15857,G36413,n15858);
  nand U16824(n15858,G36168,n15859);
  or U16825(n15856,n15859,G36168);
  nand U16826(n15852,G16,n15649);
  nand U16827(G7333,n15860,n15861,n15862);
  nand U16828(n15862,n14965,G7317);
  nand U16829(n14965,n15863,n15864);
  nand U16830(n15864,n15634,n15865);
  xnor U16831(n15865,n15859,n15866);
  xor U16832(n15866,G36413,G36168);
  and U16833(n15859,n15867,n15868);
  nand U16834(n15868,G36412,n15869);
  nand U16835(n15869,G36167,n15870);
  or U16836(n15867,n15870,G36167);
  nand U16837(n15863,n15649,G17);
  nand U16838(n15861,G36478,n15871);
  nand U16839(n15871,n15728,n15872);
  nand U16840(n15872,n15631,n15873);
  nand U16841(n15860,n15631,n14976,n14975);
  nand U16842(G7332,n15874,n15875,n15876);
  nand U16843(n15876,n15653,G36477);
  or U16844(n15875,n15011,n15823);
  nand U16845(n15011,n14976,n15877);
  nand U16846(n15877,G36477,n15048);
  not U16847(n14976,n15873);
  nand U16848(n15874,n15012,G7317);
  not U16849(n15012,n15002);
  nor U16850(n15002,n15878,n15879);
  and U16851(n15878,n15880,n15634);
  xnor U16852(n15880,n15870,n15881);
  xor U16853(n15881,G36412,G36167);
  and U16854(n15870,n15882,n15883);
  nand U16855(n15883,G36411,n15884);
  or U16856(n15884,n15885,n15886);
  nand U16857(n15882,n15886,n15885);
  nand U16858(G7331,n15887,n15888,n15889);
  nand U16859(n15889,n15039,G7317);
  nand U16860(n15039,n15890,n15891);
  nand U16861(n15891,n15634,n15892);
  xor U16862(n15892,n15886,n15893);
  xor U16863(n15893,G36411,G36166);
  nand U16864(n15886,n15894,n15895);
  nand U16865(n15895,G36410,n15896);
  nand U16866(n15896,G36165,n15897);
  or U16867(n15894,n15897,G36165);
  nand U16868(n15890,G19,n15649);
  nand U16869(n15888,G36476,n15898);
  nand U16870(n15898,n15728,n15899);
  nand U16871(n15899,n15631,n15900);
  nand U16872(n15887,n15631,n15050,n15049);
  nand U16873(G7330,n15901,n15902,n15903);
  nand U16874(n15903,n15653,G36475);
  or U16875(n15902,n15084,n15823);
  nand U16876(n15084,n15050,n15904);
  nand U16877(n15904,G36475,n15117);
  not U16878(n15050,n15900);
  nand U16879(n15901,n15075,G7317);
  nand U16880(n15075,n15905,n15906);
  nand U16881(n15906,n15634,n15907);
  xnor U16882(n15907,n15897,n15908);
  xor U16883(n15908,G36410,G36165);
  and U16884(n15897,n15909,n15910);
  nand U16885(n15910,G36409,n15911);
  nand U16886(n15911,G36164,n15912);
  or U16887(n15909,n15912,G36164);
  nand U16888(n15905,G20,n15649);
  nand U16889(G7329,n15913,n15914,n15915);
  nand U16890(n15915,n15112,G7317);
  nand U16891(n15112,n15916,n15917);
  nand U16892(n15917,n15634,n15918);
  xnor U16893(n15918,n15912,n15919);
  xor U16894(n15919,G36409,G36164);
  and U16895(n15912,n15920,n15921);
  nand U16896(n15921,G36408,n15922);
  nand U16897(n15922,G36163,n15923);
  or U16898(n15920,n15923,G36163);
  nand U16899(n15916,n15649,G21);
  nand U16900(n15914,G36474,n15924);
  nand U16901(n15924,n15728,n15925);
  nand U16902(n15925,n15631,n15926);
  nand U16903(n15913,n15631,n15119,n15118);
  nand U16904(G7328,n15927,n15928,n15929);
  nand U16905(n15929,n15653,G36473);
  or U16906(n15928,n15170,n15823);
  nand U16907(n15170,n15119,n15930);
  nand U16908(n15930,G36473,n15201);
  not U16909(n15119,n15926);
  nand U16910(n15927,n15171,G7317);
  not U16911(n15171,n15165);
  nor U16912(n15165,n15931,n15932);
  and U16913(n15931,n15933,n15634);
  xnor U16914(n15933,n15923,n15934);
  xor U16915(n15934,G36408,G36163);
  and U16916(n15923,n15935,n15936);
  nand U16917(n15936,G36407,n15937);
  or U16918(n15937,n15938,n15939);
  nand U16919(n15935,n15939,n15938);
  nand U16920(G7327,n15940,n15941,n15942);
  nand U16921(n15942,n15192,G7317);
  nand U16922(n15192,n15943,n15944);
  nand U16923(n15944,n15634,n15945);
  xor U16924(n15945,n15939,n15946);
  xor U16925(n15946,G36407,G36162);
  nand U16926(n15939,n15947,n15948);
  nand U16927(n15948,G36406,n15949);
  or U16928(n15949,n15950,n15951);
  nand U16929(n15947,n15951,n15950);
  nand U16930(n15943,G23,n15649);
  nand U16931(n15941,G36472,n15952);
  nand U16932(n15952,n15728,n15953);
  nand U16933(n15953,n15631,n15954);
  nand U16934(n15940,n15631,n15203,n15202);
  nand U16935(G7326,n15955,n15956,n15957);
  nand U16936(n15957,n15653,G36471);
  or U16937(n15956,n15236,n15823);
  nand U16938(n15236,n15203,n15958);
  nand U16939(n15958,G36471,n15273);
  not U16940(n15203,n15954);
  nand U16941(n15955,n15227,G7317);
  nand U16942(n15227,n15959,n15960);
  nand U16943(n15960,n15634,n15961);
  xor U16944(n15961,n15951,n15962);
  xor U16945(n15962,G36406,G36161);
  nand U16946(n15951,n15963,n15964);
  nand U16947(n15964,G36405,n15965);
  nand U16948(n15965,n15966,G36160);
  or U16949(n15963,n15966,G36160);
  nand U16950(n15959,G24,n15649);
  nand U16951(G7325,n15967,n15968,n15969);
  nand U16952(n15969,n15264,G7317);
  nand U16953(n15264,n15970,n15971);
  nand U16954(n15971,n15634,n15972);
  xnor U16955(n15972,n15966,n15973);
  xor U16956(n15973,G36405,G36160);
  and U16957(n15966,n15974,n15975);
  nand U16958(n15975,G36404,n15976);
  nand U16959(n15976,G36159,n15977);
  or U16960(n15974,n15977,G36159);
  nand U16961(n15970,G25,n15649);
  nand U16962(n15968,G36470,n15978);
  nand U16963(n15978,n15728,n15979);
  nand U16964(n15979,n15631,n15980);
  nand U16965(n15967,n15631,n15275,n15274);
  nand U16966(G7324,n15981,n15982,n15983);
  nand U16967(n15983,n15653,G36469);
  or U16968(n15982,n15309,n15823);
  nand U16969(n15309,n15275,n15984);
  nand U16970(n15984,G36469,n15345);
  not U16971(n15275,n15980);
  nand U16972(n15981,n15310,G7317);
  not U16973(n15310,n15300);
  nor U16974(n15300,n15985,n15986);
  and U16975(n15985,n15987,n15634);
  xnor U16976(n15987,n15977,n15988);
  xor U16977(n15988,G36404,G36159);
  and U16978(n15977,n15989,n15990);
  nand U16979(n15990,G36403,n15991);
  nand U16980(n15991,G36158,n15992);
  or U16981(n15989,n15992,G36158);
  nand U16982(G7323,n15993,n15994,n15995);
  nand U16983(n15995,n15348,G7317);
  not U16984(n15348,n15336);
  nor U16985(n15336,n15996,n15997);
  and U16986(n15996,n15998,n15634);
  xnor U16987(n15998,n15992,n15999);
  xor U16988(n15999,G36403,G36158);
  and U16989(n15992,n16000,n16001);
  nand U16990(n16001,G36402,n16002);
  nand U16991(n16002,G36157,n16003);
  or U16992(n16000,n16003,G36157);
  nand U16993(n15994,G36468,n16004);
  nand U16994(n16004,n15728,n16005);
  nand U16995(n16005,n15631,n16006);
  nand U16996(n15993,n15631,n15347,n15346);
  nand U16997(G7322,n16007,n16008,n16009);
  nand U16998(n16009,n15653,G36467);
  or U16999(n16008,n15383,n15823);
  nand U17000(n15383,n15347,n16010);
  nand U17001(n16010,G36467,n15419);
  not U17002(n15347,n16006);
  nand U17003(n16007,n15384,G7317);
  not U17004(n15384,n15374);
  nor U17005(n15374,n16011,n16012);
  and U17006(n16011,n16013,n15634);
  xnor U17007(n16013,n16003,n16014);
  xor U17008(n16014,G36402,G36157);
  and U17009(n16003,n16015,n16016);
  nand U17010(n16016,G36401,n16017);
  or U17011(n16017,n16018,n16019);
  nand U17012(n16015,n16019,n16018);
  nand U17013(G7321,n16020,n16021,n16022);
  nand U17014(n16022,n15410,G7317);
  nand U17015(n15410,n16023,n16024);
  nand U17016(n16024,n15634,n16025);
  xor U17017(n16025,n16019,n16026);
  xor U17018(n16026,G36401,G36156);
  nand U17019(n16019,n16027,n16028);
  or U17020(n16027,n16029,n16030);
  nand U17021(n16023,G29,n15649);
  nand U17022(n16021,G36466,n16031);
  nand U17023(n16031,n15728,n16032);
  nand U17024(n16032,n15631,n16033);
  nand U17025(n16020,n15631,n15421,n15420);
  nand U17026(G7320,n16034,n16035,n16036);
  nand U17027(n16036,n15653,G36465);
  or U17028(n16035,n15455,n15823);
  nand U17029(n15455,n15421,n16037);
  nand U17030(n16037,G36465,n16038);
  nand U17031(n16038,n15493,n13671);
  not U17032(n15421,n16033);
  nand U17033(n16034,n15446,G7317);
  nand U17034(n15446,n16039,n16040);
  nand U17035(n16040,n15634,n16041);
  xor U17036(n16041,n16029,n16042);
  nor U17037(n16042,n16030,n16043);
  not U17038(n16043,n16028);
  nand U17039(n16028,G36400,n16044);
  nor U17040(n16030,n16044,G36400);
  not U17041(n16044,G36155);
  nand U17042(n16029,n16045,n16046);
  nand U17043(n16046,n16047,n16048);
  nand U17044(n16047,n16049,n16050);
  nand U17045(n16045,G36154,n16051);
  nand U17046(n16039,G30,n15649);
  nand U17047(G7319,n16052,n16053,n16054);
  nand U17048(n16054,n15653,G36464);
  not U17049(n15653,n15728);
  nand U17050(n16053,n15631,n15494);
  xor U17051(n15494,n15493,n13671);
  not U17052(n13671,G36463);
  not U17053(n15493,G36464);
  nand U17054(n16052,n15490,G7317);
  nand U17055(n15490,n16055,n16056);
  nand U17056(n16056,n15649,G31);
  nand U17057(n16055,n16057,n15634);
  xor U17058(n16057,n16049,n16058);
  xor U17059(n16058,G36399,G36154);
  nand U17060(G7318,n16059,n16060);
  nand U17061(n16060,G36463,n16061);
  nand U17062(n16061,n15728,n15823);
  nand U17063(n15823,n15728,G36705);
  nand U17064(n15728,G36705,n14904);
  nand U17065(n16059,n15527,G7317);
  nand U17066(n15527,n16062,n16063);
  nand U17067(n16063,n15634,n16064);
  nand U17068(n16064,n16051,n16065);
  nand U17069(n16065,G36153,n16066);
  not U17070(n16051,n16049);
  nor U17071(n16049,n16066,G36153);
  nand U17072(n16062,n15649,G32);
  not U17073(G7316,n14018);
  nand U17074(n14018,n16067,n12448);
  nand U17075(n14017,n15525,n13318);
  nor U17076(n15525,n15612,n15611,n15614);
  nand U17077(n15614,n16068,n16069,n16070);
  nand U17078(n16069,n15732,n14904);
  nand U17079(n16068,G36488,n15731,G36494);
  not U17080(n15611,n15627);
  nand U17081(n15627,n16071,n16072);
  nand U17082(n16072,G36487,n14904);
  nand U17083(n16071,n15736,n15731,G36494);
  not U17084(n15731,n15730);
  nand U17085(n15736,G36487,n16073);
  nand U17086(n16073,n15760,n15762);
  not U17087(n15762,G36486);
  nand U17088(n15612,n16074,n16075);
  or U17089(n16075,G36489,G36494);
  nand U17090(n16074,G36494,n16076);
  nand U17091(n16076,n15705,n15704);
  nand U17092(n15704,G36489,n16070);
  nand U17093(n16067,n16077,G36705);
  nand U17094(n16077,n16078,n14516);
  nor U17095(n13661,n15572,n16079);
  nor U17096(n16079,G36491,G36494);
  nor U17097(n15572,n14904,n15473);
  and U17098(n15473,n15667,n16080);
  nand U17099(n16080,G36491,n16081);
  or U17100(n15667,n16081,G36491);
  nor U17101(n13660,n16082,n15569);
  nor U17102(n15569,n15475,G36494);
  not U17103(n15475,G36490);
  nor U17104(n16082,n15474,n14904);
  not U17105(n14904,G36494);
  nand U17106(n15474,n16081,n16083);
  nand U17107(n16083,G36490,n15705);
  or U17108(n16081,n15705,G36490);
  or U17109(n15705,n16070,G36489);
  nand U17110(n16070,n15730,n15732);
  not U17111(n15732,G36488);
  nor U17112(n15730,G36486,G36487,n15761);
  nand U17113(n16078,n12934,n13318);
  xor U17114(n13318,n16084,G36486);
  nand U17115(n16084,G36494,n15761);
  not U17116(n12934,n13029);
  nand U17117(n13029,n12950,n13026);
  not U17118(n13026,n12946);
  nand U17119(n12946,n16085,n16086);
  or U17120(n16086,G36485,G36494);
  nand U17121(n16085,G36494,n16087);
  nand U17122(n16087,n15761,n15766);
  nand U17123(n15766,G36485,n15780);
  not U17124(n15761,n15760);
  nor U17125(n15760,n15780,G36485);
  not U17126(n12950,n13025);
  nand U17127(n13025,n16088,n16089);
  or U17128(n16089,G36484,G36494);
  nand U17129(n16088,G36494,n16090);
  nand U17130(n16090,n15780,n15779);
  nand U17131(n15779,G36484,n15622);
  or U17132(n15780,n15622,G36484);
  nand U17133(n15622,n15804,n15623);
  not U17134(n15623,G36483);
  not U17135(n15804,n15617);
  nand U17136(n15617,n15819,n15618);
  not U17137(n15618,G36482);
  nor U17138(n15819,n14902,G36481);
  nand U17139(n14902,n15847,n14903);
  not U17140(n14903,G36480);
  nor U17141(n15847,n14974,G36479);
  nand U17142(n14974,n15873,n14975);
  not U17143(n14975,G36478);
  nor U17144(n15873,n15048,G36477);
  nand U17145(n15048,n15900,n15049);
  not U17146(n15049,G36476);
  nor U17147(n15900,n15117,G36475);
  nand U17148(n15117,n15926,n15118);
  not U17149(n15118,G36474);
  nor U17150(n15926,n15201,G36473);
  nand U17151(n15201,n15954,n15202);
  not U17152(n15202,G36472);
  nor U17153(n15954,n15273,G36471);
  nand U17154(n15273,n15980,n15274);
  not U17155(n15274,G36470);
  nor U17156(n15980,n15345,G36469);
  nand U17157(n15345,n16006,n15346);
  not U17158(n15346,G36468);
  nor U17159(n16006,n15419,G36467);
  nand U17160(n15419,n16033,n15420);
  not U17161(n15420,G36466);
  nor U17162(n16033,G36464,G36465,G36463);
  nand U17163(G4836,n16091,n16092);
  nand U17164(n16092,G36429,n16093);
  nand U17165(n16091,G4591,n16094);
  nand U17166(G4835,n16095,n16096);
  nand U17167(n16096,G36428,n16093);
  nand U17168(n16095,G4591,n16097);
  nand U17169(G4834,n16098,n16099);
  nand U17170(n16099,G36427,n16093);
  nand U17171(n16098,G4591,n16100);
  nand U17172(G4833,n16101,n16102);
  nand U17173(n16102,G36426,n16093);
  nand U17174(n16101,G4591,n16103);
  nand U17175(G4832,n16104,n16105);
  nand U17176(n16105,G36425,n16093);
  nand U17177(n16104,G4591,n16106);
  nand U17178(G4831,n16107,n16108);
  nand U17179(n16108,G36424,n16093);
  nand U17180(n16107,G4591,n16109);
  nand U17181(G4830,n16110,n16111);
  nand U17182(n16111,G36423,n16093);
  nand U17183(n16110,G4591,n16112);
  nand U17184(G4829,n16113,n16114);
  nand U17185(n16114,G36422,n16093);
  nand U17186(n16113,G4591,n16115);
  nand U17187(G4828,n16116,n16117);
  nand U17188(n16117,G36421,n16093);
  nand U17189(n16116,G4591,n16118);
  nand U17190(G4827,n16119,n16120);
  nand U17191(n16120,G36420,n16093);
  nand U17192(n16119,G4591,n16121);
  nand U17193(G4826,n16122,n16123);
  nand U17194(n16123,G36419,n16093);
  nand U17195(n16122,G4591,n16124);
  nand U17196(G4825,n16125,n16126);
  nand U17197(n16126,G36418,n16093);
  nand U17198(n16125,G4591,n16127);
  nand U17199(G4824,n16128,n16129);
  nand U17200(n16129,G36417,n16093);
  nand U17201(n16128,G4591,n16130);
  nand U17202(G4823,n16131,n16132);
  nand U17203(n16132,G36416,n16093);
  nand U17204(n16131,G4591,n16133);
  nand U17205(G4822,n16134,n16135);
  nand U17206(n16135,G36415,n16093);
  nand U17207(n16134,G4591,n16136);
  nand U17208(G4821,n16137,n16138);
  nand U17209(n16138,G36414,n16093);
  nand U17210(n16137,G4591,n16139);
  nand U17211(G4820,n16140,n16141);
  nand U17212(n16141,G36413,n16093);
  nand U17213(n16140,G4591,n16142);
  nand U17214(G4819,n16143,n16144);
  nand U17215(n16144,G36412,n16093);
  nand U17216(n16143,G4591,n16145);
  nand U17217(G4818,n16146,n16147);
  nand U17218(n16147,G36411,n16093);
  nand U17219(n16146,G4591,n16148);
  nand U17220(G4817,n16149,n16150);
  nand U17221(n16150,G36410,n16093);
  nand U17222(n16149,G4591,n16151);
  nand U17223(G4816,n16152,n16153);
  nand U17224(n16153,G36409,n16093);
  nand U17225(n16152,G4591,n16154);
  nand U17226(G4815,n16155,n16156);
  nand U17227(n16156,G36408,n16093);
  nand U17228(n16155,G4591,n16157);
  nand U17229(G4814,n16158,n16159);
  nand U17230(n16159,G36407,n16093);
  nand U17231(n16158,G4591,n16160);
  nand U17232(G4813,n16161,n16162);
  nand U17233(n16162,G36406,n16093);
  nand U17234(n16161,G4591,n16163);
  nand U17235(G4812,n16164,n16165);
  nand U17236(n16165,G36405,n16093);
  nand U17237(n16164,G4591,n16166);
  nand U17238(G4811,n16167,n16168);
  nand U17239(n16168,G36404,n16093);
  nand U17240(n16167,G4591,n16169);
  nand U17241(G4810,n16170,n16171);
  nand U17242(n16171,G36403,n16093);
  nand U17243(n16170,G4591,n16172);
  nand U17244(G4809,n16173,n16174);
  nand U17245(n16174,G36402,n16093);
  nand U17246(n16173,G4591,n16175);
  nand U17247(G4808,n16176,n16177);
  nand U17248(n16177,G36401,n16093);
  nand U17249(n16176,G4591,n16178);
  nand U17250(G4807,n16179,n16180);
  nand U17251(n16180,G36400,n16093);
  nand U17252(n16179,G4591,n16181);
  nand U17253(G4806,n16182,n16183);
  nand U17254(n16183,G36399,n16093);
  nand U17255(n16182,G4591,n16184);
  nand U17256(G4805,n16185,n16186);
  nand U17257(n16186,G36398,n16093);
  nand U17258(n16185,G4591,n16187);
  nand U17259(G4804,n16188,n16189);
  nand U17260(n16189,n16190,n16191);
  nand U17261(n16188,G36345,n16192);
  nand U17262(G4803,n16193,n16194);
  nand U17263(n16194,G36344,n16192);
  nand U17264(n16193,n16190,n16195);
  nand U17265(G4802,n16196,n16197);
  nand U17266(n16197,G36343,n16192);
  nand U17267(n16196,n16190,n16198);
  nand U17268(G4801,n16199,n16200);
  nand U17269(n16200,G36342,n16192);
  nand U17270(n16199,n16190,n16201);
  nand U17271(G4800,n16202,n16203);
  nand U17272(n16203,G36341,n16192);
  nand U17273(n16202,n16190,n16204);
  nand U17274(G4799,n16205,n16206);
  nand U17275(n16206,G36340,n16192);
  nand U17276(n16205,n16190,n16207);
  nand U17277(G4798,n16208,n16209);
  nand U17278(n16209,G36339,n16192);
  nand U17279(n16208,n16190,n16210);
  nand U17280(G4797,n16211,n16212);
  nand U17281(n16212,G36338,n16192);
  nand U17282(n16211,n16190,n16213);
  nand U17283(G4796,n16214,n16215);
  nand U17284(n16215,G36337,n16192);
  nand U17285(n16214,n16190,n16216);
  nand U17286(G4795,n16217,n16218);
  nand U17287(n16218,G36336,n16192);
  nand U17288(n16217,n16190,n16219);
  nand U17289(G4794,n16220,n16221);
  nand U17290(n16221,G36335,n16192);
  nand U17291(n16220,n16190,n16222);
  nand U17292(G4793,n16223,n16224);
  nand U17293(n16224,G36334,n16192);
  nand U17294(n16223,n16190,n16225);
  nand U17295(G4792,n16226,n16227);
  nand U17296(n16227,G36333,n16192);
  nand U17297(n16226,n16190,n16228);
  nand U17298(G4791,n16229,n16230);
  nand U17299(n16230,G36332,n16192);
  nand U17300(n16229,n16190,n16231);
  nand U17301(G4790,n16232,n16233);
  nand U17302(n16233,G36331,n16192);
  nand U17303(n16232,n16190,n16234);
  nand U17304(G4789,n16235,n16236);
  nand U17305(n16236,G36330,n16192);
  nand U17306(n16235,n16190,n16237);
  nand U17307(G4788,n16238,n16239);
  nand U17308(n16239,G36329,n16192);
  nand U17309(n16238,n16190,n16240);
  nand U17310(G4787,n16241,n16242);
  nand U17311(n16242,G36328,n16192);
  nand U17312(n16241,n16190,n16243);
  nand U17313(G4786,n16244,n16245);
  nand U17314(n16245,G36327,n16192);
  nand U17315(n16244,n16190,n16246);
  nand U17316(G4785,n16247,n16248);
  nand U17317(n16248,G36326,n16192);
  nand U17318(n16247,n16190,n16249);
  nand U17319(G4784,n16250,n16251);
  nand U17320(n16251,G36325,n16192);
  nand U17321(n16250,n16190,n16252);
  nand U17322(G4783,n16253,n16254);
  nand U17323(n16254,G36324,n16192);
  nand U17324(n16253,n16190,n16255);
  nand U17325(G4782,n16256,n16257);
  nand U17326(n16257,G36323,n16192);
  nand U17327(n16256,n16190,n16258);
  nand U17328(G4781,n16259,n16260);
  nand U17329(n16260,G36322,n16192);
  nand U17330(n16259,n16190,n16261);
  nand U17331(G4780,n16262,n16263);
  nand U17332(n16263,G36321,n16192);
  nand U17333(n16262,n16190,n16264);
  nand U17334(G4779,n16265,n16266);
  nand U17335(n16266,G36320,n16192);
  nand U17336(n16265,n16190,n16267);
  nand U17337(G4778,n16268,n16269);
  nand U17338(n16269,G36319,n16192);
  nand U17339(n16268,n16190,n16270);
  nand U17340(G4777,n16271,n16272);
  nand U17341(n16272,G36318,n16192);
  nand U17342(n16271,n16190,n16273);
  nand U17343(G4776,n16274,n16275);
  nand U17344(n16275,G36317,n16192);
  nand U17345(n16274,n16190,n16276);
  nand U17346(G4775,n16277,n16278);
  nand U17347(n16278,G36316,n16192);
  nand U17348(n16277,n16190,n16279);
  nand U17349(G4774,n16280,n16281);
  nand U17350(n16281,G36315,n16192);
  nand U17351(n16280,n16190,n16282);
  nand U17352(G4773,n16283,n16284);
  nand U17353(n16284,G36314,n16192);
  nand U17354(n16283,n16190,n16285);
  nand U17355(G4772,n16288,n16289);
  nand U17356(n16289,n16290,n16191);
  nand U17357(n16191,n16291,n16292,n16293);
  nand U17358(n16293,n16294,n16295);
  nand U17359(n16291,n16296,n16297);
  nand U17360(n16288,G36313,n16298);
  nand U17361(G4771,n16299,n16300);
  nand U17362(n16300,n16290,n16195);
  nand U17363(n16195,n16301,n16292,n16302);
  nand U17364(n16302,n16303,n16296);
  nand U17365(n16301,n16304,n16294);
  nand U17366(n16299,G36312,n16298);
  nand U17367(G4770,n16305,n16306);
  nand U17368(n16306,n16290,n16198);
  nand U17369(n16198,n16307,n16308,n16309,n16310);
  nand U17370(n16309,n16311,n16294);
  nand U17371(n16308,n16312,n16313);
  nand U17372(n16307,n16314,n16315);
  nand U17373(n16305,G36311,n16298);
  nand U17374(G4769,n16316,n16317);
  nand U17375(n16317,n16290,n16201);
  nand U17376(n16201,n16318,n16319,n16320,n16321);
  nor U17377(n16321,n16322,n16323);
  nor U17378(n16323,n16324,n16325);
  nor U17379(n16322,n16326,n16327);
  nand U17380(n16320,n16328,n16315);
  nand U17381(n16319,n16329,n16294);
  nand U17382(n16318,n16330,n16313);
  nand U17383(n16316,G36310,n16298);
  nand U17384(G4768,n16331,n16332);
  nand U17385(n16332,n16290,n16204);
  nand U17386(n16204,n16333,n16334,n16335,n16336);
  nor U17387(n16336,n16337,n16338);
  nor U17388(n16338,n16339,n16325);
  nor U17389(n16337,n16340,n16327);
  nand U17390(n16335,n16341,n16315);
  nand U17391(n16334,n16342,n16294);
  nand U17392(n16333,n16343,n16313);
  nand U17393(n16331,G36309,n16298);
  nand U17394(G4767,n16344,n16345);
  nand U17395(n16345,n16290,n16207);
  nand U17396(n16207,n16346,n16347,n16348,n16349);
  nor U17397(n16349,n16350,n16351);
  nor U17398(n16351,n16352,n16325);
  nor U17399(n16350,n16324,n16327);
  nand U17400(n16348,n16353,n16315);
  nand U17401(n16347,n16354,n16294);
  nand U17402(n16346,n16355,n16313);
  nand U17403(n16344,G36308,n16298);
  nand U17404(G4766,n16356,n16357);
  nand U17405(n16357,n16290,n16210);
  nand U17406(n16210,n16358,n16359,n16360,n16361);
  nor U17407(n16361,n16362,n16363);
  nor U17408(n16363,n16364,n16325);
  nor U17409(n16362,n16339,n16327);
  nand U17410(n16360,n16365,n16315);
  nand U17411(n16359,n16366,n16294);
  nand U17412(n16358,n16367,n16313);
  nand U17413(n16356,G36307,n16298);
  nand U17414(G4765,n16368,n16369);
  nand U17415(n16369,n16290,n16213);
  nand U17416(n16213,n16370,n16371,n16372,n16373);
  nor U17417(n16373,n16374,n16375);
  nor U17418(n16375,n16376,n16325);
  nor U17419(n16374,n16352,n16327);
  nand U17420(n16372,n16377,n16315);
  nand U17421(n16371,n16378,n16294);
  nand U17422(n16370,n16379,n16313);
  nand U17423(n16368,G36306,n16298);
  nand U17424(G4764,n16380,n16381);
  nand U17425(n16381,n16290,n16216);
  nand U17426(n16216,n16382,n16383,n16384,n16385);
  nor U17427(n16385,n16386,n16387);
  nor U17428(n16387,n16388,n16325);
  nor U17429(n16386,n16364,n16327);
  nand U17430(n16384,n16389,n16315);
  nand U17431(n16383,n16390,n16294);
  nand U17432(n16382,n16391,n16313);
  nand U17433(n16380,G36305,n16298);
  nand U17434(G4763,n16392,n16393);
  nand U17435(n16393,n16290,n16219);
  nand U17436(n16219,n16394,n16395,n16396,n16397);
  nor U17437(n16397,n16398,n16399);
  nor U17438(n16399,n16400,n16325);
  nor U17439(n16398,n16376,n16327);
  nand U17440(n16396,n16401,n16315);
  nand U17441(n16395,n16402,n16294);
  nand U17442(n16394,n16403,n16313);
  nand U17443(n16392,G36304,n16298);
  nand U17444(G4762,n16404,n16405);
  nand U17445(n16405,n16290,n16222);
  nand U17446(n16222,n16406,n16407,n16408,n16409);
  nor U17447(n16409,n16410,n16411);
  nor U17448(n16411,n16412,n16325);
  nor U17449(n16410,n16388,n16327);
  nand U17450(n16408,n16413,n16315);
  nand U17451(n16407,n16414,n16294);
  nand U17452(n16406,n16415,n16313);
  nand U17453(n16404,G36303,n16298);
  nand U17454(G4761,n16416,n16417);
  nand U17455(n16417,n16290,n16225);
  nand U17456(n16225,n16418,n16419,n16420,n16421);
  nor U17457(n16421,n16422,n16423);
  nor U17458(n16423,n16424,n16325);
  nor U17459(n16422,n16400,n16327);
  nand U17460(n16420,n16425,n16315);
  nand U17461(n16419,n16426,n16294);
  nand U17462(n16418,n16427,n16313);
  nand U17463(n16416,G36302,n16298);
  nand U17464(G4760,n16428,n16429);
  nand U17465(n16429,n16290,n16228);
  nand U17466(n16228,n16430,n16431,n16432,n16433);
  nor U17467(n16433,n16434,n16435);
  nor U17468(n16435,n16436,n16325);
  nor U17469(n16434,n16412,n16327);
  nand U17470(n16432,n16437,n16315);
  nand U17471(n16431,n16438,n16294);
  nand U17472(n16430,n16439,n16313);
  nand U17473(n16428,G36301,n16298);
  nand U17474(G4758,n16440,n16441);
  nand U17475(n16441,n16290,n16231);
  nand U17476(n16231,n16442,n16443,n16444,n16445);
  nor U17477(n16445,n16446,n16447);
  nor U17478(n16447,n16448,n16325);
  nor U17479(n16446,n16424,n16327);
  nand U17480(n16444,n16449,n16315);
  nand U17481(n16443,n16450,n16294);
  nand U17482(n16442,n16451,n16313);
  nand U17483(n16440,G36300,n16298);
  nand U17484(G4755,n16452,n16453);
  nand U17485(n16453,n16290,n16234);
  nand U17486(n16234,n16454,n16455,n16456,n16457);
  nor U17487(n16457,n16458,n16459);
  nor U17488(n16459,n16460,n16325);
  nor U17489(n16458,n16436,n16327);
  nand U17490(n16456,n16461,n16315);
  nand U17491(n16455,n16462,n16294);
  nand U17492(n16454,n16463,n16313);
  nand U17493(n16452,G36299,n16298);
  nand U17494(G4752,n16464,n16465);
  nand U17495(n16465,n16290,n16237);
  nand U17496(n16237,n16466,n16467,n16468,n16469);
  nor U17497(n16469,n16470,n16471);
  nor U17498(n16471,n16472,n16325);
  nor U17499(n16470,n16448,n16327);
  nand U17500(n16468,n16473,n16315);
  nand U17501(n16467,n16474,n16294);
  nand U17502(n16466,n16475,n16313);
  nand U17503(n16464,G36298,n16298);
  nand U17504(G4749,n16476,n16477);
  nand U17505(n16477,n16290,n16240);
  nand U17506(n16240,n16478,n16479,n16480,n16481);
  nor U17507(n16481,n16482,n16483);
  nor U17508(n16483,n16484,n16325);
  nor U17509(n16482,n16460,n16327);
  nand U17510(n16480,n16485,n16315);
  nand U17511(n16479,n16486,n16294);
  nand U17512(n16478,n16487,n16313);
  nand U17513(n16476,G36297,n16298);
  nand U17514(G4746,n16488,n16489);
  nand U17515(n16489,n16290,n16243);
  nand U17516(n16243,n16490,n16491,n16492,n16493);
  nor U17517(n16493,n16494,n16495);
  nor U17518(n16495,n16496,n16325);
  nor U17519(n16494,n16472,n16327);
  nand U17520(n16492,n16497,n16315);
  nand U17521(n16491,n16498,n16294);
  nand U17522(n16490,n16499,n16313);
  nand U17523(n16488,G36296,n16298);
  nand U17524(G4743,n16500,n16501);
  nand U17525(n16501,n16290,n16246);
  nand U17526(n16246,n16502,n16503,n16504,n16505);
  nor U17527(n16505,n16506,n16507);
  nor U17528(n16507,n16508,n16325);
  nor U17529(n16506,n16484,n16327);
  nand U17530(n16504,n16509,n16315);
  nand U17531(n16503,n16510,n16294);
  nand U17532(n16502,n16511,n16313);
  nand U17533(n16500,G36295,n16298);
  nand U17534(G4740,n16512,n16513);
  nand U17535(n16513,n16290,n16249);
  nand U17536(n16249,n16514,n16515,n16516,n16517);
  nor U17537(n16517,n16518,n16519);
  nor U17538(n16519,n16520,n16325);
  nor U17539(n16518,n16496,n16327);
  nand U17540(n16516,n16521,n16315);
  nand U17541(n16515,n16522,n16294);
  nand U17542(n16514,n16523,n16313);
  nand U17543(n16512,G36294,n16298);
  nand U17544(G4737,n16524,n16525);
  nand U17545(n16525,n16290,n16252);
  nand U17546(n16252,n16526,n16527,n16528,n16529);
  nor U17547(n16529,n16530,n16531);
  nor U17548(n16531,n16532,n16325);
  nor U17549(n16530,n16508,n16327);
  nand U17550(n16528,n16533,n16315);
  nand U17551(n16527,n16534,n16294);
  nand U17552(n16526,n16535,n16313);
  nand U17553(n16524,G36293,n16298);
  nand U17554(G4734,n16536,n16537);
  nand U17555(n16537,n16290,n16255);
  nand U17556(n16255,n16538,n16539,n16540,n16541);
  nor U17557(n16541,n16542,n16543);
  nor U17558(n16543,n16544,n16325);
  nor U17559(n16542,n16520,n16327);
  nand U17560(n16540,n16545,n16315);
  nand U17561(n16539,n16546,n16294);
  nand U17562(n16538,n16547,n16313);
  nand U17563(n16536,G36292,n16298);
  nand U17564(G4731,n16548,n16549);
  nand U17565(n16549,n16290,n16258);
  nand U17566(n16258,n16550,n16551,n16552,n16553);
  nor U17567(n16553,n16554,n16555);
  nor U17568(n16555,n16556,n16325);
  nor U17569(n16554,n16532,n16327);
  nand U17570(n16552,n16557,n16315);
  nand U17571(n16551,n16558,n16294);
  nand U17572(n16550,n16559,n16313);
  nand U17573(n16548,G36291,n16298);
  nand U17574(G4728,n16560,n16561);
  nand U17575(n16561,n16290,n16261);
  nand U17576(n16261,n16562,n16563,n16564,n16565);
  nor U17577(n16565,n16566,n16567);
  nor U17578(n16567,n16568,n16325);
  nor U17579(n16566,n16544,n16327);
  nand U17580(n16564,n16569,n16315);
  nand U17581(n16563,n16570,n16294);
  nand U17582(n16562,n16571,n16313);
  nand U17583(n16560,G36290,n16298);
  nand U17584(G4725,n16572,n16573);
  nand U17585(n16573,n16290,n16264);
  nand U17586(n16264,n16574,n16575,n16576,n16577);
  nor U17587(n16577,n16578,n16579);
  nor U17588(n16579,n16580,n16325);
  nor U17589(n16578,n16556,n16327);
  nand U17590(n16576,n16581,n16315);
  nand U17591(n16575,n16582,n16294);
  nand U17592(n16574,n16583,n16313);
  nand U17593(n16572,G36289,n16298);
  nand U17594(G4722,n16584,n16585);
  nand U17595(n16585,n16290,n16267);
  nand U17596(n16267,n16586,n16587,n16588,n16589);
  nor U17597(n16589,n16590,n16591);
  nor U17598(n16591,n16592,n16325);
  nor U17599(n16590,n16568,n16327);
  nand U17600(n16588,n16593,n16315);
  nand U17601(n16587,n16594,n16294);
  nand U17602(n16586,n16595,n16313);
  nand U17603(n16584,G36288,n16298);
  nand U17604(G4719,n16596,n16597);
  nand U17605(n16597,n16290,n16270);
  nand U17606(n16270,n16598,n16599,n16600,n16601);
  nor U17607(n16601,n16602,n16603);
  nor U17608(n16603,n16604,n16325);
  nor U17609(n16602,n16580,n16327);
  nand U17610(n16600,n16605,n16315);
  nand U17611(n16599,n16606,n16294);
  nand U17612(n16598,n16607,n16313);
  nand U17613(n16596,G36287,n16298);
  nand U17614(G4716,n16608,n16609);
  nand U17615(n16609,n16290,n16273);
  nand U17616(n16273,n16610,n16611,n16612,n16613);
  nor U17617(n16613,n16614,n16615);
  nor U17618(n16615,n16616,n16325);
  nor U17619(n16614,n16592,n16327);
  nand U17620(n16612,n16617,n16315);
  nand U17621(n16611,n16618,n16294);
  nand U17622(n16610,n16619,n16313);
  nand U17623(n16608,G36286,n16298);
  nand U17624(G4713,n16620,n16621);
  nand U17625(n16621,n16290,n16276);
  nand U17626(n16276,n16622,n16623,n16624,n16625);
  nor U17627(n16625,n16626,n16627);
  nor U17628(n16627,n16628,n16325);
  nor U17629(n16626,n16604,n16327);
  nand U17630(n16624,n16629,n16315);
  nand U17631(n16623,n16630,n16294);
  nand U17632(n16622,n16631,n16313);
  nand U17633(n16620,G36285,n16298);
  nand U17634(G4710,n16632,n16633);
  nand U17635(n16633,n16290,n16279);
  nand U17636(n16279,n16634,n16635,n16636,n16637);
  nor U17637(n16637,n16638,n16639);
  nor U17638(n16639,n16640,n16325);
  nor U17639(n16638,n16616,n16327);
  nand U17640(n16636,n16641,n16315);
  nand U17641(n16635,n16642,n16294);
  nand U17642(n16634,n16643,n16313);
  nand U17643(n16632,G36284,n16298);
  nand U17644(G4707,n16644,n16645);
  nand U17645(n16645,n16290,n16282);
  nand U17646(n16282,n16646,n16647,n16648,n16649);
  nor U17647(n16649,n16650,n16651);
  nor U17648(n16651,n16628,n16327);
  and U17649(n16650,n16187,n16652);
  nand U17650(n16648,n16653,n16315);
  nand U17651(n16647,n16654,n16294);
  nand U17652(n16646,n16655,n16313);
  nand U17653(n16644,G36283,n16298);
  nand U17654(G4704,n16656,n16657);
  nand U17655(n16657,n16290,n16285);
  nand U17656(n16285,n16658,n16659,n16660,n16661);
  nand U17657(n16661,n16662,n16294);
  nand U17658(n16660,n16665,n16313);
  nand U17659(n16313,n16666,n16667,n16668);
  nand U17660(n16659,n16669,n16315);
  nand U17661(n16315,n16670,n16671,n16672);
  nand U17662(n16670,n16673,n16674);
  nand U17663(n16658,n16675,n16184);
  nand U17664(n16656,G36282,n16298);
  and U17665(n16286,n16677,n16678,n16679,n16680);
  nand U17666(n16679,n16296,n16681);
  nand U17667(G4693,n16682,n16683);
  nand U17668(n16683,G36251,n16684);
  nand U17669(n16682,n16685,n16686);
  nand U17670(G4692,n16687,n16688);
  nand U17671(n16688,n16685,n16689);
  nand U17672(n16687,G36250,n16684);
  nand U17673(G4533,n16690,n16691,n16692,n16693);
  nor U17674(n16693,n16694,n16695,n16696,n16697);
  nor U17675(n16697,n16580,n16698);
  nor U17676(n16696,n16556,n16699);
  nor U17677(n16695,n16700,n16701);
  nor U17678(n16694,n16702,n16703);
  nand U17679(n16692,G36459,G4389);
  nand U17680(n16691,n16704,n16581);
  nand U17681(n16690,n16705,n16583);
  nand U17682(G4532,n16706,n16707,n16708,n16709);
  nor U17683(n16709,n16710,n16711,n16712,n16713);
  nor U17684(n16713,n16339,n16698);
  nor U17685(n16712,n16340,n16699);
  nor U17686(n16711,n16700,n16714);
  nor U17687(n16710,n16715,n16703);
  nand U17688(n16708,G36458,G4389);
  nand U17689(n16707,n16704,n16341);
  nand U17690(n16706,n16705,n16343);
  nand U17691(G4531,n16716,n16717,n16718,n16719);
  nor U17692(n16719,n16720,n16721,n16722,n16723);
  nor U17693(n16723,n16496,n16698);
  nor U17694(n16722,n16472,n16699);
  nor U17695(n16721,n16700,n16724);
  nor U17696(n16720,n16725,n16703);
  nand U17697(n16718,G36457,G4389);
  nand U17698(n16717,n16704,n16497);
  nand U17699(n16716,n16705,n16499);
  nand U17700(G4530,n16726,n16727,n16728,n16729);
  nor U17701(n16729,n16730,n16731,n16732,n16733);
  nor U17702(n16733,n16388,n16698);
  nor U17703(n16732,n16364,n16699);
  nor U17704(n16731,n16700,n16734);
  nor U17705(n16730,n16735,n16703);
  nand U17706(n16728,G36456,G4389);
  nand U17707(n16727,n16704,n16389);
  nand U17708(n16726,n16705,n16391);
  nand U17709(G4529,n16736,n16737,n16738,n16739);
  nor U17710(n16739,n16740,n16741,n16742,n16743);
  nor U17711(n16743,n16544,n16698);
  nor U17712(n16742,n16520,n16699);
  nor U17713(n16741,n16700,n16744);
  nor U17714(n16740,n16745,n16703);
  nand U17715(n16738,G36455,G4389);
  nand U17716(n16737,n16704,n16545);
  nand U17717(n16736,n16705,n16547);
  nand U17718(G4528,n16746,n16747,n16748,n16749);
  nor U17719(n16749,n16750,n16751,n16752,n16753);
  nor U17720(n16753,n16754,n16755);
  nor U17721(n16752,n16756,n16757);
  nor U17722(n16751,G36454,n16700);
  nand U17723(n16748,n16758,n16181);
  or U17724(n16747,n16703,n16759);
  or U17725(n16746,n16699,n16604);
  nand U17726(G4527,n16760,n16761,n16762,n16763);
  nor U17727(n16763,n16764,n16765,n16766,n16767);
  nor U17728(n16767,n16436,n16698);
  nor U17729(n16766,n16412,n16699);
  nor U17730(n16765,n16700,n16768);
  nor U17731(n16764,n16769,n16703);
  nand U17732(n16762,G36453,G4389);
  nand U17733(n16761,n16704,n16437);
  nand U17734(n16760,n16705,n16439);
  nand U17735(G4526,n16770,n16771,n16772,n16773);
  nor U17736(n16773,n16774,n16775,n16776,n16777);
  nor U17737(n16777,n16324,n16698);
  nor U17738(n16776,n16326,n16699);
  nor U17739(n16775,n16700,n16778);
  not U17740(n16778,n16779);
  nor U17741(n16774,n16780,n16703);
  nand U17742(n16772,G36452,G4389);
  nand U17743(n16771,n16704,n16328);
  nand U17744(n16770,n16705,n16330);
  nand U17745(G4525,n16781,n16782,n16783,n16784);
  nor U17746(n16784,n16785,n16786,n16787,n16788);
  nor U17747(n16788,n16568,n16698);
  nor U17748(n16787,n16544,n16699);
  nor U17749(n16786,n16700,n16789);
  nor U17750(n16785,n16790,n16703);
  nand U17751(n16783,G36451,G4389);
  nand U17752(n16782,n16704,n16569);
  nand U17753(n16781,n16705,n16571);
  nand U17754(G4524,n16791,n16792,n16793,n16794);
  nor U17755(n16794,n16795,n16796,n16797);
  nor U17756(n16797,n16798,n16703);
  nor U17757(n16796,n16799,n16800);
  nor U17758(n16795,n16628,n16699);
  not U17759(n16628,n16181);
  nand U17760(n16793,n16705,n16655);
  nand U17761(n16792,n16758,n16187);
  nand U17762(n16791,n16704,n16653);
  nand U17763(G4523,n16801,n16802,n16803,n16804);
  nor U17764(n16804,n16805,n16806,n16807,n16808);
  nor U17765(n16808,n16412,n16698);
  nor U17766(n16807,n16388,n16699);
  nor U17767(n16806,n16700,n16809);
  not U17768(n16809,n16810);
  nor U17769(n16805,n16811,n16703);
  nand U17770(n16803,G36449,G4389);
  nand U17771(n16802,n16704,n16413);
  nand U17772(n16801,n16705,n16415);
  nand U17773(G4522,n16812,n16813,n16814,n16815);
  nor U17774(n16815,n16816,n16817,n16818,n16819);
  nor U17775(n16819,n16520,n16698);
  nor U17776(n16818,n16496,n16699);
  nor U17777(n16817,n16700,n16820);
  not U17778(n16820,n16821);
  nor U17779(n16816,n16822,n16703);
  nand U17780(n16814,G36448,G4389);
  nand U17781(n16813,n16704,n16521);
  nand U17782(n16812,n16705,n16523);
  nand U17783(G4521,n16823,n16824,n16825,n16826);
  nor U17784(n16826,n16827,n16828,n16829,n16830);
  nor U17785(n16830,n16364,n16698);
  nor U17786(n16829,n16339,n16699);
  nor U17787(n16828,n16700,n16831);
  not U17788(n16831,n16832);
  nor U17789(n16827,n16833,n16703);
  nand U17790(n16825,G36447,G4389);
  nand U17791(n16824,n16704,n16365);
  nand U17792(n16823,n16705,n16367);
  nand U17793(G4520,n16834,n16835,n16836,n16837);
  nor U17794(n16837,n16838,n16839,n16840,n16841);
  nor U17795(n16841,n16472,n16698);
  nor U17796(n16840,n16448,n16699);
  nor U17797(n16839,n16700,n16842);
  nor U17798(n16838,n16843,n16703);
  nand U17799(n16836,G36446,G4389);
  nand U17800(n16835,n16704,n16473);
  nand U17801(n16834,n16705,n16475);
  nand U17802(G4519,n16844,n16845,n16846,n16847);
  nor U17803(n16847,n16848,n16849,n16850,n16851);
  nor U17804(n16851,n16604,n16698);
  nor U17805(n16850,n16580,n16699);
  nor U17806(n16849,n16700,n16852);
  nor U17807(n16848,n16853,n16703);
  nand U17808(n16846,G36445,G4389);
  nand U17809(n16845,n16704,n16605);
  nand U17810(n16844,n16705,n16607);
  nand U17811(G4518,n16854,n16855,n16856,n16857);
  nor U17812(n16857,n16858,n16859,n16860,n16861);
  nor U17813(n16861,n16460,n16698);
  nor U17814(n16860,n16436,n16699);
  nor U17815(n16859,n16700,n16862);
  not U17816(n16862,n16863);
  nor U17817(n16858,n16864,n16703);
  nand U17818(n16856,G36444,G4389);
  nand U17819(n16855,n16704,n16461);
  nand U17820(n16854,n16705,n16463);
  nand U17821(G4517,n16865,n16866,n16867,n16868);
  nor U17822(n16868,n16869,n16870,n16871,n16872);
  nor U17823(n16872,n16376,n16698);
  nor U17824(n16871,n16352,n16699);
  nor U17825(n16870,n16700,n16873);
  nor U17826(n16869,n16874,n16703);
  nand U17827(n16867,G36443,G4389);
  nand U17828(n16866,n16704,n16377);
  nand U17829(n16865,n16705,n16379);
  nand U17830(G4516,n16875,n16876,n16877,n16878);
  nor U17831(n16878,n16879,n16880,n16881,n16882);
  nor U17832(n16882,n16616,n16698);
  nor U17833(n16881,n16592,n16699);
  nor U17834(n16880,n16883,n16703);
  nor U17835(n16879,n16700,n16884);
  nand U17836(n16877,G36442,G4389);
  nand U17837(n16876,n16704,n16617);
  nand U17838(n16875,n16705,n16619);
  nand U17839(G4515,n16885,n16886,n16887,n16888);
  nor U17840(n16888,n16889,n16890,n16891,n16892);
  nor U17841(n16892,n16556,n16698);
  nor U17842(n16891,n16532,n16699);
  nor U17843(n16890,n16700,n16893);
  not U17844(n16893,n16894);
  nor U17845(n16889,n16895,n16703);
  nand U17846(n16887,G36441,G4389);
  nand U17847(n16886,n16704,n16557);
  nand U17848(n16885,n16705,n16559);
  nand U17849(G4514,n16896,n16897,n16898);
  nor U17850(n16898,n16899,n16900,n16901);
  nor U17851(n16901,n16902,n16703);
  nor U17852(n16900,n16799,n16903);
  nor U17853(n16899,n16640,n16699);
  not U17854(n16640,n16184);
  nand U17855(n16897,n16704,n16669);
  nand U17856(n16896,n16705,n16665);
  nand U17857(G4513,n16904,n16905,n16906,n16907);
  nor U17858(n16907,n16908,n16909,n16910,n16911);
  nor U17859(n16911,n16424,n16698);
  nor U17860(n16910,n16400,n16699);
  nor U17861(n16909,n16700,n16912);
  nor U17862(n16908,n16913,n16703);
  nand U17863(n16906,G36439,G4389);
  nand U17864(n16905,n16704,n16425);
  nand U17865(n16904,n16705,n16427);
  nand U17866(G4512,n16914,n16915,n16916,n16917);
  nor U17867(n16917,n16918,n16919,n16920,n16921);
  nor U17868(n16921,n16508,n16698);
  nor U17869(n16920,n16484,n16699);
  nor U17870(n16919,n16700,n16922);
  nor U17871(n16918,n16923,n16703);
  nand U17872(n16916,G36438,G4389);
  nand U17873(n16915,n16704,n16509);
  nand U17874(n16914,n16705,n16511);
  nand U17875(G4511,n16924,n16925,n16926,n16927);
  nor U17876(n16927,n16928,n16929,n16930,n16931);
  nor U17877(n16931,n16400,n16698);
  nor U17878(n16930,n16376,n16699);
  nor U17879(n16929,n16700,n16932);
  not U17880(n16932,n16933);
  nor U17881(n16928,n16934,n16703);
  nand U17882(n16926,G36437,G4389);
  nand U17883(n16925,n16704,n16401);
  nand U17884(n16924,n16705,n16403);
  nand U17885(G4510,n16935,n16936,n16937,n16938);
  nor U17886(n16938,n16939,n16940,n16941,n16942);
  nor U17887(n16942,n16532,n16698);
  nor U17888(n16941,n16508,n16699);
  nor U17889(n16940,n16700,n16943);
  nor U17890(n16939,n16944,n16703);
  nand U17891(n16937,G36436,G4389);
  nand U17892(G4509,n16945,n16946,n16947,n16948);
  nor U17893(n16948,n16949,n16950,n16951);
  nor U17894(n16951,n16952,n16703);
  nor U17895(n16950,n16799,n16953);
  and U17896(n16799,n16700,G36460);
  nor U17897(n16949,n16616,n16699);
  nand U17898(n16947,n16705,n16643);
  nand U17899(n16946,n16758,n16184);
  not U17900(n16758,n16698);
  nand U17901(n16945,n16704,n16641);
  nand U17902(G4508,n16954,n16955,n16956,n16957);
  nor U17903(n16957,n16958,n16959,n16960,n16961);
  nor U17904(n16961,n16448,n16698);
  nor U17905(n16960,n16424,n16699);
  nor U17906(n16959,n16700,n16962);
  not U17907(n16962,n16963);
  nor U17908(n16958,n16964,n16703);
  nand U17909(n16956,G36434,G4389);
  nand U17910(n16955,n16704,n16449);
  nand U17911(n16954,n16705,n16451);
  nand U17912(G4507,n16965,n16966,n16967,n16968);
  nor U17913(n16968,n16969,n16970,n16971,n16972);
  nor U17914(n16972,n16592,n16698);
  nor U17915(n16971,n16568,n16699);
  nor U17916(n16970,n16700,n16973);
  nor U17917(n16969,n16974,n16703);
  nand U17918(n16967,G36433,G4389);
  nand U17919(n16966,n16704,n16593);
  nand U17920(n16965,n16705,n16595);
  nand U17921(G4506,n16975,n16976,n16977,n16978);
  nor U17922(n16978,n16979,n16980,n16981,n16982);
  nor U17923(n16982,n16352,n16698);
  nor U17924(n16981,n16324,n16699);
  nor U17925(n16980,n16700,n16983);
  nor U17926(n16979,n16984,n16703);
  nand U17927(n16977,G36432,G4389);
  nand U17928(n16976,n16704,n16353);
  nand U17929(n16975,n16705,n16355);
  nand U17930(G4505,n16985,n16986,n16987,n16988);
  nor U17931(n16988,n16989,n16990,n16991,n16992);
  nor U17932(n16992,n16484,n16698);
  nand U17933(n16698,n16993,n16994,n16995);
  nor U17934(n16991,n16460,n16699);
  nand U17935(n16699,n16993,n16996,n16995);
  nor U17936(n16990,n16700,n16997);
  and U17937(n16700,n16998,n16999,n17000,n16093);
  nand U17938(n16999,n16677,n17001);
  nand U17939(n17001,n17002,n17003);
  or U17940(n17003,n17004,n16993);
  nor U17941(n17004,n17005,n17006,n17007);
  nand U17942(n16998,n16995,n17008);
  and U17943(n16995,n16677,n17009,n17010);
  nor U17944(n16989,n17011,n16703);
  nand U17945(n16703,n16677,n17012);
  nand U17946(n17012,n17013,n17014);
  nand U17947(n17014,n16993,n17006);
  nand U17948(n16987,G36431,G4389);
  nand U17949(n16986,n16704,n16485);
  not U17950(n16704,n16757);
  nand U17951(n16757,n16677,n17007,n16993);
  nand U17952(n17007,n17015,n17016,n17017,n17018);
  nand U17953(n17018,n17019,n17020);
  nor U17954(n17017,n17021,n17022);
  not U17955(n17021,n17023);
  nand U17956(n17016,n17024,n17025);
  nand U17957(n16985,n16705,n16487);
  not U17958(n16705,n16755);
  nand U17959(n16755,n16677,n17005,n16993);
  not U17960(n16993,n17008);
  nand U17961(n17008,n17026,n17027);
  nand U17962(n17005,n17028,n16667);
  nand U17963(G4504,n17029,n17030);
  nand U17964(n17030,n17031,n17032);
  nand U17965(n17032,n17033,n17034,n17035,n17036);
  nand U17966(n17036,n17037,n17038,n17039);
  nand U17967(n17038,n16663,n17023);
  or U17968(n17035,n17020,n17040,n17039);
  nand U17969(n17039,n17041,n17042,n17043,n17044);
  nor U17970(n17044,n17045,n17046,n17047,n17048);
  nand U17971(n17048,n17049,n17050,n17051,n17052);
  xor U17972(n17052,n16178,n16759);
  xor U17973(n17051,n16181,n16952);
  xor U17974(n17050,n16184,n16798);
  xor U17975(n17049,n16187,n16902);
  nand U17976(n17047,n17053,n17054,n17055,n17056);
  xor U17977(n17056,n16166,n16702);
  xor U17978(n17055,n16169,n16974);
  xor U17979(n17054,n16172,n16853);
  xor U17980(n17053,n16175,n16883);
  nand U17981(n17046,n17057,n17058,n17059,n17060);
  xor U17982(n17060,n16534,n16520);
  xor U17983(n17059,n16546,n16532);
  xor U17984(n17058,n16558,n16544);
  xor U17985(n17057,n16163,n16790);
  nand U17986(n17045,n17061,n17062,n17063,n17064);
  xor U17987(n17064,n16486,n16472);
  xor U17988(n17063,n16498,n16484);
  xor U17989(n17062,n16510,n16496);
  xor U17990(n17061,n16522,n16508);
  nor U17991(n17043,n17065,n17066,n17067,n17068);
  xor U17992(n17068,n16121,n16402);
  xor U17993(n17067,n16118,n16390);
  nand U17994(n17066,n17069,n17070);
  xor U17995(n17070,n16414,n16400);
  xor U17996(n17069,n16426,n16412);
  nand U17997(n17065,n17071,n17072,n17073,n17074);
  xor U17998(n17074,n16438,n16424);
  xor U17999(n17073,n16450,n16436);
  xor U18000(n17072,n16462,n16448);
  xor U18001(n17071,n16474,n16460);
  nor U18002(n17042,n17075,n17076,n17077,n17078);
  xor U18003(n17078,n16103,n16329);
  xor U18004(n17077,n16100,n16311);
  xor U18005(n17076,n16097,n16304);
  xor U18006(n17075,n16094,n16295);
  nor U18007(n17041,n17079,n17080,n17081,n17082);
  xor U18008(n17082,n16115,n16378);
  xor U18009(n17081,n16112,n16366);
  xor U18010(n17080,n16109,n16354);
  xor U18011(n17079,n16106,n16342);
  nand U18012(n17034,n17083,n17084);
  nand U18013(n17084,n17085,n16671);
  xor U18014(n17083,n16673,n17086);
  nand U18015(n17033,n17087,n17088,n16674);
  nand U18016(n17088,n17089,n17090);
  nand U18017(n17087,n17086,n17091);
  nand U18018(n17091,n17092,n17020);
  not U18019(n17086,n17089);
  nand U18020(n17089,n17093,n17094);
  nand U18021(n17094,n17095,n17096);
  nand U18022(n17093,n17097,n17098,n17099);
  nand U18023(n17099,n17100,n17101);
  nand U18024(n17098,n17102,n17103,n17104);
  or U18025(n17104,n17101,n17100);
  and U18026(n17100,n17105,n17106,n17107);
  nand U18027(n17107,n17108,n16097);
  nand U18028(n17106,n17109,n16304);
  nand U18029(n17105,n17110,n17111);
  nand U18030(n17101,n17112,n17113);
  nand U18031(n17113,n17109,n16097);
  nand U18032(n17112,n17114,n16304);
  nand U18033(n17103,n17115,n17116,n17117);
  nand U18034(n17117,n17118,n17119);
  nand U18035(n17116,n17120,n17121,n17122,n17123);
  or U18036(n17123,n17119,n17118);
  and U18037(n17118,n17124,n17125);
  nand U18038(n17125,n17126,n17127);
  nand U18039(n17124,n17128,n17129,n17130);
  nand U18040(n17130,n17131,n17132);
  nand U18041(n17129,n17133,n17134,n17135);
  nand U18042(n17135,n17136,n17137);
  nand U18043(n17134,n17138,n17139,n17140);
  or U18044(n17140,n17137,n17136);
  and U18045(n17136,n17141,n17142);
  nand U18046(n17142,n17109,n16112);
  nand U18047(n17141,n17114,n16366);
  nand U18048(n17137,n17143,n17144,n17145);
  nand U18049(n17145,n17108,n16112);
  nand U18050(n17144,n16365,n17146);
  nand U18051(n17143,n17109,n16366);
  nand U18052(n17139,n17147,n17148,n17149);
  nand U18053(n17149,n17150,n17151);
  nand U18054(n17148,n17152,n17153,n17154);
  or U18055(n17154,n17151,n17150);
  and U18056(n17150,n17155,n17156);
  nand U18057(n17156,n17109,n16118);
  nand U18058(n17155,n17114,n16390);
  nand U18059(n17151,n17157,n17158,n17159);
  nand U18060(n17159,n17108,n16118);
  nand U18061(n17158,n16389,n17146);
  nand U18062(n17157,n17109,n16390);
  nand U18063(n17153,n17160,n17161,n17162);
  nand U18064(n17162,n17163,n17164);
  nand U18065(n17161,n17165,n17166,n17167);
  or U18066(n17167,n17164,n17163);
  and U18067(n17163,n17168,n17169);
  nand U18068(n17169,n17109,n16124);
  nand U18069(n17168,n17114,n16414);
  nand U18070(n17164,n17170,n17171,n17172);
  nand U18071(n17172,n17108,n16124);
  nand U18072(n17171,n16413,n17146);
  nand U18073(n17170,n17109,n16414);
  nand U18074(n17166,n17173,n17174,n17175);
  nand U18075(n17175,n17176,n17177);
  nand U18076(n17174,n17178,n17179,n17180);
  or U18077(n17180,n17177,n17176);
  and U18078(n17176,n17181,n17182);
  nand U18079(n17182,n17109,n16130);
  nand U18080(n17181,n17114,n16438);
  nand U18081(n17177,n17183,n17184,n17185);
  nand U18082(n17185,n17108,n16130);
  nand U18083(n17184,n16437,n17146);
  nand U18084(n17183,n17109,n16438);
  nand U18085(n17179,n17186,n17187,n17188);
  nand U18086(n17188,n17189,n17190);
  nand U18087(n17187,n17191,n17192,n17193);
  or U18088(n17193,n17190,n17189);
  and U18089(n17189,n17194,n17195);
  nand U18090(n17195,n17109,n16136);
  nand U18091(n17194,n17114,n16462);
  nand U18092(n17190,n17196,n17197,n17198);
  nand U18093(n17198,n17108,n16136);
  nand U18094(n17197,n16461,n17146);
  nand U18095(n17196,n17109,n16462);
  nand U18096(n17192,n17199,n17200,n17201);
  nand U18097(n17201,n17202,n17203);
  nand U18098(n17200,n17204,n17205,n17206);
  or U18099(n17206,n17203,n17202);
  and U18100(n17202,n17207,n17208);
  nand U18101(n17208,n17109,n16142);
  nand U18102(n17207,n17114,n16486);
  nand U18103(n17203,n17209,n17210,n17211);
  nand U18104(n17211,n17108,n16142);
  nand U18105(n17210,n16485,n17146);
  nand U18106(n17209,n17109,n16486);
  nand U18107(n17205,n17212,n17213,n17214);
  nand U18108(n17214,n17215,n17216);
  nand U18109(n17213,n17217,n17218,n17219);
  or U18110(n17219,n17216,n17215);
  and U18111(n17215,n17220,n17221);
  nand U18112(n17221,n17109,n16148);
  nand U18113(n17220,n17114,n16510);
  nand U18114(n17216,n17222,n17223,n17224);
  nand U18115(n17224,n17108,n16148);
  nand U18116(n17223,n16509,n17146);
  nand U18117(n17222,n17109,n16510);
  nand U18118(n17218,n17225,n17226,n17227);
  nand U18119(n17227,n17228,n17229);
  nand U18120(n17226,n17230,n17231,n17232);
  or U18121(n17232,n17229,n17228);
  and U18122(n17228,n17233,n17234);
  nand U18123(n17234,n17109,n16154);
  nand U18124(n17233,n17114,n16534);
  nand U18125(n17229,n17235,n17236,n17237);
  nand U18126(n17237,n17108,n16154);
  nand U18127(n17236,n16533,n17146);
  nand U18128(n17235,n17109,n16534);
  nand U18129(n17231,n17238,n17239,n17240);
  nand U18130(n17240,n17241,n17242);
  nand U18131(n17239,n17243,n17244,n17245);
  or U18132(n17245,n17242,n17241);
  and U18133(n17241,n17246,n17247);
  nand U18134(n17247,n17109,n16160);
  nand U18135(n17246,n17114,n16558);
  nand U18136(n17242,n17248,n17249,n17250,n17251);
  nand U18137(n17251,n16557,n17146);
  nand U18138(n17249,n17109,n16558);
  nand U18139(n17248,n17108,n16160);
  nand U18140(n17244,n17252,n17253,n17254);
  nand U18141(n17254,n17255,n17256);
  nand U18142(n17253,n17257,n17258,n17259);
  or U18143(n17259,n17256,n17255);
  and U18144(n17255,n17260,n17261);
  nand U18145(n17261,n17109,n16166);
  nand U18146(n17260,n17114,n16582);
  nand U18147(n17256,n17262,n17263,n17250,n17264);
  nand U18148(n17264,n16581,n17146);
  nand U18149(n17263,n17109,n16582);
  nand U18150(n17262,n17108,n16166);
  nand U18151(n17258,n17265,n17266,n17267);
  nand U18152(n17267,n17268,n17269);
  nand U18153(n17266,n17270,n17271,n17272);
  or U18154(n17272,n17269,n17268);
  and U18155(n17268,n17273,n17274);
  nand U18156(n17274,n17109,n16172);
  nand U18157(n17273,n17114,n16606);
  nand U18158(n17269,n17275,n17276,n17250,n17277);
  nand U18159(n17277,n16605,n17146);
  nand U18160(n17276,n17109,n16606);
  nand U18161(n17275,n17108,n16172);
  nand U18162(n17271,n17278,n17279,n17280);
  nand U18163(n17280,n17281,n17282);
  nand U18164(n17279,n17283,n17284,n17285);
  or U18165(n17285,n17282,n17281);
  and U18166(n17281,n17286,n17287);
  nand U18167(n17287,n17109,n16178);
  nand U18168(n17286,n17114,n16630);
  nand U18169(n17282,n17288,n17289,n17250,n17290);
  nand U18170(n17290,n16629,n17146);
  nand U18171(n17289,n17109,n16630);
  nand U18172(n17288,n17108,n16178);
  nand U18173(n17284,n17291,n17292,n17293);
  nand U18174(n17293,n17294,n17295);
  nand U18175(n17292,n17296,n17297,n17298);
  nand U18176(n17298,n17250,n17299,n17300);
  nand U18177(n17297,n17301,n17302,n17250,n17303);
  nor U18178(n17303,n17304,n17025,n17037);
  or U18179(n17302,n17299,n17300);
  and U18180(n17300,n17305,n17306,n17307);
  nand U18181(n17307,n17108,n16187);
  nand U18182(n17306,n17109,n16662);
  nand U18183(n17305,n17110,n16669);
  nand U18184(n17299,n17308,n17309);
  nand U18185(n17309,n17109,n16187);
  nand U18186(n17308,n17114,n16662);
  nand U18187(n17301,n17310,n17311);
  or U18188(n17296,n17295,n17294);
  and U18189(n17294,n17312,n17313);
  nand U18190(n17313,n17109,n16184);
  nand U18191(n17312,n17114,n16654);
  nand U18192(n17295,n17314,n17315,n17250,n17316);
  nand U18193(n17316,n16653,n17146);
  nand U18194(n17315,n17109,n16654);
  nand U18195(n17314,n17108,n16184);
  nand U18196(n17291,n17317,n17318);
  or U18197(n17283,n17318,n17317);
  and U18198(n17317,n17319,n17320);
  nand U18199(n17320,n17109,n16181);
  nand U18200(n17319,n17114,n16642);
  nand U18201(n17318,n17250,n17321,n17322,n17323);
  nand U18202(n17323,n17109,n16642);
  nand U18203(n17322,n17110,n16641);
  nand U18204(n17321,n17108,n16181);
  nand U18205(n17278,n17324,n17325);
  or U18206(n17270,n17325,n17324);
  and U18207(n17324,n17326,n17327);
  nand U18208(n17327,n17109,n16175);
  nand U18209(n17326,n17114,n16618);
  nand U18210(n17325,n17250,n17328,n17329,n17330);
  nand U18211(n17330,n17109,n16618);
  nand U18212(n17329,n17110,n16617);
  nand U18213(n17328,n17108,n16175);
  nand U18214(n17265,n17331,n17332);
  or U18215(n17257,n17332,n17331);
  and U18216(n17331,n17333,n17334);
  nand U18217(n17334,n17109,n16169);
  nand U18218(n17333,n17114,n16594);
  nand U18219(n17332,n17250,n17335,n17336,n17337);
  nand U18220(n17337,n17109,n16594);
  nand U18221(n17336,n17110,n16593);
  nand U18222(n17335,n17108,n16169);
  nand U18223(n17252,n17338,n17339);
  or U18224(n17243,n17339,n17338);
  and U18225(n17338,n17340,n17341);
  nand U18226(n17341,n17109,n16163);
  nand U18227(n17340,n17114,n16570);
  nand U18228(n17339,n17250,n17342,n17343,n17344);
  nand U18229(n17344,n17109,n16570);
  nand U18230(n17343,n17110,n16569);
  nand U18231(n17342,n17108,n16163);
  nand U18232(n17238,n17345,n17346);
  or U18233(n17230,n17346,n17345);
  and U18234(n17345,n17347,n17348);
  nand U18235(n17348,n17109,n16157);
  nand U18236(n17347,n17114,n16546);
  nand U18237(n17346,n17349,n17350,n17351);
  nand U18238(n17351,n17108,n16157);
  nand U18239(n17350,n17109,n16546);
  nand U18240(n17349,n17110,n16545);
  nand U18241(n17225,n17352,n17353);
  or U18242(n17217,n17353,n17352);
  and U18243(n17352,n17354,n17355);
  nand U18244(n17355,n17109,n16151);
  nand U18245(n17354,n17114,n16522);
  nand U18246(n17353,n17356,n17357,n17358);
  nand U18247(n17358,n17108,n16151);
  nand U18248(n17357,n17109,n16522);
  nand U18249(n17356,n17110,n16521);
  nand U18250(n17212,n17359,n17360);
  or U18251(n17204,n17360,n17359);
  and U18252(n17359,n17361,n17362);
  nand U18253(n17362,n17109,n16145);
  nand U18254(n17361,n17114,n16498);
  nand U18255(n17360,n17363,n17364,n17365);
  nand U18256(n17365,n17108,n16145);
  nand U18257(n17364,n17109,n16498);
  nand U18258(n17363,n17110,n16497);
  nand U18259(n17199,n17366,n17367);
  or U18260(n17191,n17367,n17366);
  and U18261(n17366,n17368,n17369);
  nand U18262(n17369,n17109,n16139);
  nand U18263(n17368,n17114,n16474);
  nand U18264(n17367,n17370,n17371,n17372);
  nand U18265(n17372,n17108,n16139);
  nand U18266(n17371,n17109,n16474);
  nand U18267(n17370,n17110,n16473);
  nand U18268(n17186,n17373,n17374);
  or U18269(n17178,n17374,n17373);
  and U18270(n17373,n17375,n17376);
  nand U18271(n17376,n17109,n16133);
  nand U18272(n17375,n17114,n16450);
  nand U18273(n17374,n17377,n17378,n17379);
  nand U18274(n17379,n17108,n16133);
  nand U18275(n17378,n17109,n16450);
  nand U18276(n17377,n17110,n16449);
  nand U18277(n17173,n17380,n17381);
  or U18278(n17165,n17381,n17380);
  and U18279(n17380,n17382,n17383);
  nand U18280(n17383,n17109,n16127);
  nand U18281(n17382,n17114,n16426);
  nand U18282(n17381,n17384,n17385,n17386);
  nand U18283(n17386,n17108,n16127);
  nand U18284(n17385,n17109,n16426);
  nand U18285(n17384,n17110,n16425);
  nand U18286(n17160,n17387,n17388);
  or U18287(n17152,n17388,n17387);
  and U18288(n17387,n17389,n17390);
  nand U18289(n17390,n17109,n16121);
  nand U18290(n17389,n17114,n16402);
  nand U18291(n17388,n17391,n17392,n17393);
  nand U18292(n17393,n17108,n16121);
  nand U18293(n17392,n17109,n16402);
  nand U18294(n17391,n17110,n16401);
  nand U18295(n17147,n17394,n17395);
  or U18296(n17138,n17395,n17394);
  and U18297(n17394,n17396,n17397);
  nand U18298(n17397,n17109,n16115);
  nand U18299(n17396,n17114,n16378);
  nand U18300(n17395,n17398,n17399,n17400);
  nand U18301(n17400,n17108,n16115);
  nand U18302(n17399,n17109,n16378);
  nand U18303(n17398,n17110,n16377);
  or U18304(n17133,n17132,n17131);
  and U18305(n17131,n17401,n17402,n17403);
  nand U18306(n17403,n17108,n16109);
  nand U18307(n17402,n17109,n16354);
  nand U18308(n17401,n17110,n16353);
  nand U18309(n17132,n17404,n17405);
  nand U18310(n17405,n17109,n16109);
  nand U18311(n17404,n17114,n16354);
  or U18312(n17128,n17127,n17126);
  and U18313(n17126,n17406,n17407);
  nand U18314(n17407,n17109,n16106);
  nand U18315(n17406,n17114,n16342);
  nand U18316(n17127,n17408,n17409,n17410);
  nand U18317(n17410,n17108,n16106);
  nand U18318(n17409,n16341,n17146);
  nand U18319(n17408,n17109,n16342);
  nand U18320(n17119,n17411,n17412);
  nand U18321(n17412,n17109,n16103);
  nand U18322(n17411,n17114,n16329);
  nand U18323(n17122,n17109,n16329);
  nand U18324(n17121,n17110,n16328);
  nand U18325(n17120,n17108,n16103);
  nand U18326(n17115,n17413,n17414);
  or U18327(n17102,n17414,n17413);
  and U18328(n17413,n17415,n17416,n17417);
  nand U18329(n17417,n17108,n16100);
  nand U18330(n17416,n16314,n17146);
  nand U18331(n17146,n17250,n17418);
  nand U18332(n17415,n17109,n16311);
  nand U18333(n17414,n17419,n17420);
  nand U18334(n17420,n17109,n16100);
  nand U18335(n17419,n17114,n16311);
  or U18336(n17097,n17096,n17095);
  and U18337(n17095,n17421,n17422,n17423);
  nand U18338(n17423,n17108,n16094);
  nand U18339(n17424,n17425,n16097,n17426);
  nand U18340(n17422,n17110,n17427);
  xor U18341(n17427,n17428,n17429);
  xnor U18342(n17429,n17111,n17430);
  and U18343(n17111,n17431,n17432);
  nand U18344(n17431,n17433,n17434);
  not U18345(n17110,n17418);
  nand U18346(n17418,n16097,n17435,n17425);
  not U18347(n17425,n16094);
  nand U18348(n17421,n17109,n16295);
  nand U18349(n17096,n17436,n17437);
  nand U18350(n17437,n17109,n16094);
  nand U18351(n17438,n17009,n17250,n17010);
  nand U18352(n17015,n17439,n17092);
  nand U18353(n17436,n17114,n16295);
  and U18354(n17426,n17441,n16667,n17020);
  nand U18355(n17441,n17439,n17310);
  not U18356(n17440,n17435);
  nand U18357(n17435,n17442,n17443,n17040);
  nor U18358(n17040,n17019,n17444);
  nand U18359(n17442,n17025,n17037);
  nand U18360(n17029,n17445,n17446,G36430);
  nand U18361(n17446,n17447,n16652,n17010,n16677);
  not U18362(n16652,n16325);
  nand U18363(n17445,n17031,n17092);
  not U18364(n17031,n17000);
  nand U18365(G4503,n17448,n17449,n17450,n17451);
  nor U18366(n17451,n17452,n17453);
  and U18367(n17453,n17454,G36397);
  and U18368(n17452,n17455,n16669);
  nand U18369(n17450,G36440,G4389);
  nand U18370(n17449,G36218,n17456);
  nand U18371(n17456,n17457,n17458);
  or U18372(n17458,n17459,n17460);
  nand U18373(n17448,n17461,n17459,n17462);
  nand U18374(G4502,n17463,n17464,n17465,n17466);
  nand U18375(n17466,n16653,n17455);
  nand U18376(n17465,G36396,n17454);
  nand U18377(n17464,G36450,G4389);
  nor U18378(n17463,n17467,n17468);
  nor U18379(n17468,n17469,n17460,n17470);
  nor U18380(n17467,n17471,n17472);
  nor U18381(n17471,n17473,n17474);
  and U18382(n17473,n17470,n17461);
  nand U18383(n17470,n17475,n17476);
  nand U18384(G4501,n17477,n17478,n17479,n17480);
  nor U18385(n17480,n17481,n17482);
  nor U18386(n17482,G36460,n16953);
  not U18387(n16953,G36435);
  nor U18388(n17481,n17483,n17484);
  nand U18389(n17479,n16641,n17455);
  nand U18390(n17478,n17461,n17485);
  xnor U18391(n17485,n17486,n17487);
  xor U18392(n17487,n17488,n17489);
  nand U18393(n17477,n17474,n17490);
  nand U18394(G4500,n17491,n17492,n17493,n17494);
  nor U18395(n17494,n17495,n16750);
  nor U18396(n16750,G36460,n17496);
  nor U18397(n17495,n17483,n17497);
  nand U18398(n17493,n16629,n17455);
  nand U18399(n17492,n17498,n17461);
  xor U18400(n17498,n17499,n17500);
  xor U18401(n17500,n17501,n17502);
  nand U18402(n17491,n17474,n17502);
  nand U18403(G4499,n17503,n17504,n17505,n17506);
  nor U18404(n17506,n17507,n17508);
  nor U18405(n17508,G36460,n17509);
  and U18406(n17507,n17454,G36393);
  nand U18407(n17505,n16617,n17455);
  nand U18408(n17504,n17461,n17510);
  xor U18409(n17510,n17511,n17512);
  and U18410(n17512,n17513,n17514);
  nand U18411(n17503,n17474,n17515);
  nand U18412(G4498,n17516,n17517,n17518,n17519);
  nor U18413(n17519,n17520,n17521);
  and U18414(n17521,G4389,G36445);
  and U18415(n17520,n17454,G36392);
  nand U18416(n17518,n16605,n17455);
  nand U18417(n17517,n17522,n17461);
  xor U18418(n17522,n17523,n17524);
  and U18419(n17524,n17525,n17526);
  nand U18420(n17516,n17474,n17527);
  nand U18421(G4497,n17528,n17529,n17530,n17531);
  nor U18422(n17531,n17532,n17533);
  nor U18423(n17533,G36460,n17534);
  and U18424(n17532,n17454,G36391);
  nand U18425(n17530,n16593,n17455);
  nand U18426(n17529,n17535,n17461);
  xor U18427(n17535,n17536,n17537);
  and U18428(n17537,n17538,n17539);
  nand U18429(n17528,n17474,n17540);
  nand U18430(G4496,n17541,n17542,n17543,n17544);
  nor U18431(n17544,n17545,n17546);
  nor U18432(n17546,G36460,n17547);
  nor U18433(n17545,n17483,n17548);
  nand U18434(n17543,n16581,n17455);
  nand U18435(n17542,n17549,n17461);
  xor U18436(n17549,n17550,n17551);
  xor U18437(n17551,n17552,n17553);
  nand U18438(n17541,n17474,n17553);
  nand U18439(G4495,n17554,n17555,n17556,n17557);
  nor U18440(n17557,n17558,n17559);
  and U18441(n17559,G4389,G36451);
  nor U18442(n17558,n17483,n17560);
  nand U18443(n17556,n16569,n17455);
  nand U18444(n17555,n17461,n17561);
  xnor U18445(n17561,n17562,n17563);
  xor U18446(n17563,n17564,n17565);
  nand U18447(n17554,n17474,n17566);
  nand U18448(G4494,n17567,n17568,n17569,n17570);
  nor U18449(n17570,n17571,n17572);
  nor U18450(n17572,G36460,n17573);
  nor U18451(n17571,n17483,n17574);
  nand U18452(n17569,n16557,n17455);
  nand U18453(n17568,n17575,n17461);
  xnor U18454(n17575,n17576,n17577);
  xor U18455(n17577,n17578,n17579);
  nand U18456(n17567,n17474,n17580);
  nand U18457(G4493,n17581,n17582,n17583,n17584);
  nor U18458(n17584,n17585,n17586);
  and U18459(n17586,G4389,G36455);
  nor U18460(n17585,n17483,n17587);
  nand U18461(n17583,n16545,n17455);
  nand U18462(n17582,n17461,n17588);
  xnor U18463(n17588,n17589,n17590);
  nand U18464(n17590,n17591,n17592);
  nand U18465(n17581,n17474,n17593);
  nand U18466(G4492,n17594,n17595,n17596,n17597);
  nor U18467(n17597,n17598,n17599);
  nor U18468(n17599,G36460,n17600);
  nor U18469(n17598,n17483,n17601);
  nand U18470(n17596,n16533,n17455);
  nand U18471(n17595,n17602,n17603,n17461);
  nand U18472(n17603,n17604,n17591,n17605);
  xor U18473(n17605,n17606,n17607);
  nand U18474(n17602,n17608,n17609);
  not U18475(n17608,n17610);
  nand U18476(n17594,n17474,n17611);
  nand U18477(G4491,n17612,n17613,n17614,n17615);
  nor U18478(n17615,n17616,n17617);
  nor U18479(n17617,G36460,n17618);
  nor U18480(n17616,n17483,n17619);
  nand U18481(n17614,n16521,n17455);
  nand U18482(n17613,n17461,n17620);
  xnor U18483(n17620,n17621,n17622);
  xor U18484(n17622,n17623,n17624);
  nand U18485(n17612,n17474,n17625);
  nand U18486(G4490,n17626,n17627,n17628,n17629);
  nor U18487(n17629,n17630,n17631);
  and U18488(n17631,G4389,G36438);
  nor U18489(n17630,n17483,n17632);
  nand U18490(n17628,n16509,n17455);
  nand U18491(n17627,n17633,n17461);
  xor U18492(n17633,n17634,n17635);
  xor U18493(n17635,n17636,n17637);
  nand U18494(n17626,n17474,n17637);
  nand U18495(G4489,n17638,n17639,n17640,n17641);
  nor U18496(n17641,n17642,n17643);
  nor U18497(n17643,G36460,n17644);
  nor U18498(n17642,n17483,n17645);
  nand U18499(n17640,n16497,n17455);
  nand U18500(n17639,n17646,n17461);
  xnor U18501(n17646,n17647,n17648);
  xnor U18502(n17647,n17649,n17650);
  nand U18503(n17638,n17474,n17650);
  nand U18504(G4488,n17651,n17652,n17653,n17654);
  nor U18505(n17654,n17655,n17656);
  and U18506(n17656,G4389,G36431);
  nor U18507(n17655,n17483,n17657);
  nand U18508(n17653,n16485,n17455);
  nand U18509(n17652,n17658,n17461);
  xor U18510(n17658,n17659,n17660);
  and U18511(n17660,n17661,n17662);
  nand U18512(n17651,n17474,n17663);
  nand U18513(G4487,n17664,n17665,n17666,n17667);
  nor U18514(n17667,n17668,n17669);
  nor U18515(n17669,G36460,n17670);
  nor U18516(n17668,n17483,n17671);
  nand U18517(n17666,n16473,n17455);
  nand U18518(n17665,n17461,n17672);
  xnor U18519(n17672,n17673,n17674);
  xnor U18520(n17674,n17675,n17676);
  nand U18521(n17664,n17474,n17676);
  nand U18522(G4486,n17677,n17678,n17679,n17680);
  nor U18523(n17680,n17681,n17682);
  nor U18524(n17682,G36460,n17683);
  and U18525(n17681,n17454,G36380);
  not U18526(n17454,n17483);
  nand U18527(n17679,n16461,n17455);
  nand U18528(n17678,n17684,n17461);
  xor U18529(n17684,n17685,n17686);
  xor U18530(n17686,n17687,n17688);
  nand U18531(n17677,n17474,n17688);
  nand U18532(G4485,n17689,n17690,n17691,n17692);
  nor U18533(n17692,n17693,n17694);
  nor U18534(n17694,G36460,n17695);
  nor U18535(n17693,n17483,n17696);
  nand U18536(n17691,n16449,n17455);
  nand U18537(n17690,n17697,n17698,n17461);
  nand U18538(n17698,n17699,n17700,n17701);
  nand U18539(n17697,n17702,n17703);
  xnor U18540(n17702,n17704,n17705);
  nand U18541(n17689,n17474,n17701);
  nand U18542(G4484,n17706,n17707,n17708,n17709);
  nor U18543(n17709,n17710,n17711);
  and U18544(n17711,G4389,G36453);
  nor U18545(n17710,n17712,n17483);
  nand U18546(n17708,n16437,n17455);
  nand U18547(n17455,n17713,n17714);
  nand U18548(n17714,n16677,n17715,n16994,n17483);
  nand U18549(n17713,G4591,n16994);
  nand U18550(n17707,n17716,n17717,n17461);
  not U18551(n17461,n17460);
  nand U18552(n17460,n16994,n17483,n17718);
  nand U18553(n17718,n17000,n17719);
  nand U18554(n17719,n16677,n17720);
  nand U18555(n17717,n17721,n17700,n17722);
  not U18556(n17722,n17723);
  nand U18557(n17721,n17701,n17699);
  nand U18558(n17716,n17724,n17699,n17723);
  nand U18559(n17723,n17725,n17726);
  nand U18560(n17726,n17727,n17447);
  xor U18561(n17727,G36365,n16673);
  nand U18562(n17725,n17728,n17729);
  xor U18563(n17728,G36333,n16673);
  or U18564(n17699,n17704,n17705);
  nand U18565(n17724,n17703,n17700);
  nand U18566(n17700,n17705,n17704);
  nand U18567(n17704,n17730,n17731);
  nand U18568(n17731,n17688,n17732);
  or U18569(n17732,n17685,n17687);
  nand U18570(n17730,n17685,n17687);
  nand U18571(n17687,n17733,n17734);
  nand U18572(n17734,n17676,n17735);
  or U18573(n17735,n17673,n17675);
  nand U18574(n17733,n17673,n17675);
  nand U18575(n17675,n17661,n17736);
  nand U18576(n17736,n17662,n17659);
  nand U18577(n17659,n17737,n17738);
  nand U18578(n17738,n17650,n17739);
  or U18579(n17739,n17648,n17649);
  nand U18580(n17737,n17649,n17648);
  nand U18581(n17648,n17740,n17741);
  nand U18582(n17741,n17447,G36360);
  nand U18583(n17740,n17729,G36328);
  and U18584(n17649,n17742,n17743);
  nand U18585(n17743,n17744,n17745);
  nand U18586(n17744,n17634,n17636);
  or U18587(n17742,n17634,n17636);
  nand U18588(n17636,n17746,n17747);
  nand U18589(n17747,n17625,n17748);
  or U18590(n17748,n17621,n17623);
  nand U18591(n17746,n17621,n17623);
  nand U18592(n17623,n17610,n17609);
  nand U18593(n17609,n17611,n17607);
  nand U18594(n17610,n17749,n17750);
  nand U18595(n17750,n17604,n17591);
  nand U18596(n17591,n17751,n17752,n17593);
  or U18597(n17752,n17447,G36324);
  or U18598(n17751,n17729,G36356);
  nand U18599(n17604,n17589,n17592);
  nand U18600(n17592,n17753,n17754,n17755);
  nand U18601(n17754,n17447,G36356);
  nand U18602(n17753,n17729,G36324);
  and U18603(n17589,n17756,n17757);
  nand U18604(n17757,n17758,n17578);
  or U18605(n17758,n17576,n17579);
  nand U18606(n17756,n17576,n17579);
  nand U18607(n17579,n17759,n17760);
  nand U18608(n17760,n17565,n17761);
  nand U18609(n17761,n17562,n17564);
  or U18610(n17759,n17562,n17564);
  nand U18611(n17564,n17762,n17763);
  nand U18612(n17763,n17553,n17764);
  or U18613(n17764,n17550,n17552);
  nand U18614(n17762,n17550,n17552);
  nand U18615(n17552,n17538,n17765);
  nand U18616(n17765,n17539,n17536);
  nand U18617(n17536,n17525,n17766);
  nand U18618(n17766,n17526,n17523);
  nand U18619(n17523,n17513,n17767);
  nand U18620(n17767,n17511,n17514);
  nand U18621(n17514,n17768,n17769,n17770);
  nand U18622(n17769,n17447,G36350);
  nand U18623(n17768,n17729,G36318);
  and U18624(n17511,n17771,n17772);
  nand U18625(n17772,n17773,n17774);
  nand U18626(n17773,n17499,n17501);
  or U18627(n17771,n17499,n17501);
  nand U18628(n17501,n17775,n17776);
  nand U18629(n17776,n17490,n17777);
  or U18630(n17777,n17486,n17488);
  nand U18631(n17775,n17486,n17488);
  nand U18632(n17488,n17475,n17778);
  nand U18633(n17778,n17469,n17476);
  nand U18634(n17476,n17779,n17780);
  nand U18635(n17780,G36218,n17459);
  not U18636(n17779,n17781);
  nand U18637(n17475,n17781,n17459,G36218);
  nand U18638(n17459,n17782,n17783);
  nand U18639(n17783,n17447,G36346);
  nand U18640(n17782,n17729,G36314);
  nand U18641(n17781,n17784,n17785);
  nand U18642(n17785,n17447,G36347);
  nand U18643(n17784,n17729,G36315);
  nand U18644(n17486,n17786,n17787);
  nand U18645(n17787,n17447,G36348);
  nand U18646(n17786,n17729,G36316);
  nand U18647(n17499,n17788,n17789);
  nand U18648(n17789,n17447,G36349);
  nand U18649(n17788,n17729,G36317);
  nand U18650(n17513,n17790,n17791,n17515);
  or U18651(n17791,n17447,G36318);
  or U18652(n17790,n17729,G36350);
  nand U18653(n17526,n17792,n17793,n17794);
  nand U18654(n17793,n17447,G36351);
  nand U18655(n17792,n17729,G36319);
  nand U18656(n17525,n17795,n17796,n17527);
  or U18657(n17796,n17447,G36319);
  or U18658(n17795,n17729,G36351);
  nand U18659(n17539,n17797,n17798,n17799);
  nand U18660(n17798,n17447,G36352);
  nand U18661(n17797,n17729,G36320);
  nand U18662(n17538,n17800,n17801,n17540);
  or U18663(n17801,n17447,G36320);
  or U18664(n17800,n17729,G36352);
  nand U18665(n17550,n17802,n17803);
  nand U18666(n17803,n17447,G36353);
  nand U18667(n17802,n17729,G36321);
  nand U18668(n17562,n17804,n17805);
  nand U18669(n17805,n17447,G36354);
  nand U18670(n17804,n17729,G36322);
  nand U18671(n17576,n17806,n17807);
  or U18672(n17807,n17447,G36323);
  or U18673(n17806,n17729,G36355);
  or U18674(n17749,n17607,n17611);
  nand U18675(n17607,n17808,n17809);
  nand U18676(n17809,n17447,G36357);
  nand U18677(n17808,n17729,G36325);
  nand U18678(n17621,n17810,n17811);
  nand U18679(n17811,n17447,G36358);
  nand U18680(n17810,n17729,G36326);
  nand U18681(n17634,n17812,n17813);
  nand U18682(n17813,n17447,G36359);
  nand U18683(n17812,n17729,G36327);
  nand U18684(n17662,n17814,n17815,n17816);
  nand U18685(n17815,n17447,G36361);
  nand U18686(n17814,n17729,G36329);
  nand U18687(n17661,n17817,n17818,n17663);
  nand U18688(n17818,n17729,n17819);
  nand U18689(n17817,n17447,n17820);
  nand U18690(n17673,n17821,n17822);
  nand U18691(n17822,n17447,G36362);
  nand U18692(n17821,n17729,G36330);
  nand U18693(n17685,n17823,n17824);
  nand U18694(n17824,n17447,G36363);
  nand U18695(n17823,n17729,G36331);
  nand U18696(n17705,n17825,n17826);
  nand U18697(n17826,n17447,G36364);
  nand U18698(n17825,n17729,G36332);
  nand U18699(n17706,n17474,n16673);
  not U18700(n17474,n17457);
  nand U18701(n17457,n16996,n17827);
  nand U18702(n17827,n17828,n16093);
  nand U18703(n17828,n17483,n17830);
  nand U18704(n17830,n17831,n17000);
  nand U18705(n17000,n17250,G36460);
  nand U18706(n17831,n16677,n17832);
  or U18707(n17832,n17715,n17720);
  nand U18708(n17720,n17833,n17443,n16671,n17834);
  nand U18709(n17715,n17835,n16668);
  nand U18710(n17483,n17836,n17829,n17837);
  nand U18711(n17836,n17838,n17090);
  nand U18712(G4483,n17839,n17840,n17841);
  nand U18713(n17841,n17842,n16295);
  nand U18714(n17840,G36377,n17843);
  nand U18715(n17839,n17844,n17845);
  nand U18716(n17845,n16292,n17846);
  nand U18717(n17846,n17847,n16297);
  xnor U18718(n16297,n16295,n17848);
  nand U18719(n16295,n17849,n17850);
  nand U18720(n17850,n17851,G36184);
  nand U18721(n17849,n17852,n17853);
  nand U18722(G4482,n17854,n17855,n17856);
  nand U18723(n17856,n17842,n16304);
  nand U18724(n17855,G36376,n17843);
  nand U18725(n17854,n17844,n17857);
  nand U18726(n17857,n16292,n17858);
  nand U18727(n17858,n17847,n16303);
  nor U18728(n16303,n17859,n17848);
  nor U18729(n17848,n17860,n17861);
  and U18730(n17861,n17862,n17863);
  and U18731(n17859,n17860,n17862);
  nand U18732(n17862,n17864,n17865);
  nand U18733(n17864,n16304,n17866);
  nand U18734(n16304,n17867,n17868);
  nand U18735(n17868,n17851,G36183);
  nand U18736(n17867,n17852,n17869);
  nand U18737(n17860,n17870,n17871);
  not U18738(n17847,n17872);
  nand U18739(n16292,n16094,n17873);
  nand U18740(n17873,n17874,n17875);
  nand U18741(n17875,n16675,n17876);
  nand U18742(n17874,n17877,n17009);
  nand U18743(n16094,n17878,n17879,n17880);
  nand U18744(n17880,G36313,n17881);
  nand U18745(n17879,G36377,n17882);
  nand U18746(n17878,G36345,n17883);
  nand U18747(G4481,n17884,n17885,n17886,n17887);
  nor U18748(n17887,n17888,n17889,n17890);
  nor U18749(n17890,n17843,n16310);
  nand U18750(n16310,n17891,n17892,n17009);
  nand U18751(n17892,n17893,n16996);
  nand U18752(n17893,n16097,n17894);
  nand U18753(n17894,G36430,n17838);
  nand U18754(n16097,n17895,n17896,n17897);
  nand U18755(n17897,G36312,n17881);
  nand U18756(n17896,G36376,n17882);
  nand U18757(n17895,G36344,n17883);
  nand U18758(n17891,n16340,n16994);
  and U18759(n17889,n17843,G36375);
  and U18760(n17888,n16311,n17842);
  nand U18761(n17886,n17898,n16314);
  xor U18762(n16314,n17433,n17899);
  and U18763(n17899,n17434,n17432);
  nand U18764(n17432,n17900,n17901);
  nand U18765(n17901,n17430,n17902);
  not U18766(n17900,n17428);
  nand U18767(n17434,n17428,n17902,n17430);
  and U18768(n17430,n17903,n17904,n17905,n17906);
  nor U18769(n17906,n17907,n17908);
  and U18770(n17907,n16100,n17909);
  nand U18771(n17905,n17910,n16329);
  nand U18772(n17904,n16311,n17911);
  nand U18773(n17903,n17912,n16103);
  nand U18774(n17902,n17250,n16100);
  xor U18775(n17428,n17913,n17914);
  nand U18776(n17913,n17915,n17916,n17917,n17918);
  nor U18777(n17918,n17919,n17920);
  nor U18778(n17920,n16340,n17921);
  nor U18779(n17919,n16780,n17922);
  nand U18780(n17917,n17909,n16311);
  nand U18781(n17915,n17911,n16100);
  nand U18782(n17911,n17923,n17924);
  nand U18783(n17433,n17925,n17926);
  nand U18784(n17926,n17927,n17928);
  nand U18785(n17884,n17931,n16312);
  xor U18786(n16312,n17871,n17932);
  nor U18787(n17932,n17933,n17934);
  not U18788(n17934,n17870);
  nand U18789(n17870,n17865,n17863,n17935);
  nand U18790(n17935,n17936,n17937);
  nand U18791(n17936,n17866,n16311);
  nor U18792(n17933,n17863,n17865);
  nand U18793(n17865,n17938,n16100);
  nand U18794(n17863,n16311,n17938);
  nand U18795(n17938,n17939,n17940);
  nand U18796(n16311,n17941,n17942);
  nand U18797(n17942,n17851,G36182);
  nand U18798(n17941,n17852,n17943);
  nand U18799(n17871,n17944,n17945);
  nand U18800(n17945,n17946,n17947);
  nand U18801(G4480,n17948,n17949,n17950,n17951);
  nor U18802(n17951,n17952,n17953,n17954,n17955);
  nor U18803(n17955,n16780,n17956);
  not U18804(n16780,n16329);
  and U18805(n17954,n16330,n17931);
  xor U18806(n16330,n17947,n17957);
  and U18807(n17957,n17946,n17944);
  nand U18808(n17944,n16329,n17085,n17958);
  nand U18809(n17946,n17959,n17960);
  nand U18810(n17960,n16329,n17085);
  xor U18811(n17959,n17085,n17958);
  nand U18812(n17958,n17961,n17962);
  nand U18813(n17962,n16329,n17937);
  nand U18814(n17961,n16103,n17085);
  nand U18815(n17947,n17963,n17964);
  nand U18816(n17964,n17965,n17966);
  and U18817(n17953,n16328,n17898);
  xor U18818(n16328,n17928,n17967);
  and U18819(n17967,n17927,n17925);
  nand U18820(n17925,n17968,n17969);
  or U18821(n17927,n17968,n17969);
  nand U18822(n17969,n17970,n17971,n17972);
  nand U18823(n17971,n16329,n17973);
  nand U18824(n17970,n17974,n16103);
  xor U18825(n17968,n17975,n17976);
  nand U18826(n17975,n17977,n17916,n17978);
  nand U18827(n17978,n16103,n17973);
  nand U18828(n17977,n16329,n17979);
  nand U18829(n16329,n17980,n17981);
  nand U18830(n17981,n17851,G36181);
  nand U18831(n17980,n17852,n17982);
  nand U18832(n17928,n17983,n17984);
  nand U18833(n17984,n17985,n17986);
  nor U18834(n17952,n16326,n17987);
  not U18835(n16326,n16100);
  nand U18836(n16100,n17988,n17989,n17990,n17991);
  nand U18837(n17991,n17930,n17992);
  nand U18838(n17990,G36375,n17882);
  nand U18839(n17989,G36343,n17883);
  nand U18840(n17988,G36311,n17881);
  nand U18841(n17950,G36374,n17843);
  nand U18842(G4479,n17994,n17995,n17996,n17997);
  nor U18843(n17997,n17998,n17999,n18000,n18001);
  nor U18844(n18001,n16715,n17956);
  not U18845(n16715,n16342);
  and U18846(n18000,n16343,n17931);
  xor U18847(n16343,n17966,n18002);
  and U18848(n18002,n17965,n17963);
  nand U18849(n17963,n16342,n17085,n18003);
  nand U18850(n17965,n18004,n18005);
  nand U18851(n18005,n16342,n17085);
  xor U18852(n18004,n17085,n18003);
  nand U18853(n18003,n18006,n18007);
  nand U18854(n18007,n16342,n17937);
  nand U18855(n18006,n16106,n17085);
  nand U18856(n17966,n18008,n18009);
  nand U18857(n18009,n18010,n18011);
  and U18858(n17999,n16341,n17898);
  xor U18859(n16341,n17986,n18012);
  and U18860(n18012,n17985,n17983);
  nand U18861(n17983,n18013,n18014);
  or U18862(n17985,n18013,n18014);
  nand U18863(n18014,n18015,n18016,n17972);
  nand U18864(n18016,n16342,n17973);
  nand U18865(n18015,n17974,n16106);
  xor U18866(n18013,n18017,n17976);
  nand U18867(n18017,n18018,n17916,n18019);
  nand U18868(n18019,n16106,n17973);
  nand U18869(n18018,n16342,n17979);
  nand U18870(n16342,n18020,n18021);
  nand U18871(n18021,n17851,G36180);
  nand U18872(n18020,n18022,n17852);
  nand U18873(n17986,n18023,n18024);
  nand U18874(n18024,n18025,n18026);
  nor U18875(n17998,n16340,n17987);
  not U18876(n16340,n16103);
  nand U18877(n16103,n18027,n18028,n18029,n18030);
  nand U18878(n18030,n16779,n17992);
  nor U18879(n16779,n17930,n18031);
  and U18880(n18031,n18032,n18033);
  nor U18881(n17930,n18033,n18032);
  not U18882(n18033,G36452);
  nand U18883(n18029,G36374,n17882);
  nand U18884(n18028,G36342,n17883);
  nand U18885(n18027,G36310,n17881);
  nand U18886(n17996,G36373,n17843);
  nand U18887(G4478,n18035,n18036,n18037,n18038);
  nor U18888(n18038,n18039,n18040,n18041,n18042);
  nor U18889(n18042,n16984,n17956);
  not U18890(n16984,n16354);
  and U18891(n18041,n16355,n17931);
  xor U18892(n16355,n18011,n18043);
  and U18893(n18043,n18010,n18008);
  nand U18894(n18008,n16354,n17085,n18044);
  nand U18895(n18010,n18045,n18046);
  nand U18896(n18046,n16354,n17085);
  xor U18897(n18045,n17085,n18044);
  nand U18898(n18044,n18047,n18048);
  nand U18899(n18048,n16354,n17937);
  nand U18900(n18047,n16109,n17085);
  nand U18901(n18011,n18049,n18050);
  nand U18902(n18050,n18051,n18052);
  and U18903(n18040,n16353,n17898);
  xor U18904(n16353,n18026,n18053);
  and U18905(n18053,n18025,n18023);
  nand U18906(n18023,n18054,n18055);
  or U18907(n18025,n18054,n18055);
  nand U18908(n18055,n18056,n18057,n17972);
  nand U18909(n18057,n16354,n17973);
  nand U18910(n18056,n17974,n16109);
  xor U18911(n18054,n18058,n17976);
  nand U18912(n18058,n18059,n17916,n18060);
  nand U18913(n18060,n16109,n17973);
  nand U18914(n18059,n16354,n17979);
  nand U18915(n16354,n18061,n18062);
  nand U18916(n18062,n17851,G36179);
  nand U18917(n18061,n18063,n17852);
  nand U18918(n18026,n18064,n18065);
  nand U18919(n18065,n18066,n18067);
  nor U18920(n18039,n16324,n17987);
  not U18921(n16324,n16106);
  nand U18922(n16106,n18068,n18069,n18070,n18071);
  nand U18923(n18071,n18034,n17992);
  not U18924(n18034,n16714);
  nand U18925(n16714,n18072,n18032);
  or U18926(n18032,n18073,n18074);
  nand U18927(n18072,n18073,n18074);
  nand U18928(n18074,G36432,n18075,G36447);
  not U18929(n18073,G36458);
  nand U18930(n18070,G36373,n17882);
  nand U18931(n18069,G36341,n17883);
  nand U18932(n18068,G36309,n17881);
  nand U18933(n18037,G36372,n17843);
  nand U18934(G4477,n18077,n18078,n18079,n18080);
  nor U18935(n18080,n18081,n18082,n18083,n18084);
  nor U18936(n18084,n16833,n17956);
  not U18937(n16833,n16366);
  and U18938(n18083,n16367,n17931);
  xor U18939(n16367,n18052,n18085);
  and U18940(n18085,n18051,n18049);
  nand U18941(n18049,n16366,n17085,n18086);
  nand U18942(n18051,n18087,n18088);
  nand U18943(n18088,n16366,n17085);
  xor U18944(n18087,n17085,n18086);
  nand U18945(n18086,n18089,n18090);
  nand U18946(n18090,n16366,n17937);
  nand U18947(n18089,n16112,n17085);
  nand U18948(n18052,n18091,n18092);
  nand U18949(n18092,n18093,n18094);
  and U18950(n18082,n16365,n17898);
  xor U18951(n16365,n18067,n18095);
  and U18952(n18095,n18066,n18064);
  nand U18953(n18064,n18096,n18097);
  or U18954(n18066,n18096,n18097);
  nand U18955(n18097,n18098,n18099,n17972);
  nand U18956(n18099,n16366,n17973);
  nand U18957(n18098,n17974,n16112);
  xor U18958(n18096,n18100,n17976);
  nand U18959(n18100,n18101,n17916,n18102);
  nand U18960(n18102,n16112,n17973);
  nand U18961(n18101,n16366,n17979);
  nand U18962(n16366,n18103,n18104);
  nand U18963(n18104,n17851,G36178);
  nand U18964(n18103,n18105,n17852);
  nand U18965(n18067,n18106,n18107);
  nand U18966(n18107,n18108,n18109);
  nor U18967(n18081,n16339,n17987);
  not U18968(n16339,n16109);
  nand U18969(n16109,n18110,n18111,n18112,n18113);
  nand U18970(n18113,n18076,n17992);
  not U18971(n18076,n16983);
  xor U18972(n16983,n18114,G36432);
  nand U18973(n18114,G36447,n18075);
  nand U18974(n18112,G36372,n17882);
  nand U18975(n18111,G36340,n17883);
  nand U18976(n18110,G36308,n17881);
  nand U18977(n18079,G36371,n17843);
  nand U18978(G4476,n18115,n18116,n18117,n18118);
  nor U18979(n18118,n18119,n18120,n18121,n18122);
  nor U18980(n18122,n16874,n17956);
  not U18981(n16874,n16378);
  and U18982(n18121,n16379,n17931);
  xor U18983(n16379,n18094,n18123);
  and U18984(n18123,n18093,n18091);
  nand U18985(n18091,n16378,n17085,n18124);
  nand U18986(n18093,n18125,n18126);
  nand U18987(n18126,n16378,n17085);
  xor U18988(n18125,n17085,n18124);
  nand U18989(n18124,n18127,n18128);
  nand U18990(n18128,n16378,n17937);
  nand U18991(n18127,n16115,n17085);
  nand U18992(n18094,n18129,n18130);
  nand U18993(n18130,n18131,n18132);
  and U18994(n18120,n16377,n17898);
  xor U18995(n16377,n18109,n18133);
  and U18996(n18133,n18108,n18106);
  nand U18997(n18106,n18134,n18135);
  or U18998(n18108,n18134,n18135);
  nand U18999(n18135,n18136,n18137,n17972);
  nand U19000(n18137,n16378,n17973);
  nand U19001(n18136,n17974,n16115);
  xor U19002(n18134,n18138,n17976);
  nand U19003(n18138,n18139,n17916,n18140);
  nand U19004(n18140,n16115,n17973);
  nand U19005(n18139,n16378,n17979);
  nand U19006(n16378,n18141,n18142);
  nand U19007(n18142,n17851,G36177);
  nand U19008(n18141,n18143,n17852);
  nand U19009(n18109,n18144,n18145);
  nand U19010(n18145,n18146,n18147);
  nor U19011(n18119,n16352,n17987);
  not U19012(n16352,n16112);
  nand U19013(n16112,n18148,n18149,n18150,n18151);
  nand U19014(n18151,n16832,n17992);
  xor U19015(n16832,G36447,n18075);
  not U19016(n18075,n18152);
  nand U19017(n18150,G36371,n17882);
  nand U19018(n18149,G36339,n17883);
  nand U19019(n18148,G36307,n17881);
  nand U19020(n18117,G36370,n17843);
  nand U19021(G4475,n18154,n18155,n18156,n18157);
  nor U19022(n18157,n18158,n18159,n18160,n18161);
  nor U19023(n18161,n16735,n17956);
  not U19024(n16735,n16390);
  and U19025(n18160,n16391,n17931);
  xor U19026(n16391,n18132,n18162);
  and U19027(n18162,n18131,n18129);
  nand U19028(n18129,n16390,n17085,n18163);
  nand U19029(n18131,n18164,n18165);
  nand U19030(n18165,n16390,n17085);
  xor U19031(n18164,n17085,n18163);
  nand U19032(n18163,n18166,n18167);
  nand U19033(n18167,n16390,n17937);
  nand U19034(n18166,n16118,n17085);
  nand U19035(n18132,n18168,n18169);
  nand U19036(n18169,n18170,n18171);
  and U19037(n18159,n16389,n17898);
  xor U19038(n16389,n18147,n18172);
  and U19039(n18172,n18146,n18144);
  nand U19040(n18144,n18173,n18174);
  or U19041(n18146,n18173,n18174);
  nand U19042(n18174,n18175,n18176,n17972);
  nand U19043(n18176,n16390,n17973);
  nand U19044(n18175,n17974,n16118);
  xor U19045(n18173,n18177,n17976);
  nand U19046(n18177,n18178,n17916,n18179);
  nand U19047(n18179,n16118,n17973);
  nand U19048(n18178,n16390,n17979);
  nand U19049(n16390,n18180,n18181);
  nand U19050(n18181,n17851,G36176);
  nand U19051(n18180,n18182,n17852);
  nand U19052(n18147,n18183,n18184);
  nand U19053(n18184,n18185,n18186);
  nor U19054(n18158,n16364,n17987);
  not U19055(n16364,n16115);
  nand U19056(n16115,n18187,n18188,n18189,n18190);
  nand U19057(n18190,n18153,n17992);
  not U19058(n18153,n16873);
  nand U19059(n16873,n18191,n18152);
  nand U19060(n18152,G36443,n18192,G36456);
  nand U19061(n18191,n18193,n18194);
  nand U19062(n18194,G36456,n18192);
  not U19063(n18193,G36443);
  nand U19064(n18189,G36370,n17882);
  nand U19065(n18188,G36338,n17883);
  nand U19066(n18187,G36306,n17881);
  nand U19067(n18156,G36369,n17843);
  nand U19068(G4474,n18196,n18197,n18198,n18199);
  nor U19069(n18199,n18200,n18201,n18202,n18203);
  nor U19070(n18203,n16934,n17956);
  not U19071(n16934,n16402);
  and U19072(n18202,n16403,n17931);
  xor U19073(n16403,n18171,n18204);
  and U19074(n18204,n18170,n18168);
  nand U19075(n18168,n16402,n17085,n18205);
  nand U19076(n18170,n18206,n18207);
  nand U19077(n18207,n16402,n17085);
  xor U19078(n18206,n17085,n18205);
  nand U19079(n18205,n18208,n18209);
  nand U19080(n18209,n16402,n17937);
  nand U19081(n18208,n16121,n17085);
  nand U19082(n18171,n18210,n18211);
  nand U19083(n18211,n18212,n18213);
  and U19084(n18201,n16401,n17898);
  xor U19085(n16401,n18186,n18214);
  and U19086(n18214,n18185,n18183);
  nand U19087(n18183,n18215,n18216);
  or U19088(n18185,n18215,n18216);
  nand U19089(n18216,n18217,n18218,n17972);
  nand U19090(n18218,n16402,n17973);
  nand U19091(n18217,n17974,n16121);
  xor U19092(n18215,n18219,n17976);
  nand U19093(n18219,n18220,n17916,n18221);
  nand U19094(n18221,n16121,n17973);
  nand U19095(n18220,n16402,n17979);
  nand U19096(n16402,n18222,n18223);
  nand U19097(n18223,n17851,G36175);
  nand U19098(n18222,n18224,n17852);
  nand U19099(n18186,n18225,n18226);
  nand U19100(n18226,n18227,n18228);
  nor U19101(n18200,n16376,n17987);
  not U19102(n16376,n16118);
  nand U19103(n16118,n18229,n18230,n18231,n18232);
  nand U19104(n18232,n18195,n17992);
  not U19105(n18195,n16734);
  xnor U19106(n16734,n18192,G36456);
  nand U19107(n18231,G36369,n17882);
  nand U19108(n18230,G36337,n17883);
  nand U19109(n18229,G36305,n17881);
  nand U19110(n18198,G36368,n17843);
  nand U19111(G4473,n18233,n18234,n18235,n18236);
  nor U19112(n18236,n18237,n18238,n18239,n18240);
  nor U19113(n18240,n16811,n17956);
  not U19114(n16811,n16414);
  and U19115(n18239,n16415,n17931);
  xor U19116(n16415,n18213,n18241);
  and U19117(n18241,n18212,n18210);
  nand U19118(n18210,n16414,n17085,n18242);
  nand U19119(n18212,n18243,n18244);
  nand U19120(n18244,n16414,n17085);
  xor U19121(n18243,n17085,n18242);
  nand U19122(n18242,n18245,n18246);
  nand U19123(n18246,n16414,n17937);
  nand U19124(n18245,n16124,n17085);
  nand U19125(n18213,n18247,n18248);
  nand U19126(n18248,n18249,n18250);
  and U19127(n18238,n16413,n17898);
  xor U19128(n16413,n18228,n18251);
  and U19129(n18251,n18227,n18225);
  nand U19130(n18225,n18252,n18253);
  or U19131(n18227,n18252,n18253);
  nand U19132(n18253,n18254,n18255,n17972);
  nand U19133(n18255,n16414,n17973);
  nand U19134(n18254,n17974,n16124);
  xor U19135(n18252,n18256,n17976);
  nand U19136(n18256,n18257,n17916,n18258);
  nand U19137(n18258,n16124,n17973);
  nand U19138(n18257,n16414,n17979);
  nand U19139(n16414,n18259,n18260);
  nand U19140(n18260,n17851,G36174);
  nand U19141(n18259,n18261,n17852);
  nand U19142(n18228,n18262,n18263);
  nand U19143(n18263,n18264,n18265);
  nor U19144(n18237,n16388,n17987);
  not U19145(n16388,n16121);
  nand U19146(n16121,n18266,n18267,n18268,n18269);
  nand U19147(n18269,n16933,n17992);
  nor U19148(n16933,n18270,n18192);
  and U19149(n18192,G36437,n18271,G36449);
  nor U19150(n18270,G36437,n18272);
  and U19151(n18272,G36449,n18271);
  nand U19152(n18268,G36368,n17882);
  nand U19153(n18267,G36336,n17883);
  nand U19154(n18266,G36304,n17881);
  nand U19155(n18235,G36367,n17843);
  nand U19156(G4472,n18273,n18274,n18275,n18276);
  nor U19157(n18276,n18277,n18278,n18279,n18280);
  nor U19158(n18280,n16913,n17956);
  not U19159(n16913,n16426);
  and U19160(n18279,n16427,n17931);
  xor U19161(n16427,n18250,n18281);
  and U19162(n18281,n18249,n18247);
  nand U19163(n18247,n16426,n17085,n18282);
  nand U19164(n18249,n18283,n18284);
  nand U19165(n18284,n16426,n17085);
  xor U19166(n18283,n17085,n18282);
  nand U19167(n18282,n18285,n18286);
  nand U19168(n18286,n16426,n17937);
  nand U19169(n18285,n16127,n17085);
  nand U19170(n18250,n18287,n18288);
  nand U19171(n18288,n18289,n18290);
  and U19172(n18278,n16425,n17898);
  xor U19173(n16425,n18265,n18291);
  and U19174(n18291,n18264,n18262);
  nand U19175(n18262,n18292,n18293);
  or U19176(n18264,n18292,n18293);
  nand U19177(n18293,n18294,n18295,n17972);
  nand U19178(n18295,n16426,n17973);
  nand U19179(n18294,n17974,n16127);
  xor U19180(n18292,n18296,n17976);
  nand U19181(n18296,n18297,n17916,n18298);
  nand U19182(n18298,n16127,n17973);
  nand U19183(n18297,n16426,n17979);
  nand U19184(n16426,n18299,n18300);
  nand U19185(n18300,n17851,G36173);
  nand U19186(n18299,n18301,n17852);
  nand U19187(n18265,n18302,n18303);
  nand U19188(n18303,n18304,n18305);
  nor U19189(n18277,n16400,n17987);
  not U19190(n16400,n16124);
  nand U19191(n16124,n18306,n18307,n18308,n18309);
  nand U19192(n18309,n16810,n17992);
  xor U19193(n16810,G36449,n18271);
  not U19194(n18271,n18310);
  nand U19195(n18308,G36367,n17882);
  nand U19196(n18307,G36335,n17883);
  nand U19197(n18306,G36303,n17881);
  nand U19198(n18275,G36366,n17843);
  nand U19199(G4471,n18312,n18313,n18314,n18315);
  nor U19200(n18315,n18316,n18317,n18318,n18319);
  nor U19201(n18319,n16769,n17956);
  not U19202(n16769,n16438);
  and U19203(n18318,n16439,n17931);
  xor U19204(n16439,n18290,n18320);
  and U19205(n18320,n18289,n18287);
  nand U19206(n18287,n16438,n17085,n18321);
  nand U19207(n18289,n18322,n18323);
  nand U19208(n18323,n16438,n17085);
  xor U19209(n18322,n17085,n18321);
  nand U19210(n18321,n18324,n18325);
  nand U19211(n18325,n16438,n17937);
  nand U19212(n18324,n16130,n17085);
  nand U19213(n18290,n18326,n18327);
  nand U19214(n18327,n18328,n18329);
  and U19215(n18317,n16437,n17898);
  xor U19216(n16437,n18305,n18330);
  and U19217(n18330,n18304,n18302);
  nand U19218(n18302,n18331,n18332);
  or U19219(n18304,n18331,n18332);
  nand U19220(n18332,n17972,n18333,n18334,n18335);
  nand U19221(n18335,n16438,n17973);
  nand U19222(n18334,n17974,n16130);
  nand U19223(n18333,n16673,n18336);
  not U19224(n17972,n17908);
  nand U19225(n17908,n18337,n18338);
  nand U19226(n18338,n18339,G36365);
  nand U19227(n18337,n18340,G36333);
  xor U19228(n18331,n18341,n17976);
  nand U19229(n18341,n18342,n17916,n18343,n18344);
  nor U19230(n18344,n18345,n18346);
  and U19231(n18346,G36365,n18347);
  and U19232(n18345,G36333,n18348);
  nand U19233(n18343,n16130,n17973);
  nand U19234(n17916,n16673,n18349);
  nand U19235(n18342,n16438,n17979);
  nand U19236(n16438,n18350,n18351,n18352);
  nand U19237(n18352,n16673,n17877);
  nand U19238(n18351,n17851,G36172);
  nand U19239(n18350,n18353,n17852);
  nand U19240(n18305,n18354,n18355);
  nand U19241(n18355,n18356,n18357);
  nor U19242(n18316,n16412,n17987);
  not U19243(n16412,n16127);
  nand U19244(n16127,n18358,n18359,n18360,n18361);
  nand U19245(n18361,n18311,n17992);
  not U19246(n18311,n16912);
  nand U19247(n16912,n18362,n18310);
  nand U19248(n18310,G36439,n18363,G36453);
  nand U19249(n18362,n18364,n18365);
  nand U19250(n18365,G36453,n18363);
  not U19251(n18364,G36439);
  nand U19252(n18360,G36366,n17882);
  nand U19253(n18359,G36334,n17883);
  nand U19254(n18358,G36302,n17881);
  nand U19255(n18314,G36365,n17843);
  nand U19256(G4470,n18367,n18368,n18369,n18370);
  nor U19257(n18370,n18371,n18372,n18373,n18374);
  nor U19258(n18374,n16964,n17956);
  not U19259(n16964,n16450);
  and U19260(n18373,n16451,n17931);
  xor U19261(n16451,n18329,n18375);
  and U19262(n18375,n18328,n18326);
  nand U19263(n18326,n16450,n17085,n18376);
  nand U19264(n18328,n18377,n18378);
  nand U19265(n18378,n16450,n17085);
  xor U19266(n18377,n17085,n18376);
  nand U19267(n18376,n18379,n18380);
  nand U19268(n18380,n16450,n17937);
  nand U19269(n18379,n16133,n17085);
  nand U19270(n18329,n18381,n18382);
  nand U19271(n18382,n18383,n18384);
  and U19272(n18372,n16449,n17898);
  xor U19273(n16449,n18357,n18385);
  and U19274(n18385,n18356,n18354);
  nand U19275(n18354,n18386,n18387);
  or U19276(n18356,n18386,n18387);
  nand U19277(n18387,n18388,n18389,n18390,n18391);
  nor U19278(n18391,n18392,n18393);
  nor U19279(n18393,n18394,n18395);
  nor U19280(n18392,n18396,n18397);
  nand U19281(n18390,n17974,n16133);
  nand U19282(n18389,n16450,n17973);
  nand U19283(n18388,n17701,n18336);
  xor U19284(n18386,n18398,n17976);
  nand U19285(n18398,n18399,n18400,n18401,n18402);
  nor U19286(n18402,n18403,n18404);
  nor U19287(n18404,n18396,n18405);
  not U19288(n18396,G36364);
  nor U19289(n18403,n18394,n18406);
  not U19290(n18394,G36332);
  nand U19291(n18401,n16133,n17973);
  nand U19292(n18400,n16450,n17979);
  nand U19293(n16450,n18407,n18408,n18409);
  nand U19294(n18409,n17701,n17877);
  nand U19295(n18408,n17851,G36171);
  nand U19296(n18407,n18410,n17852);
  nand U19297(n18399,n17701,n18349);
  not U19298(n17701,n17703);
  nand U19299(n17703,n18411,n18412);
  or U19300(n18412,G36236,G36249);
  nand U19301(n18411,G36249,n18413);
  nand U19302(n18357,n18414,n18415);
  nand U19303(n18415,n18416,n18417);
  nor U19304(n18371,n16424,n17987);
  not U19305(n16424,n16130);
  nand U19306(n16130,n18418,n18419,n18420,n18421);
  nand U19307(n18421,n18366,n17992);
  not U19308(n18366,n16768);
  xnor U19309(n16768,n18363,G36453);
  nand U19310(n18420,G36365,n17882);
  nand U19311(n18419,G36333,n17883);
  nand U19312(n18418,G36301,n17881);
  nand U19313(n18369,G36364,n17843);
  nand U19314(n18368,n17929,n16963);
  nand U19315(G4469,n18422,n18423,n18424,n18425);
  nor U19316(n18425,n18426,n18427,n18428,n18429);
  nor U19317(n18429,n16864,n17956);
  not U19318(n16864,n16462);
  and U19319(n18428,n16463,n17931);
  xor U19320(n16463,n18384,n18430);
  and U19321(n18430,n18383,n18381);
  nand U19322(n18381,n16462,n17085,n18431);
  nand U19323(n18383,n18432,n18433);
  nand U19324(n18433,n16462,n17085);
  xor U19325(n18432,n17085,n18431);
  nand U19326(n18431,n18434,n18435);
  nand U19327(n18435,n16462,n17937);
  nand U19328(n18434,n16136,n17085);
  nand U19329(n18384,n18436,n18437);
  nand U19330(n18437,n18438,n18439);
  and U19331(n18427,n16461,n17898);
  xor U19332(n16461,n18417,n18440);
  and U19333(n18440,n18416,n18414);
  nand U19334(n18414,n18441,n18442);
  or U19335(n18416,n18441,n18442);
  nand U19336(n18442,n18443,n18444,n18445,n18446);
  nor U19337(n18446,n18447,n18448);
  nor U19338(n18448,n18449,n18395);
  nor U19339(n18447,n18450,n18397);
  nand U19340(n18445,n17974,n16136);
  nand U19341(n18444,n16462,n17973);
  nand U19342(n18443,n17688,n18336);
  xor U19343(n18441,n18451,n17976);
  nand U19344(n18451,n18452,n18453,n18454,n18455);
  nor U19345(n18455,n18456,n18457);
  nor U19346(n18457,n18450,n18405);
  not U19347(n18450,G36363);
  nor U19348(n18456,n18449,n18406);
  not U19349(n18449,G36331);
  nand U19350(n18454,n16136,n17973);
  nand U19351(n18453,n16462,n17979);
  nand U19352(n16462,n18458,n18459,n18460);
  nand U19353(n18460,n17688,n17877);
  nand U19354(n18459,n17851,G36170);
  nand U19355(n18458,n18461,n17852);
  nand U19356(n18452,n17688,n18349);
  and U19357(n17688,n18462,n18463,n18464);
  nand U19358(n18463,n18465,n18466);
  nand U19359(n18462,G36235,n18467,G36249);
  nand U19360(n18417,n18468,n18469);
  nand U19361(n18469,n18470,n18471);
  nor U19362(n18426,n16436,n17987);
  not U19363(n16436,n16133);
  nand U19364(n16133,n18472,n18473,n18474,n18475);
  nand U19365(n18475,n16963,n17992);
  nor U19366(n16963,n18476,n18363);
  nor U19367(n18363,n17695,n18477,n17683);
  and U19368(n18476,n17695,n18478);
  or U19369(n18478,n17683,n18477);
  not U19370(n17695,G36434);
  nand U19371(n18474,G36364,n17882);
  nand U19372(n18473,G36332,n17883);
  nand U19373(n18472,G36300,n17881);
  nand U19374(n18424,G36363,n17843);
  nand U19375(n18423,n17929,n16863);
  nand U19376(G4468,n18479,n18480,n18481,n18482);
  nor U19377(n18482,n18483,n18484,n18485,n18486);
  nor U19378(n18486,n16843,n17956);
  not U19379(n16843,n16474);
  and U19380(n18485,n16475,n17931);
  xor U19381(n16475,n18439,n18487);
  and U19382(n18487,n18438,n18436);
  nand U19383(n18436,n16474,n17085,n18488);
  nand U19384(n18438,n18489,n18490);
  nand U19385(n18490,n16474,n17085);
  xor U19386(n18489,n17085,n18488);
  nand U19387(n18488,n18491,n18492);
  nand U19388(n18492,n16474,n17937);
  nand U19389(n18491,n16139,n17085);
  nand U19390(n18439,n18493,n18494);
  nand U19391(n18494,n18495,n18496);
  and U19392(n18484,n16473,n17898);
  xor U19393(n16473,n18471,n18497);
  and U19394(n18497,n18470,n18468);
  nand U19395(n18468,n18498,n18499);
  or U19396(n18470,n18498,n18499);
  nand U19397(n18499,n18500,n18501,n18502,n18503);
  nor U19398(n18503,n18504,n18505);
  nor U19399(n18505,n18506,n18395);
  nor U19400(n18504,n18507,n18397);
  nand U19401(n18502,n17974,n16139);
  nand U19402(n18501,n16474,n17973);
  nand U19403(n18500,n17676,n18336);
  xor U19404(n18498,n18508,n17976);
  nand U19405(n18508,n18509,n18510,n18511,n18512);
  nor U19406(n18512,n18513,n18514);
  nor U19407(n18514,n18507,n18405);
  not U19408(n18507,G36362);
  nor U19409(n18513,n18506,n18406);
  not U19410(n18506,G36330);
  nand U19411(n18511,n16139,n17973);
  nand U19412(n18510,n16474,n17979);
  nand U19413(n16474,n18515,n18516,n18517);
  nand U19414(n18517,n17676,n17877);
  nand U19415(n18516,n17851,G36169);
  nand U19416(n18515,n18518,n17852);
  nand U19417(n18509,n17676,n18349);
  and U19418(n17676,n18519,n18520);
  or U19419(n18520,G36234,G36249);
  nand U19420(n18519,G36249,n18521);
  nand U19421(n18471,n18522,n18523);
  nand U19422(n18523,n18524,n18525);
  nor U19423(n18483,n16448,n17987);
  not U19424(n16448,n16136);
  nand U19425(n16136,n18526,n18527,n18528,n18529);
  nand U19426(n18529,n16863,n17992);
  xor U19427(n16863,n17683,n18477);
  not U19428(n17683,G36444);
  nand U19429(n18528,G36363,n17882);
  nand U19430(n18527,G36331,n17883);
  nand U19431(n18526,G36299,n17881);
  nand U19432(n18481,G36362,n17843);
  nand U19433(n18480,n17929,n18530);
  nand U19434(n18479,n17993,n16142);
  nand U19435(G4467,n18531,n18532,n18533,n18534);
  nor U19436(n18534,n18535,n18536,n18537,n18538);
  nor U19437(n18538,n17011,n17956);
  not U19438(n17011,n16486);
  and U19439(n18537,n16487,n17931);
  xor U19440(n16487,n18496,n18539);
  and U19441(n18539,n18495,n18493);
  nand U19442(n18493,n16486,n17085,n18540);
  nand U19443(n18495,n18541,n18542);
  nand U19444(n18542,n16486,n17085);
  xor U19445(n18541,n17085,n18540);
  nand U19446(n18540,n18543,n18544);
  nand U19447(n18544,n17085,n16142);
  nand U19448(n18543,n16486,n17937);
  nand U19449(n18496,n18545,n18546);
  nand U19450(n18546,n18547,n18548);
  and U19451(n18536,n16485,n17898);
  xor U19452(n16485,n18525,n18549);
  and U19453(n18549,n18524,n18522);
  nand U19454(n18522,n18550,n18551);
  or U19455(n18524,n18550,n18551);
  nand U19456(n18551,n18552,n18553,n18554,n18555);
  nor U19457(n18555,n18556,n18557);
  nor U19458(n18557,n17819,n18395);
  nor U19459(n18556,n17820,n18397);
  nand U19460(n18554,n17974,n16142);
  nand U19461(n18553,n16486,n17973);
  nand U19462(n18552,n17663,n18336);
  xor U19463(n18550,n18558,n17976);
  nand U19464(n18558,n18559,n18560,n18561,n18562);
  nor U19465(n18562,n18563,n18564);
  nor U19466(n18564,n17820,n18405);
  not U19467(n17820,G36361);
  nor U19468(n18563,n17819,n18406);
  not U19469(n17819,G36329);
  nand U19470(n18561,n16142,n17973);
  nand U19471(n18560,n16486,n17979);
  nand U19472(n16486,n18565,n18566,n18567);
  nand U19473(n18567,n17663,n17877);
  nand U19474(n18566,n17851,G36168);
  nand U19475(n18565,n18568,n17852);
  nand U19476(n18559,n17663,n18349);
  not U19477(n17663,n17816);
  nand U19478(n17816,n18569,n18570,n18571);
  nand U19479(n18570,n18572,n18466);
  nand U19480(n18569,G36233,n18573,G36249);
  nand U19481(n18525,n18574,n18575);
  nand U19482(n18575,n18576,n18577);
  nor U19483(n18535,n16460,n17987);
  not U19484(n16460,n16139);
  nand U19485(n16139,n18578,n18579,n18580,n18581);
  nand U19486(n18581,n18530,n17992);
  not U19487(n18530,n16842);
  nand U19488(n16842,n18582,n18477);
  nand U19489(n18477,G36431,n18583,G36446);
  nand U19490(n18582,n17670,n18584);
  nand U19491(n18584,G36431,n18583);
  not U19492(n18583,n18585);
  not U19493(n17670,G36446);
  nand U19494(n18580,G36362,n17882);
  nand U19495(n18579,G36330,n17883);
  nand U19496(n18578,G36298,n17881);
  nand U19497(n18533,G36361,n17843);
  nand U19498(n18532,n17929,n18586);
  nand U19499(n18531,n17993,n16145);
  nand U19500(G4466,n18587,n18588,n18589,n18590);
  nor U19501(n18590,n18591,n18592,n18593,n18594);
  nor U19502(n18594,n16725,n17956);
  not U19503(n16725,n16498);
  and U19504(n18593,n16499,n17931);
  xor U19505(n16499,n18548,n18595);
  and U19506(n18595,n18545,n18547);
  nand U19507(n18547,n18596,n18597);
  nand U19508(n18597,n16498,n17085);
  xor U19509(n18596,n17085,n18598);
  nand U19510(n18545,n16498,n17085,n18598);
  nand U19511(n18598,n18599,n18600);
  nand U19512(n18600,n16498,n17937);
  nand U19513(n18599,n16145,n17085);
  nand U19514(n18548,n18601,n18602);
  nand U19515(n18602,n18603,n18604);
  and U19516(n18592,n16497,n17898);
  xor U19517(n16497,n18577,n18605);
  and U19518(n18605,n18574,n18576);
  or U19519(n18576,n18606,n18607);
  nand U19520(n18574,n18606,n18607);
  nand U19521(n18607,n18608,n18609,n18610,n18611);
  nor U19522(n18611,n18612,n18613);
  nor U19523(n18613,n18614,n18395);
  nor U19524(n18612,n18615,n18397);
  nand U19525(n18610,n17974,n16145);
  nand U19526(n18609,n16498,n17973);
  nand U19527(n18608,n17650,n18336);
  xor U19528(n18606,n18616,n17976);
  nand U19529(n18616,n18617,n18618,n18619,n18620);
  nor U19530(n18620,n18621,n18622);
  nor U19531(n18622,n18615,n18405);
  not U19532(n18615,G36360);
  nor U19533(n18621,n18614,n18406);
  not U19534(n18614,G36328);
  nand U19535(n18619,n16145,n17973);
  nand U19536(n18618,n16498,n17979);
  nand U19537(n16498,n18623,n18624,n18625);
  nand U19538(n18625,n17650,n17877);
  nand U19539(n18624,n17851,G36167);
  nand U19540(n18623,n17852,n18626);
  nand U19541(n18617,n17650,n18349);
  and U19542(n17650,n18627,n18628);
  or U19543(n18628,G36232,G36249);
  nand U19544(n18627,G36249,n18629);
  nand U19545(n18577,n18630,n18631);
  nand U19546(n18631,n18632,n18633);
  nor U19547(n18591,n16472,n17987);
  not U19548(n16472,n16142);
  nand U19549(n16142,n18634,n18635,n18636,n18637);
  nand U19550(n18637,n18586,n17992);
  not U19551(n18586,n16997);
  xor U19552(n16997,n18585,G36431);
  nand U19553(n18636,G36361,n17882);
  nand U19554(n18635,G36329,n17883);
  nand U19555(n18634,G36297,n17881);
  nand U19556(n18589,G36360,n17843);
  nand U19557(n18588,n17929,n18638);
  nand U19558(n18587,n17993,n16148);
  nand U19559(G4465,n18639,n18640,n18641,n18642);
  nor U19560(n18642,n18643,n18644,n18645,n18646);
  nor U19561(n18646,n16923,n17956);
  not U19562(n16923,n16510);
  and U19563(n18645,n16511,n17931);
  xor U19564(n16511,n18604,n18647);
  and U19565(n18647,n18603,n18601);
  nand U19566(n18601,n16510,n17085,n18648);
  nand U19567(n18603,n18649,n18650);
  nand U19568(n18650,n16510,n17085);
  xor U19569(n18649,n17085,n18648);
  nand U19570(n18648,n18651,n18652);
  nand U19571(n18652,n16510,n17937);
  nand U19572(n18651,n16148,n17085);
  nand U19573(n18604,n18653,n18654);
  nand U19574(n18654,n18655,n18656);
  and U19575(n18644,n16509,n17898);
  xor U19576(n16509,n18633,n18657);
  and U19577(n18657,n18632,n18630);
  nand U19578(n18630,n18658,n18659);
  or U19579(n18632,n18658,n18659);
  nand U19580(n18659,n18660,n18661,n18662,n18663);
  nor U19581(n18663,n18664,n18665);
  nor U19582(n18665,n18666,n18395);
  nor U19583(n18664,n18667,n18397);
  nand U19584(n18662,n17974,n16148);
  nand U19585(n18661,n16510,n17973);
  nand U19586(n18660,n17637,n18336);
  xor U19587(n18658,n18668,n17976);
  nand U19588(n18668,n18669,n18670,n18671,n18672);
  nor U19589(n18672,n18673,n18674);
  nor U19590(n18674,n18667,n18405);
  not U19591(n18667,G36359);
  nor U19592(n18673,n18666,n18406);
  not U19593(n18666,G36327);
  nand U19594(n18671,n16148,n17973);
  nand U19595(n18670,n16510,n17979);
  nand U19596(n16510,n18675,n18676,n18677);
  nand U19597(n18677,n17637,n17877);
  nand U19598(n18676,n17851,G36166);
  nand U19599(n18675,n18678,n17852);
  nand U19600(n18669,n17637,n18349);
  not U19601(n17637,n17745);
  nand U19602(n17745,n18679,n18680,n18681);
  nand U19603(n18680,n18682,n18466);
  nand U19604(n18679,G36231,n18683,G36249);
  nand U19605(n18633,n18684,n18685);
  nand U19606(n18685,n18686,n18687);
  nor U19607(n18643,n16484,n17987);
  not U19608(n16484,n16145);
  nand U19609(n16145,n18688,n18689,n18690,n18691);
  nand U19610(n18691,n18638,n17992);
  not U19611(n18638,n16724);
  nand U19612(n16724,n18692,n18585);
  nand U19613(n18585,G36438,n18693,G36457);
  nand U19614(n18692,n17644,n18694);
  nand U19615(n18694,G36438,n18693);
  not U19616(n17644,G36457);
  nand U19617(n18690,G36360,n17882);
  nand U19618(n18689,G36328,n17883);
  nand U19619(n18688,G36296,n17881);
  nand U19620(n18641,G36359,n17843);
  nand U19621(n18640,n17929,n18695);
  nand U19622(n18639,n17993,n16151);
  nand U19623(G4464,n18696,n18697,n18698,n18699);
  nor U19624(n18699,n18700,n18701,n18702,n18703);
  nor U19625(n18703,n16822,n17956);
  and U19626(n18702,n16523,n17931);
  xor U19627(n16523,n18656,n18704);
  and U19628(n18704,n18655,n18653);
  nand U19629(n18653,n16522,n17085,n18705);
  nand U19630(n18655,n18706,n18707);
  nand U19631(n18707,n16522,n17085);
  xor U19632(n18706,n17085,n18705);
  nand U19633(n18705,n18708,n18709);
  nand U19634(n18709,n16522,n17937);
  nand U19635(n18708,n16151,n17085);
  nand U19636(n18656,n18710,n18711);
  nand U19637(n18711,n18712,n18713);
  and U19638(n18701,n16521,n17898);
  xor U19639(n16521,n18687,n18714);
  and U19640(n18714,n18686,n18684);
  nand U19641(n18684,n18715,n18716);
  or U19642(n18686,n18715,n18716);
  nand U19643(n18716,n18717,n18718,n18719,n18720);
  nor U19644(n18720,n18721,n18722);
  and U19645(n18722,G36326,n18340);
  and U19646(n18721,G36358,n18339);
  nand U19647(n18719,n17974,n16151);
  nand U19648(n18718,n16522,n17973);
  nand U19649(n18717,n17625,n18336);
  xor U19650(n18715,n18723,n17976);
  nand U19651(n18723,n18724,n18725,n18726,n18727);
  nand U19652(n18727,n16151,n17973);
  nor U19653(n18726,n18728,n18729);
  nor U19654(n18729,n18730,n17624);
  nor U19655(n18728,n18731,n16822);
  not U19656(n16822,n16522);
  nand U19657(n16522,n18732,n18733,n18734);
  nand U19658(n18734,n17625,n17877);
  not U19659(n17625,n17624);
  nand U19660(n17624,n18735,n18736);
  or U19661(n18736,G36230,G36249);
  nand U19662(n18735,G36249,n18737);
  nand U19663(n18733,n17851,G36165);
  nand U19664(n18732,n18738,n17852);
  nand U19665(n18725,n18348,G36326);
  nand U19666(n18724,n18347,G36358);
  nand U19667(n18687,n18739,n18740);
  nand U19668(n18740,n18741,n18742);
  nor U19669(n18700,n16496,n17987);
  not U19670(n16496,n16148);
  nand U19671(n16148,n18743,n18744,n18745,n18746);
  nand U19672(n18746,n18695,n17992);
  not U19673(n18695,n16922);
  xnor U19674(n16922,G36438,n18693);
  nand U19675(n18745,G36359,n17882);
  nand U19676(n18744,G36327,n17883);
  nand U19677(n18743,G36295,n17881);
  nand U19678(n18698,G36358,n17843);
  nand U19679(n18697,n17929,n16821);
  nand U19680(n18696,n17993,n16154);
  nand U19681(G4463,n18747,n18748,n18749,n18750);
  nor U19682(n18750,n18751,n18752,n18753,n18754);
  nor U19683(n18754,n16944,n17956);
  and U19684(n18753,n16535,n17931);
  xor U19685(n16535,n18713,n18755);
  and U19686(n18755,n18712,n18710);
  nand U19687(n18710,n16534,n17085,n18756);
  nand U19688(n18712,n18757,n18758);
  nand U19689(n18758,n16534,n17085);
  xor U19690(n18757,n17085,n18756);
  nand U19691(n18756,n18759,n18760);
  nand U19692(n18760,n16534,n17937);
  nand U19693(n18759,n16154,n17085);
  nand U19694(n18713,n18761,n18762);
  nand U19695(n18762,n18763,n18764);
  and U19696(n18752,n16533,n17898);
  xor U19697(n16533,n18742,n18765);
  and U19698(n18765,n18741,n18739);
  nand U19699(n18739,n18766,n18767);
  or U19700(n18741,n18766,n18767);
  nand U19701(n18767,n18768,n18769,n18770,n18771);
  nand U19702(n18771,n17974,n16154);
  nor U19703(n18770,n18772,n18773);
  nor U19704(n18773,n18774,n17606);
  nor U19705(n18772,n18775,n16944);
  nand U19706(n18769,n18339,G36357);
  nand U19707(n18768,n18340,G36325);
  xor U19708(n18766,n18776,n17976);
  nand U19709(n18776,n18777,n18778,n18779,n18780);
  nand U19710(n18780,n16154,n17973);
  nor U19711(n18779,n18781,n18782);
  nor U19712(n18782,n18730,n17606);
  nor U19713(n18781,n18731,n16944);
  not U19714(n16944,n16534);
  nand U19715(n16534,n18783,n18784,n18785);
  nand U19716(n18785,n17611,n17877);
  not U19717(n17611,n17606);
  nand U19718(n17606,n18786,n18787,n18788);
  nand U19719(n18787,n18789,n18466);
  nand U19720(n18786,G36229,n18790,G36249);
  nand U19721(n18784,n17851,G36164);
  nand U19722(n18783,n18791,n17852);
  nand U19723(n18778,n18348,G36325);
  nand U19724(n18777,n18347,G36357);
  nand U19725(n18742,n18792,n18793);
  nand U19726(n18793,n18794,n18795);
  nor U19727(n18751,n16508,n17987);
  not U19728(n16508,n16151);
  nand U19729(n16151,n18796,n18797,n18798,n18799);
  nand U19730(n18799,n16821,n17992);
  nor U19731(n16821,n18800,n18693);
  nor U19732(n18693,n17618,n18801);
  and U19733(n18800,n17618,n18801);
  not U19734(n17618,G36448);
  nand U19735(n18798,G36358,n17882);
  nand U19736(n18797,G36326,n17883);
  nand U19737(n18796,G36294,n17881);
  nand U19738(n18749,G36357,n17843);
  nand U19739(n18748,n17929,n18802);
  nand U19740(n18747,n17993,n16157);
  nand U19741(G4462,n18803,n18804,n18805,n18806);
  nor U19742(n18806,n18807,n18808,n18809,n18810);
  nor U19743(n18810,n16745,n17956);
  and U19744(n18809,n16547,n17931);
  xor U19745(n16547,n18763,n18811);
  and U19746(n18811,n18761,n18764);
  nand U19747(n18764,n18812,n18813);
  nand U19748(n18813,n16546,n17085);
  xor U19749(n18812,n17085,n18814);
  nand U19750(n18761,n16546,n17085,n18814);
  nand U19751(n18814,n18815,n18816);
  nand U19752(n18816,n16546,n17937);
  nand U19753(n18815,n16157,n17085);
  nand U19754(n18763,n18817,n18818);
  nand U19755(n18818,n18819,n18820);
  and U19756(n18808,n16545,n17898);
  xor U19757(n16545,n18794,n18821);
  and U19758(n18821,n18792,n18795);
  or U19759(n18795,n18822,n18823);
  nand U19760(n18792,n18822,n18823);
  nand U19761(n18823,n18824,n18825,n18826,n18827);
  nand U19762(n18827,n17974,n16157);
  nor U19763(n18826,n18828,n18829);
  nor U19764(n18829,n18774,n17755);
  nor U19765(n18828,n18775,n16745);
  nand U19766(n18825,n18339,G36356);
  nand U19767(n18824,n18340,G36324);
  xor U19768(n18822,n18830,n17976);
  nand U19769(n18830,n18831,n18832,n18833,n18834);
  nand U19770(n18834,n16157,n17973);
  nor U19771(n18833,n18835,n18836);
  nor U19772(n18836,n18730,n17755);
  nor U19773(n18835,n18731,n16745);
  not U19774(n16745,n16546);
  nand U19775(n16546,n18837,n18838,n18839);
  nand U19776(n18839,n17593,n17877);
  not U19777(n17593,n17755);
  nand U19778(n17755,n18840,n18841);
  or U19779(n18841,G36228,G36249);
  nand U19780(n18840,G36249,n18842);
  nand U19781(n18838,n17851,G36163);
  nand U19782(n18837,n17852,n18843);
  nand U19783(n18832,n18348,G36324);
  nand U19784(n18831,n18347,G36356);
  nand U19785(n18794,n18844,n18845);
  nand U19786(n18845,n18846,n18847);
  nor U19787(n18807,n16520,n17987);
  not U19788(n16520,n16154);
  nand U19789(n16154,n18848,n18849,n18850,n18851);
  nand U19790(n18851,n18802,n17992);
  not U19791(n18802,n16943);
  nand U19792(n16943,n18801,n18852);
  nand U19793(n18852,n18853,n17600);
  not U19794(n17600,G36436);
  nand U19795(n18853,G36455,n18854);
  nand U19796(n18801,G36436,n18854,G36455);
  nand U19797(n18850,G36357,n17882);
  nand U19798(n18849,G36325,n17883);
  nand U19799(n18848,G36293,n17881);
  nand U19800(n18805,G36356,n17843);
  nand U19801(n18804,n17929,n18855);
  nand U19802(n18803,n17993,n16160);
  nand U19803(G4461,n18856,n18857,n18858,n18859);
  nor U19804(n18859,n18860,n18861,n18862,n18863);
  nor U19805(n18863,n16895,n17956);
  and U19806(n18862,n16559,n17931);
  xor U19807(n16559,n18820,n18864);
  and U19808(n18864,n18819,n18817);
  nand U19809(n18817,n16558,n17085,n18865);
  nand U19810(n18819,n18866,n18867);
  nand U19811(n18867,n16558,n17085);
  xor U19812(n18866,n17085,n18865);
  nand U19813(n18865,n18868,n18869);
  nand U19814(n18869,n16558,n17937);
  nand U19815(n18868,n16160,n17085);
  nand U19816(n18820,n18870,n18871);
  nand U19817(n18871,n18872,n18873);
  and U19818(n18861,n16557,n17898);
  xor U19819(n16557,n18847,n18874);
  and U19820(n18874,n18846,n18844);
  nand U19821(n18844,n18875,n18876);
  or U19822(n18846,n18875,n18876);
  nand U19823(n18876,n18877,n18878,n18879,n18880);
  nand U19824(n18880,n17974,n16160);
  nor U19825(n18879,n18881,n18882);
  nor U19826(n18882,n18774,n17578);
  nor U19827(n18881,n18775,n16895);
  nand U19828(n18878,n18339,G36355);
  nand U19829(n18877,n18340,G36323);
  xor U19830(n18875,n18883,n17976);
  nand U19831(n18883,n18884,n18885,n18886,n18887);
  nand U19832(n18887,n16160,n17973);
  nor U19833(n18886,n18888,n18889);
  nor U19834(n18889,n18730,n17578);
  nor U19835(n18888,n18731,n16895);
  not U19836(n16895,n16558);
  nand U19837(n16558,n18890,n18891,n18892);
  nand U19838(n18892,n17580,n17877);
  not U19839(n17580,n17578);
  nand U19840(n17578,n18893,n18894,n18895);
  nand U19841(n18894,n18896,n18466);
  nand U19842(n18893,G36227,n18897,G36249);
  nand U19843(n18891,n17851,G36162);
  nand U19844(n18890,n18898,n17852);
  nand U19845(n18885,n18348,G36323);
  nand U19846(n18884,n18347,G36355);
  nand U19847(n18847,n18899,n18900);
  nand U19848(n18900,n18901,n18902);
  nor U19849(n18860,n16532,n17987);
  not U19850(n16532,n16157);
  nand U19851(n16157,n18903,n18904,n18905,n18906);
  nand U19852(n18906,n18855,n17992);
  not U19853(n18855,n16744);
  xnor U19854(n16744,G36455,n18854);
  nand U19855(n18905,G36356,n17882);
  nand U19856(n18904,G36324,n17883);
  nand U19857(n18903,G36292,n17881);
  nand U19858(n18858,G36355,n17843);
  nand U19859(n18857,n17929,n16894);
  nand U19860(n18856,n17993,n16163);
  nand U19861(G4460,n18907,n18908,n18909,n18910);
  nor U19862(n18910,n18911,n18912,n18913,n18914);
  nor U19863(n18914,n16790,n17956);
  and U19864(n18913,n16571,n17931);
  xor U19865(n16571,n18873,n18915);
  and U19866(n18915,n18870,n18872);
  nand U19867(n18872,n18916,n18917);
  nand U19868(n18917,n16570,n17085);
  or U19869(n18870,n18916,n16790);
  and U19870(n18916,n18918,n18919);
  nand U19871(n18919,n16790,n17937);
  nand U19872(n18918,n16163,n17085);
  nand U19873(n18873,n18920,n18921);
  nand U19874(n18921,n18922,n18923);
  and U19875(n18912,n16569,n17898);
  xor U19876(n16569,n18902,n18924);
  and U19877(n18924,n18901,n18899);
  nand U19878(n18899,n18925,n18926);
  or U19879(n18901,n18925,n18926);
  nand U19880(n18926,n18927,n18928,n18929,n18930);
  nand U19881(n18930,n17974,n16163);
  nor U19882(n18929,n18931,n18932);
  nor U19883(n18932,n18774,n17565);
  nor U19884(n18931,n18775,n16790);
  nand U19885(n18928,n18339,G36354);
  nand U19886(n18927,n18340,G36322);
  xor U19887(n18925,n18933,n17976);
  nand U19888(n18933,n18934,n18935,n18936,n18937);
  nand U19889(n18937,n16163,n17973);
  nor U19890(n18936,n18938,n18939);
  nor U19891(n18939,n18730,n17565);
  nor U19892(n18938,n18731,n16790);
  not U19893(n16790,n16570);
  nand U19894(n16570,n18940,n18941,n18942);
  nand U19895(n18942,n17566,n17877);
  not U19896(n17566,n17565);
  nand U19897(n17565,n18943,n18944);
  or U19898(n18944,G36226,G36249);
  nand U19899(n18943,G36249,n18945);
  nand U19900(n18941,n17851,G36161);
  nand U19901(n18940,n18946,n17852);
  nand U19902(n18935,n18348,G36322);
  nand U19903(n18934,n18347,G36354);
  nand U19904(n18902,n18947,n18948);
  nand U19905(n18948,n18949,n18950);
  nor U19906(n18911,n16544,n17987);
  not U19907(n16544,n16160);
  nand U19908(n16160,n18951,n18952,n18953,n18954);
  nand U19909(n18954,n16894,n17992);
  nor U19910(n16894,n18854,n18955);
  and U19911(n18955,n18956,n17573);
  nor U19912(n18854,n17573,n18956);
  nand U19913(n18956,G36451,n18957);
  not U19914(n17573,G36441);
  nand U19915(n18953,G36355,n17882);
  nand U19916(n18952,G36323,n17883);
  nand U19917(n18951,G36291,n17881);
  nand U19918(n18909,G36354,n17843);
  nand U19919(n18908,n17929,n18958);
  nand U19920(n18907,n17993,n16166);
  nand U19921(G4459,n18959,n18960,n18961,n18962);
  nor U19922(n18962,n18963,n18964,n18965,n18966);
  nor U19923(n18966,n16702,n17956);
  and U19924(n18965,n16583,n17931);
  xor U19925(n16583,n18923,n18967);
  and U19926(n18967,n18922,n18920);
  nand U19927(n18920,n16582,n17085,n18968);
  nand U19928(n18922,n18969,n18970);
  nand U19929(n18970,n16582,n17085);
  xor U19930(n18969,n17085,n18968);
  nand U19931(n18968,n18971,n18972);
  nand U19932(n18972,n16582,n17937);
  nand U19933(n18971,n16166,n17085);
  nand U19934(n18923,n18973,n18974);
  nand U19935(n18974,n18975,n18976);
  and U19936(n18964,n16581,n17898);
  xor U19937(n16581,n18949,n18977);
  and U19938(n18977,n18947,n18950);
  or U19939(n18950,n18978,n18979);
  nand U19940(n18947,n18978,n18979);
  nand U19941(n18979,n18980,n18981,n18982,n18983);
  nand U19942(n18983,n17974,n16166);
  nor U19943(n18982,n18984,n18985);
  nor U19944(n18985,n18774,n18986);
  nor U19945(n18984,n18775,n16702);
  nand U19946(n18981,n18339,G36353);
  nand U19947(n18980,n18340,G36321);
  xor U19948(n18978,n18987,n17976);
  nand U19949(n18987,n18988,n18989,n18990,n18991);
  nand U19950(n18991,n16166,n17973);
  nor U19951(n18990,n18992,n18993);
  nor U19952(n18993,n18730,n18986);
  nor U19953(n18992,n18731,n16702);
  not U19954(n16702,n16582);
  nand U19955(n16582,n18994,n18995,n18996);
  nand U19956(n18996,n17553,n17877);
  not U19957(n17553,n18986);
  nand U19958(n18986,n18997,n18998,n18999);
  nand U19959(n18998,n19000,n18466);
  nand U19960(n18997,G36225,n19001,G36249);
  nand U19961(n18995,n17851,G36160);
  nand U19962(n18994,n19002,n17852);
  nand U19963(n18989,n18348,G36321);
  nand U19964(n18988,n18347,G36353);
  nand U19965(n18949,n19003,n19004);
  nand U19966(n19004,n19005,n19006);
  nor U19967(n18963,n16556,n17987);
  not U19968(n16556,n16163);
  nand U19969(n16163,n19007,n19008,n19009,n19010);
  nand U19970(n19010,n18958,n17992);
  not U19971(n18958,n16789);
  xnor U19972(n16789,G36451,n18957);
  nor U19973(n18957,n17547,n19011);
  not U19974(n17547,G36459);
  nand U19975(n19009,G36354,n17882);
  nand U19976(n19008,G36322,n17883);
  nand U19977(n19007,G36290,n17881);
  nand U19978(n18961,G36353,n17843);
  nand U19979(n18960,n17929,n19012);
  nand U19980(n18959,n17993,n16169);
  nand U19981(G4458,n19013,n19014,n19015,n19016);
  nor U19982(n19016,n19017,n19018,n19019,n19020);
  nor U19983(n19020,n16974,n17956);
  and U19984(n19019,n16595,n17931);
  xor U19985(n16595,n18975,n19021);
  and U19986(n19021,n18973,n18976);
  nand U19987(n18976,n19022,n19023);
  nand U19988(n19023,n16594,n17085);
  xor U19989(n19022,n17085,n19024);
  nand U19990(n18973,n16594,n17085,n19024);
  nand U19991(n19024,n19025,n19026);
  nand U19992(n19026,n16594,n17937);
  nand U19993(n19025,n16169,n17085);
  nand U19994(n18975,n19027,n19028);
  nand U19995(n19028,n19029,n19030);
  and U19996(n19018,n16593,n17898);
  xor U19997(n16593,n19005,n19031);
  and U19998(n19031,n19003,n19006);
  or U19999(n19006,n19032,n19033);
  nand U20000(n19003,n19032,n19033);
  nand U20001(n19033,n19034,n19035,n19036,n19037);
  nor U20002(n19036,n19038,n19039);
  nor U20003(n19039,n18774,n17799);
  nor U20004(n19038,n18775,n16974);
  nand U20005(n19035,n18339,G36352);
  nand U20006(n19034,n18340,G36320);
  xor U20007(n19032,n19040,n17976);
  nand U20008(n19040,n19041,n19042,n19043,n19044);
  nand U20009(n19044,n16169,n17973);
  nor U20010(n19043,n19045,n19046);
  nor U20011(n19046,n18730,n17799);
  nor U20012(n19045,n18731,n16974);
  not U20013(n16974,n16594);
  nand U20014(n16594,n19047,n19048,n19049);
  nand U20015(n19049,n17540,n17877);
  not U20016(n17540,n17799);
  nand U20017(n17799,n19050,n19051);
  or U20018(n19051,G36224,G36249);
  nand U20019(n19050,G36249,n19052);
  nand U20020(n19048,n17851,G36159);
  nand U20021(n19047,n19053,n17852);
  nand U20022(n19042,n18348,G36320);
  nand U20023(n19041,n18347,G36352);
  nand U20024(n19005,n19054,n19055);
  nand U20025(n19055,n19056,n19057);
  nor U20026(n19017,n16568,n17987);
  not U20027(n16568,n16166);
  nand U20028(n16166,n19058,n19059,n19060,n19061);
  nand U20029(n19061,n19012,n17992);
  not U20030(n19012,n16701);
  xor U20031(n16701,n19011,G36459);
  nand U20032(n19060,G36353,n17882);
  nand U20033(n19059,G36321,n17883);
  nand U20034(n19058,G36289,n17881);
  nand U20035(n19015,G36352,n17843);
  nand U20036(n19014,n17929,n19062);
  nand U20037(n19013,n17993,n16172);
  nand U20038(G4457,n19063,n19064,n19065,n19066);
  nor U20039(n19066,n19067,n19068,n19069,n19070);
  nor U20040(n19070,n16853,n17956);
  and U20041(n19069,n16607,n17931);
  xor U20042(n16607,n19030,n19071);
  and U20043(n19071,n19029,n19027);
  nand U20044(n19027,n16606,n17085,n19072);
  nand U20045(n19029,n19073,n19074);
  nand U20046(n19074,n16606,n17085);
  xor U20047(n19073,n17085,n19072);
  nand U20048(n19072,n19075,n19076);
  nand U20049(n19076,n16606,n17937);
  nand U20050(n19075,n16172,n17085);
  nand U20051(n19030,n19077,n19078);
  nand U20052(n19078,n19079,n19080);
  and U20053(n19068,n16605,n17898);
  xor U20054(n16605,n19057,n19081);
  and U20055(n19081,n19056,n19054);
  nand U20056(n19054,n19082,n19083);
  or U20057(n19056,n19082,n19083);
  nand U20058(n19083,n19084,n19085,n19086,n19087);
  nor U20059(n19086,n19088,n19089);
  nor U20060(n19089,n18774,n17794);
  nor U20061(n19088,n18775,n16853);
  nand U20062(n19085,n18339,G36351);
  nand U20063(n19084,n18340,G36319);
  xor U20064(n19082,n19090,n17976);
  nand U20065(n19090,n19091,n19092,n19093,n19094);
  nand U20066(n19094,n16172,n17973);
  nor U20067(n19093,n19095,n19096);
  nor U20068(n19096,n18730,n17794);
  nor U20069(n19095,n18731,n16853);
  not U20070(n16853,n16606);
  nand U20071(n16606,n19097,n19098,n19099);
  nand U20072(n19099,n17527,n17877);
  not U20073(n17527,n17794);
  nand U20074(n17794,n19100,n19101,n19102);
  nand U20075(n19101,n19103,n18466);
  nand U20076(n19100,G36223,n19104,G36249);
  nand U20077(n19098,n17851,G36158);
  nand U20078(n19097,n19105,n17852);
  nand U20079(n19092,n18348,G36319);
  nand U20080(n19091,n18347,G36351);
  nand U20081(n19057,n19106,n19107);
  nand U20082(n19107,n19108,n19109);
  nor U20083(n19067,n16580,n17987);
  not U20084(n16580,n16169);
  nand U20085(n16169,n19110,n19111,n19112,n19113);
  nand U20086(n19113,n19062,n17992);
  not U20087(n19062,n16973);
  nand U20088(n16973,n19011,n19114);
  nand U20089(n19114,n19115,n17534);
  or U20090(n19011,n17534,n19115);
  nand U20091(n19115,G36445,n19116);
  not U20092(n17534,G36433);
  nand U20093(n19112,G36352,n17882);
  nand U20094(n19111,G36320,n17883);
  nand U20095(n19110,G36288,n17881);
  nand U20096(n19065,G36351,n17843);
  nand U20097(n19064,n17929,n19117);
  nand U20098(n19063,n17993,n16175);
  nand U20099(G4456,n19118,n19119,n19120,n19121);
  nor U20100(n19121,n19122,n19123,n19124,n19125);
  and U20101(n19125,n16619,n17931);
  xor U20102(n16619,n19080,n19126);
  and U20103(n19126,n19077,n19079);
  nand U20104(n19079,n19127,n19128);
  nand U20105(n19128,n16618,n17085);
  or U20106(n19077,n19127,n16883);
  and U20107(n19127,n19129,n19130);
  nand U20108(n19130,n16883,n17937);
  nand U20109(n19129,n16175,n17085);
  nand U20110(n19080,n19131,n19132);
  nand U20111(n19132,n19133,n19134);
  and U20112(n19124,n16617,n17898);
  xor U20113(n16617,n19109,n19135);
  and U20114(n19135,n19108,n19106);
  nand U20115(n19106,n19136,n19137);
  or U20116(n19108,n19136,n19137);
  nand U20117(n19137,n19138,n19139,n19140,n19141);
  nand U20118(n19141,n17974,n16175);
  nor U20119(n19140,n19142,n19143);
  nor U20120(n19143,n18774,n17770);
  nor U20121(n19142,n18775,n16883);
  nand U20122(n19139,n18339,G36350);
  nand U20123(n19138,n18340,G36318);
  xor U20124(n19136,n19144,n17976);
  nand U20125(n19144,n19145,n19146,n19147,n19148);
  nand U20126(n19148,n16175,n17973);
  nor U20127(n19147,n19149,n19150);
  nor U20128(n19150,n18730,n17770);
  nor U20129(n19149,n18731,n16883);
  not U20130(n16883,n16618);
  nand U20131(n19146,n18348,G36318);
  nand U20132(n19145,n18347,G36350);
  nand U20133(n19109,n19151,n19152);
  nand U20134(n19152,n19153,n19154);
  nor U20135(n19123,n16592,n17987);
  not U20136(n16592,n16172);
  nand U20137(n16172,n19155,n19156,n19157,n19158);
  nand U20138(n19158,n19117,n17992);
  not U20139(n19117,n16852);
  xnor U20140(n16852,n19116,G36445);
  nand U20141(n19157,G36351,n17882);
  nand U20142(n19156,G36319,n17883);
  nand U20143(n19155,G36287,n17881);
  nor U20144(n19122,n16884,n19159);
  not U20145(n16884,n19160);
  nand U20146(n19120,G36350,n17843);
  nand U20147(n19119,n17842,n16618);
  nand U20148(n16618,n19161,n19162,n19163);
  nand U20149(n19163,n17515,n17877);
  not U20150(n17515,n17770);
  nand U20151(n17770,n19164,n19165);
  or U20152(n19165,G36222,G36249);
  nand U20153(n19164,G36249,n19166);
  nand U20154(n19162,n17851,G36157);
  nand U20155(n19161,n17852,n19167);
  not U20156(n17842,n17956);
  nand U20157(n19118,n17993,n16178);
  nand U20158(G4455,n19168,n19169,n19170,n19171);
  nor U20159(n19171,n19172,n19173,n19174,n19175);
  nor U20160(n19175,n16759,n17956);
  nor U20161(n19174,n16754,n19176);
  not U20162(n16754,n16631);
  xor U20163(n16631,n19134,n19177);
  and U20164(n19177,n19133,n19131);
  nand U20165(n19131,n16630,n17085,n19178);
  nand U20166(n19133,n19179,n19180);
  nand U20167(n19180,n16630,n17085);
  xor U20168(n19179,n17085,n19178);
  nand U20169(n19178,n19181,n19182);
  nand U20170(n19182,n16630,n17937);
  nand U20171(n19181,n16178,n17085);
  nand U20172(n19134,n19183,n19184);
  nand U20173(n19184,n19185,n19186);
  nor U20174(n19173,n16756,n19187);
  not U20175(n16756,n16629);
  xor U20176(n16629,n19154,n19188);
  and U20177(n19188,n19153,n19151);
  nand U20178(n19151,n19189,n19190);
  or U20179(n19153,n19189,n19190);
  nand U20180(n19190,n19191,n19192,n19193,n19194);
  nand U20181(n19194,n17974,n16178);
  nor U20182(n19193,n19195,n19196);
  nor U20183(n19196,n18774,n17774);
  nor U20184(n19195,n18775,n16759);
  nand U20185(n19192,n18339,G36349);
  nand U20186(n19191,n18340,G36317);
  xor U20187(n19189,n19197,n17976);
  nand U20188(n19197,n19198,n19199,n19200,n19201);
  nand U20189(n19201,n16178,n17973);
  nor U20190(n19200,n19202,n19203);
  nor U20191(n19203,n18730,n17774);
  nor U20192(n19202,n18731,n16759);
  not U20193(n16759,n16630);
  nand U20194(n16630,n19204,n19205,n19206);
  nand U20195(n19206,n17502,n17877);
  not U20196(n17502,n17774);
  nand U20197(n17774,n19207,n19208,n19209);
  nand U20198(n19208,n19210,n18466);
  nand U20199(n19207,G36221,n19211,G36249);
  nand U20200(n19205,n17851,G36156);
  nand U20201(n19204,n19212,n17852);
  nand U20202(n19199,n18348,G36317);
  nand U20203(n19198,n18347,G36349);
  nand U20204(n19154,n19213,n19214);
  nand U20205(n19214,n19215,n19216);
  nor U20206(n19172,n16604,n17987);
  not U20207(n16604,n16175);
  nand U20208(n16175,n19217,n19218,n19219,n19220);
  nand U20209(n19220,n19160,n17992);
  nor U20210(n19160,n19221,n19116);
  nor U20211(n19116,n17496,n17509);
  not U20212(n17509,G36442);
  nor U20213(n19221,G36454,G36442);
  nand U20214(n19219,G36350,n17882);
  nand U20215(n19218,G36318,n17883);
  nand U20216(n19217,G36286,n17881);
  nand U20217(n19170,G36349,n17843);
  nand U20218(n19169,n17993,n16181);
  nand U20219(n19168,n17929,n17496);
  nand U20220(G4454,n19222,n19223,n19224,n19225);
  nor U20221(n19225,n19226,n19227,n19228,n19229);
  nor U20222(n19229,n16952,n17956);
  and U20223(n19228,n16643,n17931);
  xnor U20224(n16643,n19230,n19185);
  nand U20225(n19185,n19231,n19232);
  nand U20226(n19232,n19233,n19234);
  nand U20227(n19230,n19186,n19183);
  nand U20228(n19183,n16642,n17085,n19235);
  nand U20229(n19186,n19236,n19237);
  nand U20230(n19237,n16642,n17085);
  xor U20231(n19236,n17085,n19235);
  nand U20232(n19235,n19238,n19239);
  nand U20233(n19239,n16642,n17937);
  nand U20234(n19238,n16181,n17085);
  and U20235(n19227,n16641,n17898);
  xor U20236(n16641,n19215,n19240);
  and U20237(n19240,n19213,n19216);
  or U20238(n19216,n19241,n19242);
  nand U20239(n19213,n19241,n19242);
  nand U20240(n19242,n19243,n19244,n19245,n19246);
  nand U20241(n19246,n17974,n16181);
  nor U20242(n19245,n19247,n19248);
  nor U20243(n19248,n18774,n17489);
  nor U20244(n19247,n18775,n16952);
  nand U20245(n19244,n18339,G36348);
  nand U20246(n19243,n18340,G36316);
  xor U20247(n19241,n19249,n17976);
  nand U20248(n19249,n19250,n19251,n19252,n19253);
  nand U20249(n19253,n16181,n17973);
  nor U20250(n19252,n19254,n19255);
  nor U20251(n19255,n18730,n17489);
  nor U20252(n19254,n18731,n16952);
  not U20253(n16952,n16642);
  nand U20254(n16642,n19256,n19257,n19258);
  nand U20255(n19258,n17490,n17877);
  not U20256(n17490,n17489);
  nand U20257(n17489,n19259,n19260);
  or U20258(n19260,G36220,G36249);
  nand U20259(n19259,G36249,n19261);
  nand U20260(n19257,n17851,G36155);
  nand U20261(n19256,n19262,n17852);
  nand U20262(n19251,n18348,G36316);
  nand U20263(n19250,n18347,G36348);
  nand U20264(n19215,n19263,n19264);
  nand U20265(n19264,n19265,n19266);
  nor U20266(n19226,n16616,n17987);
  not U20267(n16616,n16178);
  nand U20268(n16178,n19267,n19268,n19269,n19270);
  nand U20269(n19270,G36349,n17882);
  nand U20270(n19269,G36317,n17883);
  nand U20271(n19268,G36285,n17881);
  nand U20272(n19267,n17992,n17496);
  not U20273(n17496,G36454);
  nand U20274(n19224,G36348,n17843);
  nand U20275(n19223,n17993,n16184);
  nand U20276(n19222,n17929,G36435);
  nand U20277(G4453,n19271,n19272,n19273,n19274);
  nor U20278(n19274,n19275,n19276,n19277,n19278);
  nor U20279(n19278,n16800,n19159);
  not U20280(n16800,G36450);
  nor U20281(n19277,n16798,n17956);
  nor U20282(n19276,n17843,n19279,n19280);
  not U20283(n19280,n16653);
  xor U20284(n16653,n19266,n19281);
  and U20285(n19281,n19265,n19263);
  nand U20286(n19263,n19282,n19283);
  or U20287(n19265,n19282,n19283);
  nand U20288(n19283,n19284,n19285,n19286,n19287);
  nand U20289(n19287,n17974,n16184);
  nor U20290(n19286,n19288,n19289);
  nor U20291(n19289,n18774,n17472);
  nor U20292(n19288,n18775,n16798);
  not U20293(n18775,n17973);
  nand U20294(n19285,n18339,G36347);
  nand U20295(n19284,n18340,G36315);
  xor U20296(n19282,n19290,n17976);
  nand U20297(n19290,n19291,n19292,n19293,n19294);
  nand U20298(n19294,n16184,n17973);
  nor U20299(n19293,n19295,n19296);
  nor U20300(n19296,n18730,n17472);
  nor U20301(n19295,n18731,n16798);
  not U20302(n16798,n16654);
  nand U20303(n19292,n18348,G36315);
  nand U20304(n19291,n18347,G36347);
  nand U20305(n19266,n19297,n19298);
  nand U20306(n19298,n19299,n17976);
  nor U20307(n19279,n17024,n17439,n19300,n17022);
  not U20308(n19300,n17443);
  nand U20309(n17443,n19301,n17037);
  and U20310(n19275,n17843,G36347);
  nand U20311(n19273,n19302,n16181);
  nand U20312(n16181,n19303,n19304,n19305,n19306);
  nand U20313(n19306,G36348,n17882);
  nand U20314(n19305,G36316,n17883);
  nand U20315(n19304,G36284,n17881);
  nand U20316(n19303,G36435,n17992);
  nand U20317(n19272,n17931,n16655);
  xor U20318(n16655,n19234,n19307);
  and U20319(n19307,n19233,n19231);
  nand U20320(n19231,n16654,n17085,n19308);
  nand U20321(n19233,n19309,n19310);
  nand U20322(n19310,n16654,n17085);
  xor U20323(n19309,n17085,n19308);
  nand U20324(n19308,n19311,n19312);
  nand U20325(n19312,n16184,n17085);
  nand U20326(n19311,n16654,n17937);
  nand U20327(n16654,n19313,n19314,n19315);
  nand U20328(n19315,n17469,n17877);
  not U20329(n17469,n17472);
  nand U20330(n17472,n19316,n19317,n19318);
  nand U20331(n19317,n19319,n18466);
  nand U20332(n19316,G36219,G36218,G36249);
  nand U20333(n19314,n17851,G36154);
  nand U20334(n19313,n17852,n19320);
  nand U20335(n19234,n19321,n19322);
  nand U20336(n19322,n19323,n17937);
  nand U20337(n19271,n17993,n16187);
  nor U20338(n17993,n17843,n16325);
  nand U20339(n16325,n17009,n16994);
  not U20340(n16994,n16996);
  nand U20341(G4452,n19324,n19325,n19326,n19327);
  nor U20342(n19327,n19328,n19329,n19330);
  nor U20343(n19330,n16903,n19159);
  nor U20344(n17929,n17013,n17843);
  not U20345(n16903,G36440);
  nor U20346(n19329,n16902,n17956);
  nand U20347(n17956,n17844,n17006);
  and U20348(n19328,n17843,G36346);
  nand U20349(n19326,n17898,n16669);
  xnor U20350(n16669,n19331,n17976);
  nand U20351(n19331,n19297,n19299);
  nand U20352(n19299,n19332,n19333);
  not U20353(n19333,n19334);
  xor U20354(n19332,n19335,n17914);
  nand U20355(n19297,n19336,n19334);
  nand U20356(n19334,n19337,n19338,n19339,n19340);
  nand U20357(n19340,n16662,n17973);
  nor U20358(n19339,n19341,n19342);
  and U20359(n19342,n16187,n17974);
  nand U20360(n17974,n18731,n19343);
  nor U20361(n19341,n18774,n17462);
  not U20362(n18774,n18336);
  nand U20363(n18336,n18406,n18405);
  not U20364(n18405,n18347);
  not U20365(n18406,n18348);
  nand U20366(n19338,n18339,G36346);
  not U20367(n18339,n18397);
  nand U20368(n19337,n18340,G36314);
  not U20369(n18340,n18395);
  xor U20370(n19336,n17976,n19335);
  nand U20371(n19335,n19344,n19345,n19346,n19347);
  nand U20372(n19347,n18347,G36346);
  nor U20373(n18347,n17729,n17829);
  nor U20374(n19346,n19348,n19349);
  nor U20375(n19349,n18730,n17462);
  not U20376(n18730,n18349);
  nand U20377(n18349,n18395,n18397);
  nand U20378(n18397,n19350,n19351,n17447);
  nand U20379(n18395,n19350,n19351,n17729);
  nand U20380(n19350,n17835,n17028);
  nand U20381(n17028,n17444,n17304);
  not U20382(n17444,n16668);
  and U20383(n17835,n19352,n19353,n17872,n17013);
  nand U20384(n19353,n17010,n17020);
  not U20385(n19352,n17006);
  nand U20386(n17006,n19354,n16664);
  nand U20387(n16664,n17019,n17304);
  nor U20388(n17019,n17310,n16673,n16674);
  not U20389(n16673,n17311);
  or U20390(n19354,n16663,n16674);
  and U20391(n19348,G36314,n18348);
  nor U20392(n18348,n17829,n17447);
  not U20393(n17447,n17729);
  nand U20394(n17829,n19355,n19343);
  nand U20395(n19345,n16662,n17979);
  not U20396(n17979,n18731);
  nor U20397(n18731,n17909,n17912);
  not U20398(n17912,n17922);
  nand U20399(n17922,n17026,n19356);
  or U20400(n19356,n19357,n19358);
  not U20401(n17026,n17866);
  nand U20402(n17909,n19359,n19360);
  nand U20403(n19360,n19358,n17866);
  nand U20404(n19359,n19357,n19361);
  not U20405(n19361,n17939);
  nand U20406(n17939,n17037,n17866);
  nand U20407(n19344,n16187,n17973);
  nand U20408(n17923,n17310,n17010,n17866,n19351);
  not U20409(n17921,n17910);
  nor U20410(n17910,n17833,n19355,n17866);
  nor U20411(n17833,n17439,n19362);
  nor U20412(n19362,n16681,n17092);
  nor U20413(n17439,n17304,n17037,n17311);
  or U20414(n17924,n17940,n17311,n17037,n19355);
  nand U20415(n17940,n17020,n17866);
  nand U20416(n17866,n19363,n16287);
  nor U20417(n17914,n19358,n19357,n17250);
  nor U20418(n19357,n17023,n19355);
  nand U20419(n17023,n19301,n17304);
  and U20420(n19358,n19364,n19351);
  nand U20421(n19364,n17834,n19365);
  nand U20422(n19365,n17024,n19343);
  not U20423(n17024,n16671);
  nand U20424(n16671,n17037,n17020);
  nand U20425(n17834,n19301,n16674);
  not U20426(n17898,n19187);
  nand U20427(n19187,n17844,n19366);
  nand U20428(n19366,n16672,n19367);
  nand U20429(n19367,n17020,n16681);
  nor U20430(n16672,n17022,n19301);
  nor U20431(n19301,n17311,n17092);
  nor U20432(n17022,n17092,n17085);
  nand U20433(n19325,n17931,n16665);
  xor U20434(n16665,n19368,n17085);
  nand U20435(n19368,n19321,n19369);
  nand U20436(n19369,n19370,n19371);
  nand U20437(n19371,n16662,n17085);
  not U20438(n19370,n19323);
  nand U20439(n19321,n19323,n16662);
  nand U20440(n19323,n19372,n19373);
  nand U20441(n19373,n16187,n17085);
  nand U20442(n16187,n19374,n19375,n19376,n19377);
  nand U20443(n19377,G36346,n17882);
  nand U20444(n19376,G36314,n17883);
  nand U20445(n19375,G36282,n17881);
  nand U20446(n19374,G36440,n17992);
  nand U20447(n19372,n16902,n17937);
  not U20448(n16902,n16662);
  nand U20449(n16662,n19378,n19379,n19380);
  nand U20450(n19380,G36218,n17877);
  nand U20451(n19379,n17851,G36153);
  nand U20452(n19378,n19381,n17852);
  not U20453(n17877,n17838);
  not U20454(n17931,n19176);
  nand U20455(n19176,n17844,n19382);
  nand U20456(n19382,n16668,n16667,n17872);
  nand U20457(n17872,n16296,n17311);
  not U20458(n16296,n16666);
  nand U20459(n16666,n17092,n17937);
  nand U20460(n16667,n17010,n17092);
  not U20461(n17010,n16681);
  nand U20462(n16668,n17310,n17311,n17037);
  nand U20463(n19324,n19302,n16184);
  nand U20464(n16184,n19383,n19384,n19385,n19386);
  nand U20465(n19386,G36347,n17882);
  nand U20466(n19388,G36248,n19389,n18466);
  nand U20467(n19387,n19390,n19391,G36249);
  nand U20468(n19385,G36315,n17883);
  nand U20469(n19393,G36247,n19394,n18466);
  nand U20470(n19392,n19395,n19396,G36249);
  nand U20471(n19384,G36283,n17881);
  nand U20472(n19398,n19389,n19394,n18466);
  not U20473(n19389,G36247);
  nand U20474(n19397,n19396,n19391,G36249);
  not U20475(n19391,n19395);
  nand U20476(n19383,G36450,n17992);
  nand U20477(n17992,n19399,n19400);
  nand U20478(n19400,G36248,G36247,n18466);
  nand U20479(n19399,n19395,n19390,G36249);
  not U20480(n19302,n17987);
  nand U20481(n17987,n17844,n16675);
  not U20482(n16675,n16327);
  nand U20483(n16327,n17009,n16996);
  not U20484(n17844,n17843);
  nand U20485(n19401,n19402,n17013);
  or U20486(n17013,n16663,n17037);
  not U20487(n17037,n16674);
  nand U20488(n16663,n17025,n17304);
  nor U20489(n17025,n17311,n17310);
  nand U20490(n19402,n19363,n16678,n16676);
  not U20491(n16676,n16287);
  nand U20492(n16287,n19403,n19404);
  nand U20493(n19404,G36250,n19405);
  nand U20494(n19403,n16689,n19406);
  nand U20495(n16689,n19407,n19408);
  and U20496(n16678,n17027,n17002);
  nand U20497(n17002,n17009,n16681);
  nand U20498(n16681,n17311,n16674);
  nand U20499(n16674,n19409,n19410,n19411);
  nand U20500(n19410,n19412,n18466);
  nand U20501(n19409,G36238,n19413,G36249);
  nand U20502(n17311,n19414,n19415,n19413);
  nand U20503(n19415,n19416,n18466);
  nand U20504(n19414,G36237,n19417,G36249);
  not U20505(n17009,n17090);
  nand U20506(n17027,n19405,n19418);
  nand U20507(n19418,n19419,n19420,n19421,n19422);
  nor U20508(n19422,n19423,n19424,n19425,n19426);
  nand U20509(n19426,n19427,n19428,n19429);
  nand U20510(n19425,n19430,n19431,n19432,n19433);
  nand U20511(n19424,n19434,n19435,n19436,n19437);
  nand U20512(n19423,n19438,n19439,n19440,n19441);
  nor U20513(n19421,n19442,G36252,G36254,G36253);
  nand U20514(n19442,n19443,n19444,n19445,n19446);
  nor U20515(n19420,G36266,G36265,G36264,G36263);
  nor U20516(n19419,G36262,G36261,G36260,G36259);
  not U20517(n19405,n19406);
  not U20518(n19363,n16680);
  nand U20519(n16680,n16686,n19447);
  or U20520(n19447,n19406,G36251);
  nand U20521(n16686,n19408,n19448);
  nor U20522(G4451,n16685,n19441);
  not U20523(n19441,G36281);
  nor U20524(G4450,n16685,n19440);
  not U20525(n19440,G36280);
  nor U20526(G4449,n16685,n19439);
  not U20527(n19439,G36279);
  nor U20528(G4448,n16685,n19438);
  not U20529(n19438,G36278);
  nor U20530(G4447,n16685,n19437);
  not U20531(n19437,G36277);
  nor U20532(G4446,n16685,n19436);
  not U20533(n19436,G36276);
  nor U20534(G4445,n16685,n19435);
  not U20535(n19435,G36275);
  nor U20536(G4444,n16685,n19434);
  not U20537(n19434,G36274);
  nor U20538(G4443,n16685,n19433);
  not U20539(n19433,G36273);
  nor U20540(G4442,n16685,n19432);
  not U20541(n19432,G36272);
  nor U20542(G4441,n16685,n19431);
  not U20543(n19431,G36271);
  nor U20544(G4440,n16685,n19430);
  not U20545(n19430,G36270);
  nor U20546(G4439,n16685,n19428);
  not U20547(n19428,G36269);
  nor U20548(G4438,n16685,n19427);
  not U20549(n19427,G36268);
  nor U20550(G4437,n16685,n19429);
  not U20551(n19429,G36267);
  and U20552(G4436,n16684,G36266);
  and U20553(G4435,n16684,G36265);
  and U20554(G4434,n16684,G36264);
  and U20555(G4433,n16684,G36263);
  and U20556(G4432,n16684,G36262);
  and U20557(G4431,n16684,G36261);
  and U20558(G4430,n16684,G36260);
  and U20559(G4429,n16684,G36259);
  nor U20560(G4428,n16685,n19446);
  not U20561(n19446,G36258);
  nor U20562(G4427,n16685,n19445);
  not U20563(n19445,G36257);
  nor U20564(G4426,n16685,n19444);
  not U20565(n19444,G36256);
  nor U20566(G4425,n16685,n19443);
  not U20567(n19443,G36255);
  not U20568(n16685,n16684);
  and U20569(G4424,n16684,G36254);
  and U20570(G4423,n16684,G36253);
  and U20571(G4422,n16684,G36252);
  nand U20572(n16684,n16677,n19406);
  nand U20573(n19406,n19449,n19450,n19451);
  not U20574(n19451,n19408);
  nand U20575(n19450,n19452,n19448,n17876);
  not U20576(n17876,G36430);
  nand U20577(n19449,n19407,n19448,G36430);
  nor U20578(n16677,n19355,G4389,n17250);
  nand U20579(G4421,n19453,n19454,n19455);
  nand U20580(n19455,n19456,n17853);
  nand U20581(n19454,n19457,n19394,n19458);
  not U20582(n19394,G36248);
  nand U20583(n19453,n19459,G36184);
  nand U20584(G4420,n19460,n19461,n19462,n19463);
  nand U20585(n19463,n19458,n19390);
  not U20586(n19390,n19396);
  xor U20587(n19396,n19457,G36248);
  nand U20588(n19462,n19459,G36183);
  nand U20589(n19461,n19464,G36248);
  nand U20590(n19460,n19456,n17869);
  nand U20591(G4419,n19465,n19466,n19467,n19468);
  nand U20592(n19468,n19458,n19395);
  nor U20593(n19395,n19457,n19469);
  and U20594(n19469,G36247,n19470);
  nor U20595(n19457,n19470,G36247);
  nand U20596(n19467,n19459,G36182);
  nand U20597(n19466,n19464,G36247);
  nand U20598(n19465,n19456,n17943);
  nand U20599(G4418,n19471,n19472,n19473,n19474);
  nand U20600(n19474,G36246,n19475);
  nand U20601(n19475,n19476,n19477);
  nand U20602(n19477,n19458,n19478);
  nand U20603(n19473,n19458,n19479,n19480);
  nand U20604(n19472,n19459,G36181);
  nand U20605(n19471,n19456,n17982);
  nand U20606(G4417,n19481,n19482,n19483,n19484);
  nand U20607(n19484,n19485,n19479,n19458);
  nand U20608(n19483,n19459,G36180);
  nand U20609(n19482,n19464,G36245);
  nand U20610(n19481,n19456,n18022);
  nand U20611(G4416,n19486,n19487,n19488,n19489);
  nand U20612(n19489,n19490,n19491,n19458);
  nand U20613(n19488,n19459,G36179);
  nand U20614(n19487,n19464,G36244);
  nand U20615(n19486,n19456,n18063);
  nand U20616(G4415,n19492,n19493,n19494,n19495);
  nand U20617(n19495,G36243,n19496);
  nand U20618(n19496,n19476,n19497);
  nand U20619(n19497,n19458,n19498);
  nand U20620(n19494,n19458,n19499,n19500);
  nand U20621(n19493,n19459,G36178);
  nand U20622(n19492,n19456,n18105);
  nand U20623(G4414,n19501,n19502,n19503,n19504);
  nand U20624(n19504,n19505,n19499,n19458);
  nand U20625(n19503,n19459,G36177);
  nand U20626(n19502,n19464,G36242);
  nand U20627(n19501,n19456,n18143);
  nand U20628(G4413,n19506,n19507,n19508,n19509);
  nand U20629(n19509,G36241,n19510);
  nand U20630(n19510,n19476,n19511);
  nand U20631(n19511,n19458,n19512);
  nand U20632(n19508,n19458,n19513,n19514);
  nand U20633(n19507,n19459,G36176);
  nand U20634(n19506,n19456,n18182);
  nand U20635(G4412,n19515,n19516,n19517,n19518);
  nand U20636(n19518,n19519,n19513,n19458);
  nand U20637(n19517,n19459,G36175);
  nand U20638(n19516,n19464,G36240);
  nand U20639(n19515,n19456,n18224);
  nand U20640(G4411,n19520,n19521,n19522,n19523);
  nand U20641(n19523,n19524,n19525,n19458);
  nand U20642(n19522,n19459,G36174);
  nand U20643(n19521,n19464,G36239);
  nand U20644(n19520,n19456,n18261);
  nand U20645(G4410,n19526,n19527,n19528,n19529);
  nand U20646(n19529,G36238,n19530);
  nand U20647(n19530,n19476,n19531);
  nand U20648(n19531,n19458,n19532);
  nand U20649(n19528,n19458,n19413,n19412);
  nand U20650(n19527,n19459,G36173);
  nand U20651(n19526,n19456,n18301);
  nand U20652(G4409,n19533,n19534,n19535,n19536);
  nand U20653(n19536,G36237,n19537);
  nand U20654(n19537,n19476,n19538);
  nand U20655(n19538,n19458,n19539);
  nand U20656(n19535,n19458,n19417,n19416);
  nand U20657(n19534,n19459,G36172);
  nand U20658(n19533,n19456,n18353);
  nand U20659(G4408,n19540,n19541,n19542,n19543);
  or U20660(n19543,n18413,n19544);
  nand U20661(n18413,n19417,n19545);
  nand U20662(n19545,G36236,n18464);
  not U20663(n19417,n19539);
  nand U20664(n19542,n19459,G36171);
  nand U20665(n19541,n19464,G36236);
  nand U20666(n19540,n19456,n18410);
  nand U20667(G4407,n19546,n19547,n19548,n19549);
  nand U20668(n19549,G36235,n19550);
  nand U20669(n19550,n19476,n19551);
  nand U20670(n19551,n19458,n19552);
  nand U20671(n19548,n19458,n18467,n18465);
  nand U20672(n19547,n19459,G36170);
  nand U20673(n19546,n19456,n18461);
  nand U20674(G4406,n19553,n19554,n19555,n19556);
  or U20675(n19556,n18521,n19544);
  nand U20676(n18521,n18467,n19557);
  nand U20677(n19557,G36234,n18571);
  not U20678(n18467,n19552);
  nand U20679(n19555,n19459,G36169);
  nand U20680(n19554,n19464,G36234);
  nand U20681(n19553,n19456,n18518);
  nand U20682(G4405,n19558,n19559,n19560,n19561);
  nand U20683(n19561,G36233,n19562);
  nand U20684(n19562,n19476,n19563);
  nand U20685(n19563,n19458,n19564);
  nand U20686(n19560,n19458,n18573,n18572);
  nand U20687(n19559,n19459,G36168);
  nand U20688(n19558,n19456,n18568);
  nand U20689(G4404,n19565,n19566,n19567,n19568);
  or U20690(n19568,n18629,n19544);
  nand U20691(n18629,n18573,n19569);
  nand U20692(n19569,G36232,n18681);
  not U20693(n18573,n19564);
  nand U20694(n19567,n19459,G36167);
  nand U20695(n19566,n19464,G36232);
  nand U20696(n19565,n19456,n18626);
  nand U20697(G4403,n19570,n19571,n19572,n19573);
  nand U20698(n19573,G36231,n19574);
  nand U20699(n19574,n19476,n19575);
  nand U20700(n19575,n19458,n19576);
  nand U20701(n19572,n19458,n18683,n18682);
  nand U20702(n19571,n19459,G36166);
  nand U20703(n19570,n19456,n18678);
  nand U20704(G4402,n19577,n19578,n19579,n19580);
  or U20705(n19580,n18737,n19544);
  nand U20706(n18737,n18683,n19581);
  nand U20707(n19581,G36230,n18788);
  not U20708(n18683,n19576);
  nand U20709(n19579,n19459,G36165);
  nand U20710(n19578,n19464,G36230);
  nand U20711(n19577,n19456,n18738);
  nand U20712(G4401,n19582,n19583,n19584,n19585);
  nand U20713(n19585,G36229,n19586);
  nand U20714(n19586,n19476,n19587);
  nand U20715(n19587,n19458,n19588);
  nand U20716(n19584,n19458,n18790,n18789);
  nand U20717(n19583,n19459,G36164);
  nand U20718(n19582,n19456,n18791);
  nand U20719(G4400,n19589,n19590,n19591,n19592);
  or U20720(n19592,n18842,n19544);
  nand U20721(n18842,n18790,n19593);
  nand U20722(n19593,G36228,n18895);
  not U20723(n18790,n19588);
  nand U20724(n19591,n19459,G36163);
  nand U20725(n19590,n19464,G36228);
  nand U20726(n19589,n19456,n18843);
  nand U20727(G4399,n19594,n19595,n19596,n19597);
  nand U20728(n19597,G36227,n19598);
  nand U20729(n19598,n19476,n19599);
  nand U20730(n19599,n19458,n19600);
  nand U20731(n19596,n19458,n18897,n18896);
  nand U20732(n19595,n19459,G36162);
  nand U20733(n19594,n19456,n18898);
  nand U20734(G4398,n19601,n19602,n19603,n19604);
  or U20735(n19604,n18945,n19544);
  nand U20736(n18945,n18897,n19605);
  nand U20737(n19605,G36226,n18999);
  not U20738(n18897,n19600);
  nand U20739(n19603,n19459,G36161);
  nand U20740(n19602,n19464,G36226);
  nand U20741(n19601,n19456,n18946);
  nand U20742(G4397,n19606,n19607,n19608,n19609);
  nand U20743(n19609,G36225,n19610);
  nand U20744(n19610,n19476,n19611);
  nand U20745(n19611,n19458,n19612);
  nand U20746(n19608,n19458,n19001,n19000);
  nand U20747(n19607,n19459,G36160);
  nand U20748(n19606,n19456,n19002);
  nand U20749(G4396,n19613,n19614,n19615,n19616);
  or U20750(n19616,n19052,n19544);
  nand U20751(n19052,n19001,n19617);
  nand U20752(n19617,G36224,n19102);
  not U20753(n19001,n19612);
  nand U20754(n19615,n19459,G36159);
  nand U20755(n19614,n19464,G36224);
  nand U20756(n19613,n19456,n19053);
  nand U20757(G4395,n19618,n19619,n19620,n19621);
  nand U20758(n19621,G36223,n19622);
  nand U20759(n19622,n19476,n19623);
  nand U20760(n19623,n19458,n19624);
  nand U20761(n19620,n19458,n19104,n19103);
  nand U20762(n19619,n19459,G36158);
  nand U20763(n19618,n19456,n19105);
  nand U20764(G4394,n19625,n19626,n19627,n19628);
  or U20765(n19628,n19166,n19544);
  nand U20766(n19166,n19104,n19629);
  nand U20767(n19629,G36222,n19209);
  not U20768(n19104,n19624);
  nand U20769(n19627,n19459,G36157);
  nand U20770(n19626,n19464,G36222);
  nand U20771(n19625,n19456,n19167);
  nand U20772(G4393,n19630,n19631,n19632,n19633);
  nand U20773(n19633,G36221,n19634);
  nand U20774(n19634,n19476,n19635);
  nand U20775(n19635,n19458,n19636);
  nand U20776(n19632,n19458,n19211,n19210);
  nand U20777(n19631,n19459,G36156);
  nand U20778(n19630,n19456,n19212);
  nand U20779(G4392,n19637,n19638,n19639,n19640);
  or U20780(n19640,n19261,n19544);
  nand U20781(n19261,n19211,n19641);
  nand U20782(n19641,G36220,n19318);
  not U20783(n19211,n19636);
  nand U20784(n19639,n19459,G36155);
  nand U20785(n19638,n19464,G36220);
  not U20786(n19464,n19476);
  nand U20787(n19637,n19456,n19262);
  nand U20788(G4391,n19642,n19643,n19644,n19645);
  nand U20789(n19645,G36219,n19646);
  nand U20790(n19646,n19476,n19647);
  nand U20791(n19647,n19458,n17462);
  nand U20792(n19644,n19458,G36218,n19319);
  nand U20793(n19643,n19459,G36154);
  nand U20794(n19642,n19456,n19320);
  nand U20795(G4390,n19648,n19649,n19650);
  nand U20796(n19650,n19456,n19381);
  nand U20797(n19649,G36218,n19651);
  nand U20798(n19651,n19476,n19544);
  nand U20799(n19544,n19476,G36460);
  nand U20800(n19476,G36460,n18466);
  nand U20801(n19648,n19459,G36153);
  nand U20802(G4388,n17837,n19652);
  nand U20803(n19652,n17090,n19351,n17838);
  not U20804(n19351,n19355);
  nor U20805(n19355,n19408,n19407,n19448);
  nand U20806(n19448,n19653,n19654,n19655);
  nand U20807(n19654,n19500,n18466);
  nand U20808(n19653,G36243,n19499,G36249);
  not U20809(n19407,n19452);
  nand U20810(n19452,n19656,n19657);
  nand U20811(n19657,G36242,n18466);
  nand U20812(n19656,n19505,n19499,G36249);
  not U20813(n19499,n19498);
  nand U20814(n19505,G36242,n19658);
  nand U20815(n19658,n19512,n19514);
  not U20816(n19514,G36241);
  nand U20817(n19408,n19659,n19660);
  or U20818(n19660,G36244,G36249);
  nand U20819(n19659,G36249,n19661);
  nand U20820(n19661,n19491,n19490);
  nand U20821(n19490,G36244,n19655);
  nand U20822(n17090,n17310,n17020);
  not U20823(n17020,n17304);
  nand U20824(n17304,n19662,n19663);
  or U20825(n19663,G36239,G36249);
  nand U20826(n19662,G36249,n19664);
  nand U20827(n19664,n19525,n19524);
  nand U20828(n19524,G36239,n19411);
  not U20829(n17310,n17092);
  nand U20830(n17092,n19665,n19666);
  or U20831(n19666,G36240,G36249);
  nand U20832(n19665,G36249,n19667);
  nand U20833(n19667,n19513,n19519);
  nand U20834(n19519,G36240,n19525);
  and U20835(n17837,n19668,G36460);
  nand U20836(n19668,n17250,n17838);
  nand U20837(n17838,n17729,n16996);
  nand U20838(n16996,n19669,n19670,n19470);
  nand U20839(n19470,n19478,n19480);
  nand U20840(n19670,n19480,n18466);
  not U20841(n18466,G36249);
  not U20842(n19480,G36246);
  nand U20843(n19669,G36246,n19479,G36249);
  nand U20844(n17729,n19671,n19672);
  or U20845(n19672,G36245,G36249);
  nand U20846(n19671,G36249,n19673);
  nand U20847(n19673,n19479,n19485);
  nand U20848(n19485,G36245,n19491);
  not U20849(n19479,n19478);
  nor U20850(n19478,n19491,G36245);
  or U20851(n19491,n19655,G36244);
  nand U20852(n19655,n19498,n19500);
  not U20853(n19500,G36243);
  nor U20854(n19498,G36241,G36242,n19513);
  not U20855(n17250,n19343);
  xor U20856(n19343,n19674,G36241);
  nand U20857(n19674,G36249,n19513);
  not U20858(n19513,n19512);
  nor U20859(n19512,n19525,G36240);
  or U20860(n19525,n19411,G36239);
  nand U20861(n19411,n19532,n19412);
  not U20862(n19412,G36238);
  not U20863(n19532,n19413);
  nand U20864(n19413,n19539,n19416);
  not U20865(n19416,G36237);
  nor U20866(n19539,n18464,G36236);
  nand U20867(n18464,n19552,n18465);
  not U20868(n18465,G36235);
  nor U20869(n19552,n18571,G36234);
  nand U20870(n18571,n19564,n18572);
  not U20871(n18572,G36233);
  nor U20872(n19564,n18681,G36232);
  nand U20873(n18681,n19576,n18682);
  not U20874(n18682,G36231);
  nor U20875(n19576,n18788,G36230);
  nand U20876(n18788,n19588,n18789);
  not U20877(n18789,G36229);
  nor U20878(n19588,n18895,G36228);
  nand U20879(n18895,n19600,n18896);
  not U20880(n18896,G36227);
  nor U20881(n19600,n18999,G36226);
  nand U20882(n18999,n19612,n19000);
  not U20883(n19000,G36225);
  nor U20884(n19612,n19102,G36224);
  nand U20885(n19102,n19624,n19103);
  not U20886(n19103,G36223);
  nor U20887(n19624,n19209,G36222);
  nand U20888(n19209,n19636,n19210);
  not U20889(n19210,G36221);
  nor U20890(n19636,n19318,G36220);
  nand U20891(n19318,n17462,n19319);
  not U20892(n19319,G36219);
  not U20893(n17462,G36218);
  nand U20894(G1860,n19675,n19676);
  nand U20895(n19676,G36184,n19677);
  nand U20896(n19675,G1625,n19678);
  nand U20897(G1859,n19679,n19680);
  nand U20898(n19680,G36183,n19677);
  nand U20899(n19679,G1625,n19681);
  nand U20900(G1858,n19682,n19683);
  nand U20901(n19683,G36182,n19677);
  nand U20902(n19682,G1625,n19684);
  nand U20903(G1857,n19685,n19686);
  nand U20904(n19686,G36181,n19677);
  nand U20905(n19685,G1625,n19687);
  nand U20906(G1856,n19688,n19689);
  nand U20907(n19689,G36180,n19677);
  nand U20908(n19688,G1625,n19690);
  nand U20909(G1855,n19691,n19692);
  nand U20910(n19692,G36179,n19677);
  nand U20911(n19691,G1625,n19693);
  nand U20912(G1854,n19694,n19695);
  nand U20913(n19695,G36178,n19677);
  nand U20914(n19694,G1625,n19696);
  nand U20915(G1853,n19697,n19698);
  nand U20916(n19698,G36177,n19677);
  nand U20917(n19697,G1625,n19699);
  nand U20918(G1852,n19700,n19701);
  nand U20919(n19701,G36176,n19677);
  nand U20920(n19700,G1625,n19702);
  nand U20921(G1851,n19703,n19704);
  nand U20922(n19704,G36175,n19677);
  nand U20923(n19703,G1625,n19705);
  nand U20924(G1850,n19706,n19707);
  nand U20925(n19707,G36174,n19677);
  nand U20926(n19706,G1625,n19708);
  nand U20927(G1849,n19709,n19710);
  nand U20928(n19710,G36173,n19677);
  nand U20929(n19709,G1625,n19711);
  nand U20930(G1848,n19712,n19713);
  nand U20931(n19713,G36172,n19677);
  nand U20932(n19712,G1625,n19714);
  nand U20933(G1847,n19715,n19716);
  nand U20934(n19716,G36171,n19677);
  nand U20935(n19715,G1625,n19717);
  nand U20936(G1846,n19718,n19719);
  nand U20937(n19719,G36170,n19677);
  nand U20938(n19718,G1625,n19720);
  nand U20939(G1845,n19721,n19722);
  nand U20940(n19722,G36169,n19677);
  nand U20941(n19721,G1625,n19723);
  nand U20942(G1844,n19724,n19725);
  nand U20943(n19725,G36168,n19677);
  nand U20944(n19724,G1625,n19726);
  nand U20945(G1843,n19727,n19728);
  nand U20946(n19728,G36167,n19677);
  nand U20947(n19727,G1625,n19729);
  nand U20948(G1842,n19730,n19731);
  nand U20949(n19731,G36166,n19677);
  nand U20950(n19730,G1625,n19732);
  nand U20951(G1841,n19733,n19734);
  nand U20952(n19734,G36165,n19677);
  nand U20953(n19733,G1625,n19735);
  nand U20954(G1840,n19736,n19737);
  nand U20955(n19737,G36164,n19677);
  nand U20956(n19736,G1625,n19738);
  nand U20957(G1839,n19739,n19740);
  nand U20958(n19740,G36163,n19677);
  nand U20959(n19739,G1625,n19741);
  nand U20960(G1838,n19742,n19743);
  nand U20961(n19743,G36162,n19677);
  nand U20962(n19742,G1625,n19744);
  nand U20963(G1837,n19745,n19746);
  nand U20964(n19746,G36161,n19677);
  nand U20965(n19745,G1625,n19747);
  nand U20966(G1836,n19748,n19749);
  nand U20967(n19749,G36160,n19677);
  nand U20968(n19748,G1625,n19750);
  nand U20969(G1835,n19751,n19752);
  nand U20970(n19752,G36159,n19677);
  nand U20971(n19751,G1625,n19753);
  nand U20972(G1834,n19754,n19755);
  nand U20973(n19755,G36158,n19677);
  nand U20974(n19754,G1625,n19756);
  nand U20975(G1833,n19757,n19758);
  nand U20976(n19758,G36157,n19677);
  nand U20977(n19757,G1625,n19759);
  nand U20978(G1832,n19760,n19761);
  nand U20979(n19761,G36156,n19677);
  nand U20980(n19760,G1625,n19762);
  nand U20981(G1831,n19763,n19764);
  nand U20982(n19764,G36155,n19677);
  nand U20983(n19763,G1625,n19765);
  nand U20984(G1830,n19766,n19767);
  nand U20985(n19767,G36154,n19677);
  nand U20986(n19766,G1625,n19768);
  nand U20987(G1829,n19769,n19770);
  nand U20988(n19770,G36153,n19677);
  nand U20989(n19769,G1625,n19771);
  nand U20990(G1828,n19772,n19773,n19774,n19775);
  nor U20991(n19775,n19776,n19777,n19778,n19779);
  nor U20992(n19779,n19780,n19781);
  nor U20993(n19777,n19783,n19784,n19785);
  not U20994(n19785,n19786);
  nor U20995(n19784,n19787,n19788);
  nor U20996(n19776,n19789,n19790);
  nand U20997(n19774,n19791,n19765);
  nand U20998(n19773,n19792,n19793);
  nand U20999(n19772,n19794,n19795);
  nand U21000(G1827,n19796,n19797);
  nand U21001(n19797,n19798,n19799);
  nand U21002(n19796,G36100,n19800);
  nand U21003(G1826,n19801,n19802);
  nand U21004(n19802,G36099,n19800);
  nand U21005(n19801,n19798,n19803);
  nand U21006(G1825,n19804,n19805);
  nand U21007(n19805,G36098,n19800);
  nand U21008(n19804,n19798,n19806);
  nand U21009(G1824,n19807,n19808);
  nand U21010(n19808,G36097,n19800);
  nand U21011(n19807,n19798,n19809);
  nand U21012(G1823,n19810,n19811);
  nand U21013(n19811,G36096,n19800);
  nand U21014(n19810,n19798,n19812);
  nand U21015(G1822,n19813,n19814);
  nand U21016(n19814,G36095,n19800);
  nand U21017(n19813,n19798,n19815);
  nand U21018(G1821,n19816,n19817);
  nand U21019(n19817,G36094,n19800);
  nand U21020(n19816,n19798,n19818);
  nand U21021(G1820,n19819,n19820);
  nand U21022(n19820,G36093,n19800);
  nand U21023(n19819,n19798,n19821);
  nand U21024(G1819,n19822,n19823);
  nand U21025(n19823,G36092,n19800);
  nand U21026(n19822,n19798,n19824);
  nand U21027(G1818,n19825,n19826);
  nand U21028(n19826,G36091,n19800);
  nand U21029(n19825,n19798,n19827);
  nand U21030(G1817,n19828,n19829);
  nand U21031(n19829,G36090,n19800);
  nand U21032(n19828,n19798,n19830);
  nand U21033(G1816,n19831,n19832);
  nand U21034(n19832,G36089,n19800);
  nand U21035(n19831,n19798,n19833);
  nand U21036(G1815,n19834,n19835);
  nand U21037(n19835,G36088,n19800);
  nand U21038(n19834,n19798,n19836);
  nand U21039(G1814,n19837,n19838);
  nand U21040(n19838,G36087,n19800);
  nand U21041(n19837,n19798,n19839);
  nand U21042(G1813,n19840,n19841);
  nand U21043(n19841,G36086,n19800);
  nand U21044(n19840,n19798,n19842);
  nand U21045(G1812,n19843,n19844);
  nand U21046(n19844,G36085,n19800);
  nand U21047(n19843,n19798,n19845);
  nand U21048(G1811,n19846,n19847);
  nand U21049(n19847,G36084,n19800);
  nand U21050(n19846,n19798,n19848);
  nand U21051(G1810,n19849,n19850);
  nand U21052(n19850,G36083,n19800);
  nand U21053(n19849,n19798,n19851);
  nand U21054(G1809,n19852,n19853);
  nand U21055(n19853,G36082,n19800);
  nand U21056(n19852,n19798,n19854);
  nand U21057(G1808,n19855,n19856);
  nand U21058(n19856,G36081,n19800);
  nand U21059(n19855,n19798,n19857);
  nand U21060(G1807,n19858,n19859);
  nand U21061(n19859,G36080,n19800);
  nand U21062(n19858,n19798,n19860);
  nand U21063(G1806,n19861,n19862);
  nand U21064(n19862,G36079,n19800);
  nand U21065(n19861,n19798,n19863);
  nand U21066(G1805,n19864,n19865);
  nand U21067(n19865,G36078,n19800);
  nand U21068(n19864,n19798,n19866);
  nand U21069(G1804,n19867,n19868);
  nand U21070(n19868,G36077,n19800);
  nand U21071(n19867,n19798,n19869);
  nand U21072(G1803,n19870,n19871);
  nand U21073(n19871,G36076,n19800);
  nand U21074(n19870,n19798,n19872);
  nand U21075(G1802,n19873,n19874);
  nand U21076(n19874,G36075,n19800);
  nand U21077(n19873,n19798,n19875);
  nand U21078(G1801,n19876,n19877);
  nand U21079(n19877,G36074,n19800);
  nand U21080(n19876,n19798,n19878);
  nand U21081(G1800,n19879,n19880);
  nand U21082(n19880,G36073,n19800);
  nand U21083(n19879,n19798,n19881);
  nand U21084(G1799,n19882,n19883);
  nand U21085(n19883,G36072,n19800);
  nand U21086(n19882,n19798,n19884);
  nand U21087(G1798,n19885,n19886);
  nand U21088(n19886,G36071,n19800);
  nand U21089(n19885,n19798,n19887);
  nand U21090(G1797,n19888,n19889);
  nand U21091(n19889,G36070,n19800);
  nand U21092(n19888,n19798,n19890);
  nand U21093(G1796,n19891,n19892);
  nand U21094(n19892,G36069,n19800);
  nand U21095(n19891,n19798,n19893);
  nand U21096(G1795,n19896,n19897);
  nand U21097(n19897,n19898,n19799);
  nand U21098(n19799,n19899,n19900,n19901);
  nand U21099(n19901,n19902,n19903);
  nand U21100(n19899,n19904,n19905);
  nand U21101(n19896,G36068,n19906);
  nand U21102(G1794,n19907,n19908);
  nand U21103(n19908,n19898,n19803);
  nand U21104(n19803,n19909,n19900,n19910);
  nand U21105(n19910,n19904,n19911);
  nand U21106(n19909,n19912,n19913,n19903);
  nand U21107(n19907,G36067,n19906);
  nand U21108(G1793,n19914,n19915);
  nand U21109(n19915,n19898,n19806);
  nand U21110(n19806,n19916,n19917,n19918,n19919);
  nand U21111(n19918,n19904,n19920);
  nand U21112(n19917,n19921,n19922);
  nand U21113(n19916,n19923,n19924);
  nand U21114(n19914,G36066,n19906);
  nand U21115(G1792,n19925,n19926);
  nand U21116(n19926,n19898,n19809);
  nand U21117(n19809,n19927,n19928,n19929,n19930);
  nor U21118(n19930,n19931,n19932);
  nor U21119(n19932,n19933,n19934);
  nor U21120(n19931,n19935,n19936);
  nand U21121(n19929,n19937,n19924);
  nand U21122(n19928,n19904,n19938);
  nand U21123(n19927,n19939,n19922);
  nand U21124(n19925,G36065,n19906);
  nand U21125(G1791,n19940,n19941);
  nand U21126(n19941,n19898,n19812);
  nand U21127(n19812,n19942,n19943,n19944,n19945);
  nor U21128(n19945,n19946,n19947);
  nor U21129(n19947,n19948,n19934);
  nor U21130(n19946,n19949,n19936);
  nand U21131(n19944,n19950,n19924);
  nand U21132(n19943,n19904,n19951);
  nand U21133(n19942,n19952,n19922);
  nand U21134(n19940,G36064,n19906);
  nand U21135(G1790,n19953,n19954);
  nand U21136(n19954,n19898,n19815);
  nand U21137(n19815,n19955,n19956,n19957,n19958);
  nor U21138(n19958,n19959,n19960);
  nor U21139(n19960,n19961,n19934);
  nor U21140(n19959,n19933,n19936);
  nand U21141(n19957,n19962,n19924);
  nand U21142(n19956,n19904,n19963);
  nand U21143(n19955,n19964,n19922);
  nand U21144(n19953,G36063,n19906);
  nand U21145(G1789,n19965,n19966);
  nand U21146(n19966,n19898,n19818);
  nand U21147(n19818,n19967,n19968,n19969,n19970);
  nor U21148(n19970,n19971,n19972);
  nor U21149(n19972,n19973,n19934);
  nor U21150(n19971,n19948,n19936);
  nand U21151(n19969,n19974,n19924);
  nand U21152(n19968,n19904,n19975);
  nand U21153(n19967,n19976,n19922);
  nand U21154(n19965,G36062,n19906);
  nand U21155(G1788,n19977,n19978);
  nand U21156(n19978,n19898,n19821);
  nand U21157(n19821,n19979,n19980,n19981,n19982);
  nor U21158(n19982,n19983,n19984);
  nor U21159(n19984,n19985,n19934);
  nor U21160(n19983,n19961,n19936);
  nand U21161(n19981,n19986,n19924);
  nand U21162(n19980,n19904,n19987);
  nand U21163(n19979,n19988,n19922);
  nand U21164(n19977,G36061,n19906);
  nand U21165(G1787,n19989,n19990);
  nand U21166(n19990,n19898,n19824);
  nand U21167(n19824,n19991,n19992,n19993,n19994);
  nor U21168(n19994,n19995,n19996);
  nor U21169(n19996,n19997,n19934);
  nor U21170(n19995,n19973,n19936);
  nand U21171(n19993,n19998,n19924);
  nand U21172(n19992,n19904,n19999);
  nand U21173(n19991,n20000,n19922);
  nand U21174(n19989,G36060,n19906);
  nand U21175(G1786,n20001,n20002);
  nand U21176(n20002,n19898,n19827);
  nand U21177(n19827,n20003,n20004,n20005,n20006);
  nor U21178(n20006,n20007,n20008);
  nor U21179(n20008,n20009,n19934);
  nor U21180(n20007,n19985,n19936);
  nand U21181(n20005,n20010,n19924);
  nand U21182(n20004,n19904,n20011);
  nand U21183(n20003,n20012,n19922);
  nand U21184(n20001,G36059,n19906);
  nand U21185(G1785,n20013,n20014);
  nand U21186(n20014,n19898,n19830);
  nand U21187(n19830,n20015,n20016,n20017,n20018);
  nor U21188(n20018,n20019,n20020);
  nor U21189(n20020,n20021,n19934);
  nor U21190(n20019,n19997,n19936);
  nand U21191(n20017,n20022,n19924);
  nand U21192(n20016,n19904,n20023);
  nand U21193(n20015,n20024,n19922);
  nand U21194(n20013,G36058,n19906);
  nand U21195(G1784,n20025,n20026);
  nand U21196(n20026,n19898,n19833);
  nand U21197(n19833,n20027,n20028,n20029,n20030);
  nor U21198(n20030,n20031,n20032);
  nor U21199(n20032,n20033,n19934);
  nor U21200(n20031,n20009,n19936);
  nand U21201(n20029,n20034,n19924);
  nand U21202(n20028,n19904,n20035);
  nand U21203(n20027,n20036,n19922);
  nand U21204(n20025,G36057,n19906);
  nand U21205(G1783,n20037,n20038);
  nand U21206(n20038,n19898,n19836);
  nand U21207(n19836,n20039,n20040,n20041,n20042);
  nor U21208(n20042,n20043,n20044);
  nor U21209(n20044,n20045,n19934);
  nor U21210(n20043,n20021,n19936);
  nand U21211(n20041,n20046,n19924);
  nand U21212(n20040,n19904,n20047);
  nand U21213(n20039,n20048,n19922);
  nand U21214(n20037,G36056,n19906);
  nand U21215(G1781,n20049,n20050);
  nand U21216(n20050,n19898,n19839);
  nand U21217(n19839,n20051,n20052,n20053,n20054);
  nor U21218(n20054,n20055,n20056);
  nor U21219(n20056,n20057,n19934);
  nor U21220(n20055,n20033,n19936);
  nand U21221(n20053,n20058,n19924);
  nand U21222(n20052,n19904,n20059);
  nand U21223(n20051,n20060,n19922);
  nand U21224(n20049,G36055,n19906);
  nand U21225(G1778,n20061,n20062);
  nand U21226(n20062,n19898,n19842);
  nand U21227(n19842,n20063,n20064,n20065,n20066);
  nor U21228(n20066,n20067,n20068);
  nor U21229(n20068,n20069,n19934);
  nor U21230(n20067,n20045,n19936);
  nand U21231(n20065,n20070,n19924);
  nand U21232(n20064,n19904,n20071);
  nand U21233(n20063,n20072,n19922);
  nand U21234(n20061,G36054,n19906);
  nand U21235(G1775,n20073,n20074);
  nand U21236(n20074,n19898,n19845);
  nand U21237(n19845,n20075,n20076,n20077,n20078);
  nor U21238(n20078,n20079,n20080);
  nor U21239(n20080,n20081,n19934);
  nor U21240(n20079,n20057,n19936);
  nand U21241(n20077,n20082,n19924);
  nand U21242(n20076,n19904,n20083);
  nand U21243(n20075,n20084,n19922);
  nand U21244(n20073,G36053,n19906);
  nand U21245(G1772,n20085,n20086);
  nand U21246(n20086,n19898,n19848);
  nand U21247(n19848,n20087,n20088,n20089,n20090);
  nor U21248(n20090,n20091,n20092);
  nor U21249(n20092,n20093,n19934);
  nor U21250(n20091,n20069,n19936);
  nand U21251(n20089,n20094,n19924);
  nand U21252(n20088,n19904,n20095);
  nand U21253(n20087,n20096,n19922);
  nand U21254(n20085,G36052,n19906);
  nand U21255(G1769,n20097,n20098);
  nand U21256(n20098,n19898,n19851);
  nand U21257(n19851,n20099,n20100,n20101,n20102);
  nor U21258(n20102,n20103,n20104);
  nor U21259(n20104,n20105,n19934);
  nor U21260(n20103,n20081,n19936);
  nand U21261(n20101,n20106,n19924);
  nand U21262(n20100,n19904,n20107);
  nand U21263(n20099,n20108,n19922);
  nand U21264(n20097,G36051,n19906);
  nand U21265(G1766,n20109,n20110);
  nand U21266(n20110,n19898,n19854);
  nand U21267(n19854,n20111,n20112,n20113,n20114);
  nor U21268(n20114,n20115,n20116);
  nor U21269(n20116,n20117,n19934);
  nor U21270(n20115,n20093,n19936);
  nand U21271(n20113,n20118,n19924);
  nand U21272(n20112,n19904,n20119);
  nand U21273(n20111,n20120,n19922);
  nand U21274(n20109,G36050,n19906);
  nand U21275(G1763,n20121,n20122);
  nand U21276(n20122,n19898,n19857);
  nand U21277(n19857,n20123,n20124,n20125,n20126);
  nor U21278(n20126,n20127,n20128);
  nor U21279(n20128,n20129,n19934);
  nor U21280(n20127,n20105,n19936);
  nand U21281(n20125,n20130,n19924);
  nand U21282(n20124,n19904,n20131);
  nand U21283(n20123,n20132,n19922);
  nand U21284(n20121,G36049,n19906);
  nand U21285(G1760,n20133,n20134);
  nand U21286(n20134,n19898,n19860);
  nand U21287(n19860,n20135,n20136,n20137,n20138);
  nor U21288(n20138,n20139,n20140);
  nor U21289(n20140,n20141,n19934);
  nor U21290(n20139,n20117,n19936);
  nand U21291(n20137,n20142,n19924);
  nand U21292(n20136,n19904,n20143);
  nand U21293(n20135,n20144,n19922);
  nand U21294(n20133,G36048,n19906);
  nand U21295(G1757,n20145,n20146);
  nand U21296(n20146,n19898,n19863);
  nand U21297(n19863,n20147,n20148,n20149,n20150);
  nor U21298(n20150,n20151,n20152);
  nor U21299(n20152,n20153,n19934);
  nor U21300(n20151,n20129,n19936);
  nand U21301(n20149,n20154,n19924);
  nand U21302(n20148,n19904,n20155);
  nand U21303(n20147,n20156,n19922);
  nand U21304(n20145,G36047,n19906);
  nand U21305(G1754,n20157,n20158);
  nand U21306(n20158,n19898,n19866);
  nand U21307(n19866,n20159,n20160,n20161,n20162);
  nor U21308(n20162,n20163,n20164);
  nor U21309(n20164,n20165,n19934);
  nor U21310(n20163,n20141,n19936);
  nand U21311(n20161,n20166,n19924);
  nand U21312(n20160,n19904,n20167);
  nand U21313(n20159,n20168,n19922);
  nand U21314(n20157,G36046,n19906);
  nand U21315(G1751,n20169,n20170);
  nand U21316(n20170,n19898,n19869);
  nand U21317(n19869,n20171,n20172,n20173,n20174);
  nor U21318(n20174,n20175,n20176);
  nor U21319(n20176,n20177,n19934);
  nor U21320(n20175,n20153,n19936);
  nand U21321(n20173,n20178,n19924);
  nand U21322(n20172,n19904,n20179);
  nand U21323(n20171,n20180,n19922);
  nand U21324(n20169,G36045,n19906);
  nand U21325(G1748,n20181,n20182);
  nand U21326(n20182,n19898,n19872);
  nand U21327(n19872,n20183,n20184,n20185,n20186);
  nor U21328(n20186,n20187,n20188);
  nor U21329(n20188,n20189,n19934);
  nor U21330(n20187,n20165,n19936);
  nand U21331(n20185,n20190,n19924);
  nand U21332(n20184,n19904,n20191);
  nand U21333(n20183,n20192,n19922);
  nand U21334(n20181,G36044,n19906);
  nand U21335(G1745,n20193,n20194);
  nand U21336(n20194,n19898,n19875);
  nand U21337(n19875,n20195,n20196,n20197,n20198);
  nor U21338(n20198,n20199,n20200);
  nor U21339(n20200,n20201,n19934);
  nor U21340(n20199,n20177,n19936);
  nand U21341(n20197,n20202,n19924);
  nand U21342(n20196,n19904,n20203);
  nand U21343(n20195,n20204,n19922);
  nand U21344(n20193,G36043,n19906);
  nand U21345(G1742,n20205,n20206);
  nand U21346(n20206,n19898,n19878);
  nand U21347(n19878,n20207,n20208,n20209,n20210);
  nor U21348(n20210,n20211,n20212);
  nor U21349(n20212,n20213,n19934);
  nor U21350(n20211,n20189,n19936);
  nand U21351(n20209,n20214,n19924);
  nand U21352(n20208,n19904,n20215);
  nand U21353(n20207,n20216,n19922);
  nand U21354(n20205,G36042,n19906);
  nand U21355(G1739,n20217,n20218);
  nand U21356(n20218,n19898,n19881);
  nand U21357(n19881,n20219,n20220,n20221,n20222);
  nor U21358(n20222,n20223,n20224);
  nor U21359(n20224,n20225,n19934);
  nor U21360(n20223,n20201,n19936);
  nand U21361(n20221,n20226,n19924);
  nand U21362(n20220,n19904,n20227);
  nand U21363(n20219,n20228,n19922);
  nand U21364(n20217,G36041,n19906);
  nand U21365(G1736,n20229,n20230);
  nand U21366(n20230,n19898,n19884);
  nand U21367(n19884,n20231,n20232,n20233,n20234);
  nor U21368(n20234,n20235,n20236);
  nor U21369(n20236,n20237,n19934);
  nor U21370(n20235,n20213,n19936);
  nand U21371(n20233,n20238,n19924);
  nand U21372(n20232,n19904,n20239);
  nand U21373(n20231,n20240,n19922);
  nand U21374(n20229,G36040,n19906);
  nand U21375(G1733,n20241,n20242);
  nand U21376(n20242,n19898,n19887);
  nand U21377(n19887,n20243,n20244,n20245,n20246);
  nor U21378(n20246,n20247,n20248);
  nor U21379(n20248,n20249,n19934);
  nor U21380(n20247,n20225,n19936);
  nand U21381(n20245,n20250,n19924);
  nand U21382(n20244,n19904,n20251);
  nand U21383(n20243,n20252,n19922);
  nand U21384(n20241,G36039,n19906);
  nand U21385(G1730,n20253,n20254);
  nand U21386(n20254,n19898,n19890);
  nand U21387(n19890,n20255,n20256,n20257,n20258);
  nor U21388(n20258,n20259,n20260);
  nor U21389(n20260,n20261,n19934);
  nor U21390(n20259,n20237,n19936);
  nand U21391(n20257,n19786,n19924);
  nand U21392(n20256,n19795,n19904);
  nand U21393(n20255,n19793,n19922);
  nand U21394(n20253,G36038,n19906);
  nand U21395(G1727,n20262,n20263);
  nand U21396(n20263,n19898,n19893);
  nand U21397(n19893,n20264,n20265,n20266,n20267);
  nand U21398(n20267,n19904,n20268);
  nand U21399(n20266,n20271,n19922);
  or U21400(n19922,n19903,n20272);
  nand U21401(n20265,n20273,n19924);
  nand U21402(n19924,n20274,n20275);
  nand U21403(n20275,n20276,n20277);
  nand U21404(n20264,n20278,n19768);
  nand U21405(n20262,G36037,n19906);
  nand U21406(n19895,n20280,n20281,n20282);
  nand U21407(n20280,n20283,n20284,n20285);
  nand U21408(n20285,n20286,n20287);
  nand U21409(G1716,n20288,n20289);
  nand U21410(n20289,G36006,n20290);
  nand U21411(n20288,n20291,n20292);
  nand U21412(G1715,n20293,n20294);
  nand U21413(n20294,n20291,n20295);
  nand U21414(n20293,G36005,n20290);
  nand U21415(G1549,n20296,n20297,n20298,n20299);
  nor U21416(n20299,n20300,n20301,n20302,n20303);
  nor U21417(n20303,n20189,n20304);
  nor U21418(n20302,n20165,n20305);
  nor U21419(n20301,n20306,n20307);
  not U21420(n20307,n20308);
  nor U21421(n20300,n20309,n20310);
  nand U21422(n20298,G36214,G1406);
  nand U21423(n20297,n20311,n20190);
  nand U21424(n20296,n20312,n20192);
  nand U21425(G1548,n20313,n20314,n20315,n20316);
  nor U21426(n20316,n20317,n20318,n20319,n20320);
  nor U21427(n20320,n19948,n20304);
  nor U21428(n20319,n19949,n20305);
  nor U21429(n20318,n20306,n20321);
  nor U21430(n20317,n20322,n20310);
  nand U21431(n20315,G36213,G1406);
  nand U21432(n20314,n20311,n19950);
  nand U21433(n20313,n20312,n19952);
  nand U21434(G1547,n20323,n20324,n20325,n20326);
  nor U21435(n20326,n20327,n20328,n20329,n20330);
  nor U21436(n20330,n20105,n20304);
  nor U21437(n20329,n20081,n20305);
  nor U21438(n20328,n20306,n20331);
  nor U21439(n20327,n20332,n20310);
  nand U21440(n20325,G36212,G1406);
  nand U21441(n20324,n20311,n20106);
  nand U21442(n20323,n20312,n20108);
  nand U21443(G1546,n20333,n20334,n20335,n20336);
  nor U21444(n20336,n20337,n20338,n20339,n20340);
  nor U21445(n20340,n19997,n20304);
  nor U21446(n20339,n19973,n20305);
  nor U21447(n20338,n20306,n20341);
  nor U21448(n20337,n20342,n20310);
  nand U21449(n20335,G36211,G1406);
  nand U21450(n20334,n20311,n19998);
  nand U21451(n20333,n20312,n20000);
  nand U21452(G1545,n20343,n20344,n20345,n20346);
  nor U21453(n20346,n20347,n20348,n20349,n20350);
  nor U21454(n20350,n20153,n20304);
  nor U21455(n20349,n20129,n20305);
  nor U21456(n20348,n20306,n20351);
  not U21457(n20351,n20352);
  nor U21458(n20347,n20353,n20310);
  nand U21459(n20345,G36210,G1406);
  nand U21460(n20344,n20311,n20154);
  nand U21461(n20343,n20312,n20156);
  nand U21462(G1544,n20354,n20355,n20356,n20357);
  nor U21463(n20357,n20358,n20359,n20360,n20361);
  nor U21464(n20361,n20362,n20363);
  nor U21465(n20360,n20364,n20365);
  nor U21466(n20359,G36209,n20306);
  nand U21467(n20356,n20366,n19765);
  or U21468(n20355,n20310,n20367);
  or U21469(n20354,n20305,n20213);
  nand U21470(G1543,n20368,n20369,n20370,n20371);
  nor U21471(n20371,n20372,n20373,n20374,n20375);
  nor U21472(n20375,n20045,n20304);
  nor U21473(n20374,n20021,n20305);
  nor U21474(n20373,n20306,n20376);
  nor U21475(n20372,n20377,n20310);
  nand U21476(n20370,G36208,G1406);
  nand U21477(n20369,n20311,n20046);
  nand U21478(n20368,n20312,n20048);
  nand U21479(G1542,n20378,n20379,n20380,n20381);
  nor U21480(n20381,n20382,n20383,n20384,n20385);
  nor U21481(n20385,n19933,n20304);
  nor U21482(n20384,n19935,n20305);
  nor U21483(n20383,n20306,n20386);
  not U21484(n20386,n20387);
  nor U21485(n20382,n20388,n20310);
  nand U21486(n20380,G36207,G1406);
  nand U21487(n20379,n20311,n19937);
  nand U21488(n20378,n20312,n19939);
  nand U21489(G1541,n20389,n20390,n20391,n20392);
  nor U21490(n20392,n20393,n20394,n20395,n20396);
  nor U21491(n20396,n20177,n20304);
  nor U21492(n20395,n20153,n20305);
  nor U21493(n20394,n20306,n20397);
  nor U21494(n20393,n20398,n20310);
  nand U21495(n20391,G36206,G1406);
  nand U21496(n20390,n20311,n20178);
  nand U21497(n20389,n20312,n20180);
  nand U21498(G1540,n20399,n20400,n20401,n20402);
  nor U21499(n20402,n20403,n20404,n20405);
  nor U21500(n20405,n20406,n20310);
  nor U21501(n20404,n20407,n19780);
  nor U21502(n20403,n20237,n20305);
  nand U21503(n20401,n20312,n19793);
  nand U21504(n20400,n20366,n19771);
  nand U21505(n20399,n20311,n19786);
  nand U21506(G1539,n20408,n20409,n20410,n20411);
  nor U21507(n20411,n20412,n20413,n20414,n20415);
  nor U21508(n20415,n20021,n20304);
  nor U21509(n20414,n19997,n20305);
  nor U21510(n20413,n20306,n20416);
  nor U21511(n20412,n20417,n20310);
  nand U21512(n20410,G36204,G1406);
  nand U21513(n20409,n20311,n20022);
  nand U21514(n20408,n20312,n20024);
  nand U21515(G1538,n20418,n20419,n20420,n20421);
  nor U21516(n20421,n20422,n20423,n20424,n20425);
  nor U21517(n20425,n20129,n20304);
  nor U21518(n20424,n20105,n20305);
  nor U21519(n20423,n20306,n20426);
  nor U21520(n20422,n20427,n20310);
  nand U21521(n20420,G36203,G1406);
  nand U21522(n20419,n20311,n20130);
  nand U21523(n20418,n20312,n20132);
  nand U21524(G1537,n20428,n20429,n20430,n20431);
  nor U21525(n20431,n20432,n20433,n20434,n20435);
  nor U21526(n20435,n19973,n20304);
  nor U21527(n20434,n19948,n20305);
  nor U21528(n20433,n20306,n20436);
  not U21529(n20436,n20437);
  nor U21530(n20432,n20438,n20310);
  nand U21531(n20430,G36202,G1406);
  nand U21532(n20429,n20311,n19974);
  nand U21533(n20428,n20312,n19976);
  nand U21534(G1536,n20439,n20440,n20441,n20442);
  nor U21535(n20442,n20443,n20444,n20445,n20446);
  nor U21536(n20446,n20081,n20304);
  nor U21537(n20445,n20057,n20305);
  nor U21538(n20444,n20306,n20447);
  nor U21539(n20443,n20448,n20310);
  nand U21540(n20441,G36201,G1406);
  nand U21541(n20440,n20311,n20082);
  nand U21542(n20439,n20312,n20084);
  nand U21543(G1535,n20449,n20450,n20451,n20452);
  nor U21544(n20452,n20453,n20454,n20455,n20456);
  nor U21545(n20456,n20213,n20304);
  nor U21546(n20455,n20189,n20305);
  nor U21547(n20454,n20306,n20457);
  nor U21548(n20453,n20458,n20310);
  nand U21549(n20451,G36200,G1406);
  nand U21550(n20450,n20311,n20214);
  nand U21551(n20449,n20312,n20216);
  nand U21552(G1534,n20459,n20460,n20461,n20462);
  nor U21553(n20462,n20463,n20464,n20465,n20466);
  nor U21554(n20466,n20069,n20304);
  nor U21555(n20465,n20045,n20305);
  nor U21556(n20464,n20306,n20467);
  nor U21557(n20463,n20468,n20310);
  nand U21558(n20461,G36199,G1406);
  nand U21559(n20460,n20311,n20070);
  nand U21560(n20459,n20312,n20072);
  nand U21561(G1533,n20469,n20470,n20471,n20472);
  nor U21562(n20472,n20473,n20474,n20475,n20476);
  nor U21563(n20476,n19985,n20304);
  nor U21564(n20475,n19961,n20305);
  nor U21565(n20474,n20306,n20477);
  nor U21566(n20473,n20478,n20310);
  nand U21567(n20471,G36198,G1406);
  nand U21568(n20470,n20311,n19986);
  nand U21569(n20469,n20312,n19988);
  nand U21570(G1532,n20479,n20480,n20481,n20482);
  nor U21571(n20482,n20483,n20484,n20485,n20486);
  nor U21572(n20486,n20225,n20304);
  nor U21573(n20485,n20201,n20305);
  nor U21574(n20484,n20487,n20310);
  nor U21575(n20483,n20306,n20488);
  nand U21576(n20480,n20311,n20226);
  nand U21577(n20479,n20312,n20228);
  nand U21578(G1531,n20489,n20490,n20491,n20492);
  nor U21579(n20492,n20493,n20494,n20495,n20496);
  nor U21580(n20496,n20165,n20304);
  nor U21581(n20495,n20141,n20305);
  nor U21582(n20494,n20306,n20497);
  nor U21583(n20493,n20498,n20310);
  nand U21584(n20491,G36196,G1406);
  nand U21585(n20490,n20311,n20166);
  nand U21586(n20489,n20312,n20168);
  nand U21587(G1530,n20499,n20500,n20501);
  nor U21588(n20501,n20502,n20503,n20504);
  nor U21589(n20504,n20505,n20310);
  nor U21590(n20503,n20407,n20506);
  nor U21591(n20502,n20249,n20305);
  nand U21592(n20500,n20311,n20273);
  nand U21593(n20499,n20312,n20271);
  nand U21594(G1529,n20507,n20508,n20509,n20510);
  nor U21595(n20510,n20511,n20512,n20513,n20514);
  nor U21596(n20514,n20033,n20304);
  nor U21597(n20513,n20009,n20305);
  nor U21598(n20512,n20306,n20515);
  not U21599(n20515,n20516);
  nor U21600(n20511,n20517,n20310);
  nand U21601(n20509,G36194,G1406);
  nand U21602(n20508,n20311,n20034);
  nand U21603(n20507,n20312,n20036);
  nand U21604(G1528,n20518,n20519,n20520,n20521);
  nor U21605(n20521,n20522,n20523,n20524,n20525);
  nor U21606(n20525,n20117,n20304);
  nor U21607(n20524,n20093,n20305);
  nor U21608(n20523,n20306,n20526);
  nor U21609(n20522,n20527,n20310);
  nand U21610(n20520,G36193,G1406);
  nand U21611(n20519,n20311,n20118);
  nand U21612(n20518,n20312,n20120);
  nand U21613(G1527,n20528,n20529,n20530,n20531);
  nor U21614(n20531,n20532,n20533,n20534,n20535);
  nor U21615(n20535,n20009,n20304);
  nor U21616(n20534,n19985,n20305);
  nor U21617(n20533,n20306,n20536);
  nor U21618(n20532,n20537,n20310);
  nand U21619(n20530,G36192,G1406);
  nand U21620(n20529,n20311,n20010);
  nand U21621(n20528,n20312,n20012);
  nand U21622(G1526,n20538,n20539,n20540,n20541);
  nor U21623(n20541,n20542,n20543,n20544,n20545);
  nor U21624(n20545,n20141,n20304);
  nor U21625(n20544,n20117,n20305);
  nor U21626(n20543,n20306,n20546);
  nor U21627(n20542,n20547,n20310);
  nand U21628(n20540,G36191,G1406);
  nand U21629(G1525,n20548,n20549,n20550,n20551);
  nor U21630(n20551,n20552,n20553,n20554);
  nor U21631(n20554,n20555,n20310);
  nor U21632(n20553,n20407,n20556);
  not U21633(n20556,G36190);
  and U21634(n20407,n20306,G36215);
  nor U21635(n20552,n20225,n20305);
  nand U21636(n20550,n20312,n20252);
  nand U21637(n20549,n20366,n19768);
  not U21638(n20366,n20304);
  nand U21639(n20548,n20311,n20250);
  nand U21640(G1524,n20557,n20558,n20559,n20560);
  nor U21641(n20560,n20561,n20562,n20563,n20564);
  nor U21642(n20564,n20057,n20304);
  nor U21643(n20563,n20033,n20305);
  nor U21644(n20562,n20306,n20565);
  nor U21645(n20561,n20566,n20310);
  nand U21646(n20559,G36189,G1406);
  nand U21647(n20558,n20311,n20058);
  nand U21648(n20557,n20312,n20060);
  nand U21649(G1523,n20567,n20568,n20569,n20570);
  nor U21650(n20570,n20571,n20572,n20573,n20574);
  nor U21651(n20574,n20201,n20304);
  nor U21652(n20573,n20177,n20305);
  nor U21653(n20572,n20306,n20575);
  nor U21654(n20571,n20576,n20310);
  nand U21655(n20569,G36188,G1406);
  nand U21656(n20568,n20311,n20202);
  nand U21657(n20567,n20312,n20204);
  nand U21658(G1522,n20577,n20578,n20579,n20580);
  nor U21659(n20580,n20581,n20582,n20583,n20584);
  nor U21660(n20584,n19961,n20304);
  nor U21661(n20583,n19933,n20305);
  nor U21662(n20582,n20306,n20585);
  nor U21663(n20581,n20586,n20310);
  nand U21664(n20579,G36187,G1406);
  nand U21665(n20578,n20311,n19962);
  nand U21666(n20577,n20312,n19964);
  nand U21667(G1521,n20587,n20588,n20589,n20590);
  nor U21668(n20590,n20591,n20592,n20593,n20594);
  nor U21669(n20594,n20093,n20304);
  nand U21670(n20304,n20595,n20596,n20597);
  nor U21671(n20593,n20069,n20305);
  nand U21672(n20305,n20595,n20598,n20597);
  nor U21673(n20592,n20306,n20599);
  and U21674(n20306,n20600,n20601,n20602,n19677);
  nand U21675(n20601,n20282,n20603);
  nand U21676(n20603,n20604,n20605);
  or U21677(n20604,n20595,n20606);
  nor U21678(n20606,n20607,n20608,n20609);
  nand U21679(n20600,n20597,n20610);
  and U21680(n20597,n20611,n20282,n20612);
  nor U21681(n20591,n20613,n20310);
  nand U21682(n20310,n20282,n20614);
  nand U21683(n20614,n20615,n20616);
  nand U21684(n20616,n20595,n20608);
  nand U21685(n20589,G36186,G1406);
  nand U21686(n20588,n20311,n20094);
  not U21687(n20311,n20365);
  nand U21688(n20365,n20282,n20607,n20595);
  nand U21689(n20607,n20617,n20618);
  nand U21690(n20618,n20277,n20619);
  nand U21691(n20619,n20620,n20621);
  nand U21692(n20587,n20312,n20096);
  not U21693(n20312,n20363);
  nand U21694(n20363,n20282,n20609,n20595);
  not U21695(n20595,n20610);
  nand U21696(n20610,n20622,n20281);
  nand U21697(n20609,n20623,n20624);
  nand U21698(n20624,n20272,n20625);
  nand U21699(G1520,n20626,n20627);
  nand U21700(n20627,n20628,G36215,n20629);
  nand U21701(n20628,n20630,n20631,n20632,n20633);
  nand U21702(n20633,n20634,n20635);
  nand U21703(n20634,n20636,n20637);
  nand U21704(n20637,n20638,n20639);
  nand U21705(n20638,n20287,n20640);
  nand U21706(n20640,n20277,n20641);
  or U21707(n20636,n20642,n20284);
  nand U21708(n20632,n20643,n20642,n20644);
  nand U21709(n20642,n20645,n20646,n20647,n20648);
  nor U21710(n20648,n20649,n20650,n20651,n20652);
  nand U21711(n20652,n20653,n20654,n20655,n20656);
  xor U21712(n20656,n19759,n20487);
  xor U21713(n20655,n19762,n20367);
  xor U21714(n20654,n19765,n20555);
  xor U21715(n20653,n20261,n20268);
  not U21716(n20261,n19771);
  nand U21717(n20651,n20657,n20658,n20659,n20660);
  xor U21718(n20660,n19747,n20398);
  xor U21719(n20659,n19750,n20309);
  xor U21720(n20658,n19753,n20576);
  xor U21721(n20657,n19756,n20458);
  nand U21722(n20650,n20661,n20662,n20663,n20664);
  xor U21723(n20664,n20131,n20117);
  xor U21724(n20663,n20143,n20129);
  xor U21725(n20662,n20155,n20141);
  xor U21726(n20661,n19744,n20498);
  nand U21727(n20649,n20665,n20666,n20667,n20668);
  xor U21728(n20668,n20083,n20069);
  xor U21729(n20667,n20095,n20081);
  xor U21730(n20666,n20107,n20093);
  xor U21731(n20665,n20119,n20105);
  nor U21732(n20647,n20669,n20670,n20671,n20672);
  xor U21733(n20672,n19684,n19920);
  xor U21734(n20671,n19681,n19911);
  nand U21735(n20670,n20673,n20674,n20675);
  xor U21736(n20675,n20249,n19795);
  nand U21737(n20669,n20676,n20677,n20678,n20679);
  xor U21738(n20679,n19938,n19949);
  xor U21739(n20678,n19951,n19933);
  xor U21740(n20677,n19963,n19948);
  xor U21741(n20676,n19975,n19961);
  nor U21742(n20646,n20680,n20681,n20682,n20683);
  xor U21743(n20683,n19708,n20023);
  xor U21744(n20682,n19705,n20011);
  xor U21745(n20681,n19702,n19999);
  xor U21746(n20680,n19699,n19987);
  nor U21747(n20645,n20684,n20685,n20686,n20687);
  xor U21748(n20687,n19720,n20071);
  xor U21749(n20686,n19717,n20059);
  xor U21750(n20685,n19714,n20047);
  xor U21751(n20684,n19711,n20035);
  nand U21752(n20631,n20688,n20689,n20272);
  nand U21753(n20689,n20673,n20690);
  nand U21754(n20690,n20691,n20674);
  or U21755(n20674,n19905,n20692);
  nand U21756(n20691,n20693,n20694);
  nand U21757(n20694,n20639,n19681,n20695);
  not U21758(n20695,n19911);
  nand U21759(n20693,n20696,n20697,n20698);
  nand U21760(n20698,n20699,n19911);
  nand U21761(n20699,n19681,n20639);
  nand U21762(n20697,n20700,n20701,n20702);
  nand U21763(n20702,n20388,n19939);
  not U21764(n19939,n20703);
  nand U21765(n20701,n20704,n20705,n20706);
  nand U21766(n20706,n20707,n19951);
  nand U21767(n20705,n20708,n20709,n20710);
  nand U21768(n20710,n20586,n19964);
  not U21769(n19964,n20711);
  nand U21770(n20709,n20712,n20713,n20714);
  nand U21771(n20714,n20715,n19975);
  nand U21772(n20713,n20716,n20717,n20718);
  nand U21773(n20718,n20478,n19988);
  not U21774(n19988,n20719);
  nand U21775(n20717,n20720,n20721,n20722);
  nand U21776(n20722,n20723,n19999);
  nand U21777(n20721,n20724,n20725,n20726);
  nand U21778(n20726,n20537,n20012);
  not U21779(n20012,n20727);
  nand U21780(n20725,n20728,n20729,n20730);
  nand U21781(n20730,n20731,n20023);
  nand U21782(n20729,n20732,n20733,n20734);
  nand U21783(n20734,n20517,n20036);
  not U21784(n20036,n20735);
  nand U21785(n20733,n20736,n20737,n20738);
  nand U21786(n20738,n20739,n20047);
  nand U21787(n20737,n20740,n20741,n20742);
  nand U21788(n20742,n20566,n20060);
  not U21789(n20060,n20743);
  nand U21790(n20741,n20744,n20745,n20746);
  nand U21791(n20746,n20747,n20071);
  nand U21792(n20745,n20748,n20749,n20750);
  nand U21793(n20750,n20448,n20084);
  not U21794(n20084,n20751);
  nand U21795(n20749,n20752,n20753,n20754);
  nand U21796(n20754,n20755,n20095);
  nand U21797(n20753,n20756,n20757,n20758);
  nand U21798(n20758,n20332,n20108);
  not U21799(n20108,n20759);
  nand U21800(n20757,n20760,n20761,n20762);
  nand U21801(n20762,n20763,n20119);
  nand U21802(n20761,n20764,n20765,n20766);
  nand U21803(n20766,n20132,n19735,n20427);
  not U21804(n20132,n20767);
  nand U21805(n20765,n20768,n20769,n20770);
  nand U21806(n20770,n20771,n20143,n20129);
  nand U21807(n20769,n20772,n20773,n20774);
  nand U21808(n20774,n20156,n19741,n20353);
  not U21809(n20156,n20775);
  nand U21810(n20773,n20776,n20777,n20778);
  nand U21811(n20778,n20779,n20167,n20153);
  nand U21812(n20777,n20780,n20781,n20782);
  nand U21813(n20782,n20180,n19747,n20398);
  not U21814(n20180,n20783);
  nand U21815(n20781,n20784,n20785,n20786);
  nand U21816(n20786,n20787,n20191,n20177);
  nand U21817(n20785,n20788,n20789,n20790);
  nand U21818(n20790,n20204,n19753,n20576);
  not U21819(n20204,n20791);
  nand U21820(n20789,n20792,n20793,n20794);
  nand U21821(n20794,n20795,n20215,n20201);
  nand U21822(n20793,n20796,n20797,n20798);
  nand U21823(n20798,n20228,n19759,n20487);
  not U21824(n20228,n20799);
  nand U21825(n20797,n20800,n20801,n20802);
  nand U21826(n20802,n20362,n20239,n20225);
  nand U21827(n20801,n20803,n20804,n20805);
  nand U21828(n20805,n20252,n19765,n20555);
  not U21829(n20252,n20806);
  nand U21830(n20804,n20807,n20808,n20809);
  nand U21831(n20809,n20806,n20251,n20237);
  not U21832(n20237,n19765);
  nand U21833(n20808,n20810,n20268,n20811);
  nand U21834(n20811,n20271,n19771);
  nand U21835(n20810,n20812,n20406);
  nand U21836(n20812,n20249,n20813);
  nand U21837(n20807,n19795,n20813,n20249);
  not U21838(n20249,n19768);
  not U21839(n20813,n19793);
  xor U21840(n19793,n20814,n20815);
  nand U21841(n20814,n20816,n20817,n20818);
  nand U21842(n20818,n20819,n19768);
  nand U21843(n20803,n20240,n19762,n20367);
  not U21844(n20240,n20362);
  nand U21845(n20800,n20799,n20227,n20213);
  nand U21846(n20796,n20216,n19756,n20458);
  not U21847(n20216,n20795);
  nand U21848(n20792,n20791,n20203,n20189);
  nand U21849(n20788,n20192,n19750,n20309);
  not U21850(n20192,n20787);
  nand U21851(n20784,n20783,n20179,n20165);
  nand U21852(n20780,n20168,n19744,n20498);
  not U21853(n20168,n20779);
  nand U21854(n20776,n20775,n20155,n20141);
  nand U21855(n20772,n20144,n19738,n20547);
  not U21856(n20144,n20771);
  nand U21857(n20768,n20767,n20131,n20117);
  nand U21858(n20764,n20527,n20120);
  not U21859(n20120,n20763);
  nand U21860(n20760,n20759,n20107);
  nand U21861(n20756,n20613,n20096);
  not U21862(n20096,n20755);
  nand U21863(n20752,n20751,n20083);
  nand U21864(n20748,n20468,n20072);
  not U21865(n20072,n20747);
  nand U21866(n20744,n20743,n20059);
  nand U21867(n20740,n20377,n20048);
  not U21868(n20048,n20739);
  nand U21869(n20736,n20735,n20035);
  nand U21870(n20732,n20417,n20024);
  not U21871(n20024,n20731);
  nand U21872(n20728,n20727,n20011);
  nand U21873(n20724,n20342,n20000);
  not U21874(n20000,n20723);
  nand U21875(n20720,n20719,n19987);
  nand U21876(n20716,n20438,n19976);
  not U21877(n19976,n20715);
  nand U21878(n20712,n20711,n19963);
  nand U21879(n20708,n20322,n19952);
  not U21880(n19952,n20707);
  nand U21881(n20704,n20703,n19938);
  nand U21882(n20700,n20820,n19921);
  or U21883(n20696,n19921,n20820);
  nand U21884(n20673,n20692,n19905);
  nor U21885(n20630,n20821,n20822);
  and U21886(n20822,n20639,n20625,n20276);
  nor U21887(n20821,n20823,n20639);
  nand U21888(n20639,n20824,n20825);
  nand U21889(n20825,n20826,n20827);
  nand U21890(n20824,n20828,n20829,n20830);
  nand U21891(n20830,n20831,n20832);
  nand U21892(n20829,n20833,n20834,n20835);
  or U21893(n20835,n20832,n20831);
  and U21894(n20831,n20836,n20837);
  nand U21895(n20837,n19911,n20838);
  nand U21896(n20836,n20839,n19681);
  nand U21897(n20832,n20840,n20841,n20842);
  nand U21898(n20842,n20843,n19911);
  nand U21899(n20841,n20844,n20845);
  nand U21900(n20840,n20846,n19681);
  nand U21901(n20834,n20847,n20848,n20849);
  nand U21902(n20849,n20850,n20851);
  nand U21903(n20848,n20852,n20853,n20854,n20855);
  or U21904(n20855,n20851,n20850);
  and U21905(n20850,n20856,n20857);
  nand U21906(n20857,n20858,n20859);
  nand U21907(n20856,n20860,n20861,n20862);
  or U21908(n20862,n20859,n20858);
  and U21909(n20858,n20863,n20864,n20865);
  nand U21910(n20865,n20843,n19951);
  nand U21911(n20864,n20844,n19950);
  nand U21912(n20863,n20846,n19690);
  nand U21913(n20859,n20866,n20867,n20868);
  nand U21914(n20868,n20839,n19690);
  nand U21915(n20867,n19950,n20869);
  nand U21916(n20866,n19951,n20838);
  nand U21917(n20861,n20870,n20871,n20872);
  nand U21918(n20870,n20873,n19962);
  nand U21919(n20860,n20874,n20875,n20876);
  nand U21920(n20876,n20877,n20878);
  nand U21921(n20878,n20872,n20879);
  nand U21922(n20879,n19962,n20869);
  and U21923(n20872,n20880,n20881);
  nand U21924(n20881,n19963,n20838);
  nand U21925(n20880,n20839,n19693);
  not U21926(n20877,n20871);
  nand U21927(n20871,n20882,n20883,n20884);
  nand U21928(n20884,n20843,n19963);
  nand U21929(n20883,n20844,n19962);
  nand U21930(n20882,n20846,n19693);
  nand U21931(n20875,n20885,n20886);
  nand U21932(n20874,n20887,n20888,n20889);
  or U21933(n20889,n20886,n20885);
  and U21934(n20885,n20890,n20891,n20892);
  nand U21935(n20892,n20843,n19975);
  nand U21936(n20891,n20844,n19974);
  nand U21937(n20890,n20846,n19696);
  nand U21938(n20886,n20893,n20894,n20895);
  nand U21939(n20895,n20839,n19696);
  nand U21940(n20894,n19974,n20869);
  nand U21941(n20893,n19975,n20838);
  nand U21942(n20888,n20896,n20897,n20898);
  nand U21943(n20896,n20873,n19986);
  nand U21944(n20887,n20899,n20900,n20901);
  nand U21945(n20901,n20902,n20903);
  nand U21946(n20903,n20898,n20904);
  nand U21947(n20904,n19986,n20869);
  and U21948(n20898,n20905,n20906);
  nand U21949(n20906,n19987,n20838);
  nand U21950(n20905,n20839,n19699);
  not U21951(n20902,n20897);
  nand U21952(n20897,n20907,n20908,n20909);
  nand U21953(n20909,n20843,n19987);
  nand U21954(n20908,n20844,n19986);
  nand U21955(n20907,n20846,n19699);
  nand U21956(n20900,n20910,n20911);
  nand U21957(n20899,n20912,n20913,n20914);
  or U21958(n20914,n20911,n20910);
  and U21959(n20910,n20915,n20916,n20917);
  nand U21960(n20917,n20843,n19999);
  nand U21961(n20916,n20844,n19998);
  nand U21962(n20915,n20846,n19702);
  nand U21963(n20911,n20918,n20919,n20920);
  nand U21964(n20920,n20839,n19702);
  nand U21965(n20919,n19998,n20869);
  nand U21966(n20918,n19999,n20838);
  nand U21967(n20913,n20921,n20922,n20923);
  nand U21968(n20921,n20873,n20010);
  nand U21969(n20912,n20924,n20925,n20926);
  nand U21970(n20926,n20927,n20928);
  nand U21971(n20928,n20923,n20929);
  nand U21972(n20929,n20010,n20869);
  and U21973(n20923,n20930,n20931);
  nand U21974(n20931,n20011,n20838);
  nand U21975(n20930,n20839,n19705);
  not U21976(n20927,n20922);
  nand U21977(n20922,n20932,n20933,n20934);
  nand U21978(n20934,n20843,n20011);
  nand U21979(n20933,n20844,n20010);
  nand U21980(n20932,n20846,n19705);
  nand U21981(n20925,n20935,n20936);
  nand U21982(n20924,n20937,n20938,n20939);
  or U21983(n20939,n20936,n20935);
  and U21984(n20935,n20940,n20941,n20942);
  nand U21985(n20942,n20843,n20023);
  nand U21986(n20941,n20844,n20022);
  nand U21987(n20940,n20846,n19708);
  nand U21988(n20936,n20943,n20944,n20945);
  nand U21989(n20945,n20839,n19708);
  nand U21990(n20944,n20022,n20869);
  nand U21991(n20943,n20023,n20838);
  nand U21992(n20938,n20946,n20947,n20948);
  nand U21993(n20946,n20873,n20034);
  nand U21994(n20937,n20949,n20950,n20951);
  nand U21995(n20951,n20952,n20953);
  nand U21996(n20953,n20948,n20954);
  nand U21997(n20954,n20034,n20869);
  and U21998(n20948,n20955,n20956);
  nand U21999(n20956,n20035,n20838);
  nand U22000(n20955,n20839,n19711);
  not U22001(n20952,n20947);
  nand U22002(n20947,n20957,n20958,n20959);
  nand U22003(n20959,n20843,n20035);
  nand U22004(n20958,n20844,n20034);
  nand U22005(n20957,n20846,n19711);
  nand U22006(n20950,n20960,n20961);
  nand U22007(n20949,n20962,n20963,n20964);
  or U22008(n20964,n20961,n20960);
  and U22009(n20960,n20965,n20966,n20967);
  nand U22010(n20967,n20843,n20047);
  nand U22011(n20966,n20844,n20046);
  nand U22012(n20965,n20846,n19714);
  nand U22013(n20961,n20968,n20969,n20970);
  nand U22014(n20970,n20839,n19714);
  nand U22015(n20969,n20046,n20869);
  nand U22016(n20968,n20047,n20838);
  nand U22017(n20963,n20971,n20972,n20973);
  nand U22018(n20971,n20873,n20058);
  nand U22019(n20962,n20974,n20975,n20976);
  nand U22020(n20976,n20977,n20978);
  nand U22021(n20978,n20973,n20979);
  nand U22022(n20979,n20058,n20869);
  and U22023(n20973,n20980,n20981);
  nand U22024(n20981,n20059,n20838);
  nand U22025(n20980,n20839,n19717);
  not U22026(n20977,n20972);
  nand U22027(n20972,n20982,n20983,n20984);
  nand U22028(n20984,n20843,n20059);
  nand U22029(n20983,n20844,n20058);
  nand U22030(n20982,n20846,n19717);
  nand U22031(n20975,n20985,n20986);
  nand U22032(n20974,n20987,n20988,n20989);
  or U22033(n20989,n20986,n20985);
  and U22034(n20985,n20990,n20991,n20992);
  nand U22035(n20992,n20843,n20071);
  nand U22036(n20991,n20844,n20070);
  nand U22037(n20990,n20846,n19720);
  nand U22038(n20986,n20993,n20994,n20995);
  nand U22039(n20995,n20839,n19720);
  nand U22040(n20994,n20070,n20869);
  nand U22041(n20993,n20071,n20838);
  nand U22042(n20988,n20996,n20997,n20998);
  nand U22043(n20996,n20873,n20082);
  nand U22044(n20987,n20999,n21000,n21001);
  nand U22045(n21001,n21002,n21003);
  nand U22046(n21003,n20998,n21004);
  nand U22047(n21004,n20082,n20869);
  and U22048(n20998,n21005,n21006);
  nand U22049(n21006,n20083,n20838);
  nand U22050(n21005,n20839,n19723);
  not U22051(n21002,n20997);
  nand U22052(n20997,n21007,n21008,n21009);
  nand U22053(n21009,n20843,n20083);
  nand U22054(n21008,n20844,n20082);
  nand U22055(n21007,n20846,n19723);
  nand U22056(n21000,n21010,n21011);
  nand U22057(n20999,n21012,n21013,n21014);
  or U22058(n21014,n21011,n21010);
  and U22059(n21010,n21015,n21016,n21017);
  nand U22060(n21017,n20843,n20095);
  nand U22061(n21016,n20844,n20094);
  nand U22062(n21015,n20846,n19726);
  nand U22063(n21011,n21018,n21019,n21020);
  nand U22064(n21020,n20839,n19726);
  nand U22065(n21019,n20094,n20869);
  nand U22066(n21018,n20095,n20838);
  nand U22067(n21013,n21021,n21022,n21023);
  nand U22068(n21021,n20873,n20106);
  nand U22069(n21012,n21024,n21025,n21026);
  nand U22070(n21026,n21027,n21028);
  nand U22071(n21028,n21023,n21029);
  nand U22072(n21029,n20106,n20869);
  and U22073(n21023,n21030,n21031);
  nand U22074(n21031,n20107,n20838);
  nand U22075(n21030,n20839,n19729);
  not U22076(n21027,n21022);
  nand U22077(n21022,n21032,n21033,n21034);
  nand U22078(n21034,n20843,n20107);
  nand U22079(n21033,n20844,n20106);
  nand U22080(n21032,n20846,n19729);
  nand U22081(n21025,n21035,n21036);
  nand U22082(n21024,n21037,n21038,n21039);
  or U22083(n21039,n21036,n21035);
  and U22084(n21035,n21040,n21041,n21042);
  nand U22085(n21042,n20843,n20119);
  nand U22086(n21041,n20844,n20118);
  nand U22087(n21040,n20846,n19732);
  nand U22088(n21036,n21043,n21044,n21045);
  nand U22089(n21045,n20839,n19732);
  nand U22090(n21044,n20118,n20869);
  nand U22091(n21043,n20119,n20838);
  nand U22092(n21038,n21046,n21047,n21048);
  nand U22093(n21046,n20873,n20130);
  nand U22094(n21037,n21049,n21050,n21051);
  nand U22095(n21051,n21052,n21053);
  nand U22096(n21053,n21048,n21054);
  nand U22097(n21054,n20130,n20869);
  and U22098(n21048,n21055,n21056);
  nand U22099(n21056,n20131,n20838);
  nand U22100(n21055,n20839,n19735);
  not U22101(n21052,n21047);
  nand U22102(n21047,n21057,n21058,n21059);
  nand U22103(n21059,n20843,n20131);
  nand U22104(n21058,n20844,n20130);
  nand U22105(n21057,n20846,n19735);
  nand U22106(n21050,n21060,n21061);
  nand U22107(n21049,n21062,n21063,n21064);
  or U22108(n21064,n21061,n21060);
  and U22109(n21060,n21065,n21066,n21067);
  nand U22110(n21067,n20843,n20143);
  nand U22111(n21066,n20844,n20142);
  nand U22112(n21065,n20846,n19738);
  nand U22113(n21061,n21068,n21069,n21070);
  nand U22114(n21070,n20839,n19738);
  nand U22115(n21069,n20142,n20869);
  nand U22116(n21068,n20143,n20838);
  nand U22117(n21063,n21071,n21072,n21073);
  nand U22118(n21071,n20873,n20154);
  nand U22119(n21062,n21074,n21075,n21076);
  nand U22120(n21076,n21077,n21078);
  nand U22121(n21078,n21073,n21079);
  nand U22122(n21079,n20154,n20869);
  and U22123(n21073,n21080,n21081);
  nand U22124(n21081,n20155,n20838);
  nand U22125(n21080,n20839,n19741);
  not U22126(n21077,n21072);
  nand U22127(n21072,n21082,n21083,n21084);
  nand U22128(n21084,n20843,n20155);
  nand U22129(n21083,n20844,n20154);
  nand U22130(n21082,n20846,n19741);
  nand U22131(n21075,n21085,n21086);
  nand U22132(n21074,n21087,n21088,n21089);
  or U22133(n21089,n21086,n21085);
  and U22134(n21085,n21090,n21091,n21092);
  nand U22135(n21092,n20843,n20167);
  nand U22136(n21091,n20844,n20166);
  nand U22137(n21090,n20846,n19744);
  nand U22138(n21086,n21093,n21094,n21095,n21096);
  nand U22139(n21095,n20166,n20869);
  nand U22140(n21094,n20167,n20838);
  nand U22141(n21093,n20839,n19744);
  nand U22142(n21088,n21097,n21098,n21099,n21096);
  nand U22143(n21098,n20873,n20178);
  nand U22144(n21087,n21100,n21101,n21102);
  nand U22145(n21102,n21103,n21104);
  nand U22146(n21104,n21097,n21105);
  nand U22147(n21105,n20178,n20869);
  and U22148(n21097,n21106,n21107);
  nand U22149(n21107,n20179,n20838);
  nand U22150(n21106,n20839,n19747);
  not U22151(n21103,n21099);
  nand U22152(n21099,n21108,n21109,n21110);
  nand U22153(n21110,n20843,n20179);
  nand U22154(n21109,n20844,n20178);
  nand U22155(n21108,n20846,n19747);
  nand U22156(n21101,n21111,n21112);
  nand U22157(n21100,n21113,n21114,n21115);
  or U22158(n21115,n21112,n21111);
  and U22159(n21111,n21116,n21117,n21118);
  nand U22160(n21118,n20843,n20191);
  nand U22161(n21117,n20844,n20190);
  nand U22162(n21116,n20846,n19750);
  nand U22163(n21112,n21119,n21120,n21121,n21096);
  nand U22164(n21121,n20190,n20869);
  nand U22165(n21120,n20191,n20838);
  nand U22166(n21119,n20839,n19750);
  nand U22167(n21114,n21122,n21123,n21124,n21096);
  nand U22168(n21123,n20873,n20202);
  nand U22169(n21113,n21125,n21126,n21127);
  nand U22170(n21127,n21128,n21129);
  nand U22171(n21129,n21122,n21130);
  nand U22172(n21130,n20202,n20869);
  and U22173(n21122,n21131,n21132);
  nand U22174(n21132,n20203,n20838);
  nand U22175(n21131,n20839,n19753);
  not U22176(n21128,n21124);
  nand U22177(n21124,n21133,n21134,n21135);
  nand U22178(n21135,n20843,n20203);
  nand U22179(n21134,n20844,n20202);
  nand U22180(n21133,n20846,n19753);
  nand U22181(n21126,n21136,n21137);
  nand U22182(n21125,n21138,n21139,n21140);
  or U22183(n21140,n21137,n21136);
  and U22184(n21136,n21141,n21142,n21143);
  nand U22185(n21143,n20843,n20215);
  nand U22186(n21142,n20844,n20214);
  nand U22187(n21141,n20846,n19756);
  nand U22188(n21137,n21144,n21145,n21146,n21096);
  nand U22189(n21146,n20214,n20869);
  nand U22190(n21145,n20215,n20838);
  nand U22191(n21144,n20839,n19756);
  nand U22192(n21139,n21147,n21148,n21149,n21096);
  nand U22193(n21148,n20873,n20226);
  nand U22194(n21138,n21150,n21151,n21152);
  nand U22195(n21152,n21153,n21154);
  nand U22196(n21154,n21147,n21155);
  nand U22197(n21155,n20226,n20869);
  and U22198(n21147,n21156,n21157);
  nand U22199(n21157,n20227,n20838);
  nand U22200(n21156,n20839,n19759);
  not U22201(n21153,n21149);
  nand U22202(n21149,n21158,n21159,n21160);
  nand U22203(n21160,n20843,n20227);
  nand U22204(n21159,n20844,n20226);
  nand U22205(n21158,n20846,n19759);
  nand U22206(n21151,n21161,n21162);
  nand U22207(n21150,n21163,n21164,n21165);
  or U22208(n21165,n21162,n21161);
  and U22209(n21161,n21166,n21167,n21168);
  nand U22210(n21168,n20843,n20239);
  nand U22211(n21167,n20844,n20238);
  nand U22212(n21166,n20846,n19762);
  nand U22213(n21162,n21169,n21170,n21171,n21096);
  nand U22214(n21171,n20238,n20869);
  nand U22215(n21170,n20239,n20838);
  nand U22216(n21169,n20839,n19762);
  nand U22217(n21164,n21172,n21173,n21174,n21096);
  nand U22218(n21173,n20873,n20250);
  nand U22219(n21163,n21175,n21176,n21177);
  nand U22220(n21177,n21178,n21179);
  nand U22221(n21179,n21172,n21180);
  nand U22222(n21180,n20250,n20869);
  and U22223(n21172,n21181,n21182);
  nand U22224(n21182,n20251,n20838);
  nand U22225(n21181,n20839,n19765);
  not U22226(n21178,n21174);
  nand U22227(n21174,n21183,n21184,n21185);
  nand U22228(n21185,n20843,n20251);
  nand U22229(n21184,n20844,n20250);
  nand U22230(n21183,n20846,n19765);
  nand U22231(n21176,n21186,n21187);
  nand U22232(n21175,n21188,n21189,n21190);
  or U22233(n21190,n21187,n21186);
  and U22234(n21186,n21191,n21192,n21193);
  nand U22235(n21193,n19795,n20843);
  nand U22236(n21192,n20844,n19786);
  nand U22237(n21191,n20846,n19768);
  nand U22238(n21187,n21194,n21195,n21196,n21096);
  nand U22239(n21196,n19786,n20869);
  nand U22240(n21195,n19795,n20838);
  nand U22241(n21194,n20839,n19768);
  nand U22242(n21189,n21197,n21198,n21199,n21200);
  nor U22243(n21200,n21201,n21202);
  nor U22244(n21201,n21203,n20688);
  nand U22245(n21199,n21204,n21205);
  or U22246(n21188,n21205,n21204);
  and U22247(n21204,n21206,n21207,n21208);
  nand U22248(n21208,n20843,n20268);
  nand U22249(n21207,n20844,n20273);
  nand U22250(n21206,n20846,n19771);
  nand U22251(n21205,n21209,n21210,n21211,n21096);
  nand U22252(n21211,n20873,n20273);
  nand U22253(n21210,n20268,n20838);
  nand U22254(n21209,n20839,n19771);
  nand U22255(n20851,n21212,n21213,n21214);
  nand U22256(n21214,n20843,n19938);
  nand U22257(n21213,n20844,n19937);
  nand U22258(n21212,n20846,n19687);
  nand U22259(n20854,n20873,n19937);
  not U22260(n20873,n21215);
  nand U22261(n20853,n19938,n20838);
  nand U22262(n20852,n20839,n19687);
  nand U22263(n20847,n21216,n21217);
  or U22264(n20833,n21217,n21216);
  and U22265(n21216,n21218,n21219,n21220);
  nand U22266(n21220,n20839,n19684);
  nand U22267(n21219,n19923,n20869);
  nand U22268(n20869,n21096,n21215);
  nand U22269(n21215,n21221,n21222);
  and U22270(n21096,n20629,n21223);
  nand U22271(n21218,n19920,n20838);
  nand U22272(n21217,n21224,n21225,n21226);
  nand U22273(n21226,n20843,n19920);
  nand U22274(n21225,n20844,n19923);
  nand U22275(n21224,n20846,n19684);
  or U22276(n20828,n20827,n20826);
  and U22277(n20826,n21227,n21228);
  nand U22278(n21228,n19905,n20838);
  nand U22279(n21227,n20839,n19678);
  nand U22280(n21231,n21232,n20269,n21221);
  nand U22281(n20827,n21233,n21234,n21235);
  nand U22282(n21235,n20843,n19905);
  nand U22283(n21232,n20625,n21236);
  nand U22284(n21236,n21237,n21198);
  not U22285(n20269,n21238);
  nand U22286(n21234,n21239,n20844);
  xor U22287(n21239,n21241,n21242);
  xnor U22288(n21242,n20845,n21243);
  and U22289(n20845,n21244,n21245);
  nand U22290(n21244,n21246,n21247);
  nand U22291(n21233,n20846,n19678);
  nor U22292(n21229,n19787,n21203,n21249);
  and U22293(n21249,n20612,n21250);
  nand U22294(n21250,n20611,n21202);
  nor U22295(n21203,n20286,n20644);
  or U22296(n21248,n21230,n21221);
  not U22297(n21221,n21240);
  nand U22298(n21240,n20692,n19681);
  not U22299(n20692,n19678);
  nand U22300(n21230,n21251,n21252);
  nand U22301(n21252,n21237,n21253);
  nand U22302(n21253,n20644,n20277);
  nand U22303(n21223,n20272,n21251);
  nor U22304(n20823,n21254,n19787,n21255);
  nor U22305(n21255,n21237,n21251,n21256);
  not U22306(n19787,n20621);
  nor U22307(n21254,n20611,n20620);
  nand U22308(n20626,G36185,n21257);
  nand U22309(n21257,n21258,n21259,n21260);
  nand U22310(n21259,n20277,n20602);
  nand U22311(n21258,n20611,n21261);
  nand U22312(n21261,n21202,G36215,n20596,n21262);
  nor U22313(n21262,n21263,n21264);
  nand U22314(G1519,n21265,n21266,n21267,n21268);
  nor U22315(n21268,n21269,n21270);
  nor U22316(n21270,G36215,n20506);
  and U22317(n21269,n21271,G36152);
  nand U22318(n21267,n21272,n20273);
  nand U22319(n21266,n21273,n21274,n21275);
  nand U22320(n21273,n21276,n21277);
  nand U22321(n21265,G35973,n21278);
  nand U22322(G1518,n21279,n21280,n21281,n21282);
  nor U22323(n21282,n21283,n21284);
  nor U22324(n21284,G36215,n19780);
  not U22325(n19780,G36205);
  nor U22326(n21283,n21285,n21286);
  nand U22327(n21281,n21287,n21278);
  nand U22328(n21280,n21288,n21275);
  xnor U22329(n21288,n21289,n21290);
  xor U22330(n21290,n21287,n21291);
  nand U22331(n21279,n21272,n19786);
  xor U22332(n19786,n21292,n21293);
  and U22333(n21293,n21294,n21295);
  nand U22334(G1517,n21296,n21297,n21298,n21299);
  nor U22335(n21299,n21300,n21301,n21302);
  nor U22336(n21302,n21303,n21304);
  xnor U22337(n21303,n21305,n21306);
  xor U22338(n21305,n21307,n21308);
  nor U22339(n21300,n21309,n21310);
  nand U22340(n21298,G36190,G1406);
  nand U22341(n21297,n21272,n20250);
  nand U22342(n21296,G36150,n21271);
  nand U22343(G1516,n21311,n21312,n21313,n21314);
  nor U22344(n21314,n21315,n20358);
  nor U22345(n20358,G36215,n21316);
  nor U22346(n21315,n21285,n21317);
  nand U22347(n21313,n21272,n20238);
  nand U22348(n21312,n21318,n21275);
  xor U22349(n21318,n21319,n21320);
  xor U22350(n21320,n21321,n21322);
  nand U22351(n21311,n21322,n21278);
  nand U22352(G1515,n21323,n21324,n20481,n21325);
  nor U22353(n21325,n21326,n21301,n21327);
  nor U22354(n21327,n21328,n21304);
  xnor U22355(n21328,n21329,n21330);
  and U22356(n21330,n21331,n21332);
  and U22357(n21301,n21333,n21334,G1625);
  nand U22358(n21334,n20598,n21277);
  or U22359(n21333,n20273,n20598);
  nor U22360(n21326,n21309,n21336);
  not U22361(n21309,n21278);
  nand U22362(n20481,G36197,G1406);
  nand U22363(n21324,n21272,n20226);
  nand U22364(n21323,G36148,n21271);
  nand U22365(G1514,n21337,n21338,n21339,n21340);
  nor U22366(n21340,n21341,n21342);
  and U22367(n21342,G1406,G36200);
  and U22368(n21341,n21271,G36147);
  nand U22369(n21339,n21272,n20214);
  nand U22370(n21338,n21343,n21275);
  xnor U22371(n21343,n21344,n21345);
  nand U22372(n21344,n21346,n21347);
  nand U22373(n21337,n21348,n21278);
  nand U22374(G1513,n21349,n21350,n21351,n21352);
  nor U22375(n21352,n21353,n21354);
  nor U22376(n21354,G36215,n21355);
  and U22377(n21353,n21271,G36146);
  nand U22378(n21351,n21272,n20202);
  nand U22379(n21350,n21356,n21275);
  xnor U22380(n21356,n21357,n21358);
  nand U22381(n21357,n21359,n21360);
  nand U22382(n21349,n21361,n21278);
  nand U22383(G1512,n21362,n21363,n21364,n21365);
  nor U22384(n21365,n21366,n21367);
  nor U22385(n21367,G36215,n21368);
  and U22386(n21366,n21271,G36145);
  nand U22387(n21364,n21272,n20190);
  nand U22388(n21363,n21275,n21369);
  xnor U22389(n21369,n21370,n21371);
  xor U22390(n21370,n21372,n21373);
  nand U22391(n21362,n21374,n21278);
  nand U22392(G1511,n21375,n21376,n21377,n21378);
  nor U22393(n21378,n21379,n21380);
  and U22394(n21380,G1406,G36206);
  nor U22395(n21379,n21285,n21381);
  nand U22396(n21377,n21272,n20178);
  nand U22397(n21376,n21275,n21382);
  xnor U22398(n21382,n21383,n21384);
  xor U22399(n21384,n21385,n21386);
  nand U22400(n21375,n21387,n21278);
  nand U22401(G1510,n21388,n21389,n21390,n21391);
  nor U22402(n21391,n21392,n21393);
  nor U22403(n21393,G36215,n21394);
  nor U22404(n21392,n21285,n21395);
  nand U22405(n21390,n21272,n20166);
  nand U22406(n21389,n21396,n21275);
  xor U22407(n21396,n21397,n21398);
  xor U22408(n21398,n21399,n21400);
  nand U22409(n21388,n21400,n21278);
  nand U22410(G1509,n21401,n21402,n21403,n21404);
  nor U22411(n21404,n21405,n21406);
  nor U22412(n21406,G36215,n21407);
  nor U22413(n21405,n21285,n21408);
  nand U22414(n21403,n21272,n20154);
  nand U22415(n21402,n21275,n21409);
  nand U22416(n21409,n21410,n21411);
  nand U22417(n21411,n21412,n21413);
  nand U22418(n21413,n21414,n21415);
  not U22419(n21414,n21416);
  nand U22420(n21410,n21417,n21418);
  nand U22421(n21401,n21419,n21278);
  nand U22422(G1508,n21420,n21421,n21422,n21423);
  nor U22423(n21423,n21424,n21425);
  and U22424(n21425,G1406,G36191);
  nor U22425(n21424,n21285,n21426);
  nand U22426(n21422,n21272,n20142);
  nand U22427(n21421,n21275,n21427);
  xnor U22428(n21427,n21428,n21429);
  xor U22429(n21428,n21430,n21417);
  nand U22430(n21420,n21431,n21278);
  nand U22431(G1507,n21432,n21433,n21434,n21435);
  nor U22432(n21435,n21436,n21437);
  nor U22433(n21437,G36215,n21438);
  and U22434(n21436,n21271,G36140);
  nand U22435(n21434,n21272,n20130);
  nand U22436(n21433,n21439,n21275);
  xor U22437(n21439,n21440,n21441);
  xor U22438(n21441,n21442,n21443);
  nand U22439(n21432,n21443,n21278);
  nand U22440(G1506,n21444,n21445,n21446,n21447);
  nor U22441(n21447,n21448,n21449);
  and U22442(n21449,G1406,G36193);
  nor U22443(n21448,n21285,n21450);
  nand U22444(n21446,n21272,n20118);
  nand U22445(n21445,n21275,n21451);
  xnor U22446(n21451,n21452,n21453);
  xor U22447(n21453,n21454,n21455);
  nand U22448(n21444,n21456,n21278);
  nand U22449(G1505,n21457,n21458,n21459,n21460);
  nor U22450(n21460,n21461,n21462);
  nor U22451(n21462,G36215,n21463);
  nor U22452(n21461,n21285,n21464);
  nand U22453(n21459,n21272,n20106);
  nand U22454(n21458,n21275,n21465);
  nand U22455(n21465,n21466,n21467);
  nand U22456(n21467,n21468,n21469);
  nand U22457(n21466,n21470,n21471);
  nand U22458(n21471,n21472,n21473);
  not U22459(n21472,n21474);
  nand U22460(n21457,n21475,n21278);
  nand U22461(G1504,n21476,n21477,n21478,n21479);
  nor U22462(n21479,n21480,n21481);
  and U22463(n21481,G1406,G36186);
  nor U22464(n21480,n21285,n21482);
  nand U22465(n21478,n21272,n20094);
  nand U22466(n21477,n21483,n21275);
  xor U22467(n21483,n21484,n21468);
  not U22468(n21468,n21485);
  nand U22469(n21484,n21486,n21487);
  nand U22470(n21476,n21488,n21278);
  nand U22471(G1503,n21489,n21490,n21491,n21492);
  nor U22472(n21492,n21493,n21494);
  nor U22473(n21494,G36215,n21495);
  nor U22474(n21493,n21285,n21496);
  nand U22475(n21491,n21272,n20082);
  nand U22476(n21490,n21497,n21275);
  xnor U22477(n21497,n21498,n21499);
  xnor U22478(n21499,n21500,n21501);
  nand U22479(n21489,n21501,n21278);
  nand U22480(G1502,n21502,n21503,n21504,n21505);
  nor U22481(n21505,n21506,n21507);
  and U22482(n21507,G1406,G36199);
  nor U22483(n21506,n21285,n21508);
  nand U22484(n21504,n21272,n20070);
  nand U22485(n21503,n21509,n21275);
  xnor U22486(n21509,n21510,n21511);
  xnor U22487(n21510,n21512,n21513);
  nand U22488(n21502,n21513,n21278);
  nand U22489(G1501,n21514,n21515,n21516,n21517);
  nor U22490(n21517,n21518,n21519);
  nor U22491(n21519,G36215,n21520);
  nor U22492(n21518,n21285,n21521);
  nand U22493(n21516,n21272,n20058);
  nand U22494(n21515,n21522,n21275);
  xnor U22495(n21522,n21523,n21524);
  xor U22496(n21524,n21525,n21526);
  nand U22497(n21514,n21527,n21278);
  nand U22498(G1500,n21528,n21529,n21530,n21531);
  nor U22499(n21531,n21532,n21533);
  nor U22500(n21533,G36215,n21534);
  nor U22501(n21532,n21535,n21285);
  nand U22502(n21530,n21272,n20046);
  and U22503(n21272,n20282,n21536,n21285,n21537);
  not U22504(n21537,n21538);
  nand U22505(n21529,n21275,n21539);
  xor U22506(n21539,n21540,n21541);
  nor U22507(n21541,n21542,n21543);
  nor U22508(n21543,n21544,n21545);
  xor U22509(n21545,n20635,G36088);
  nor U22510(n21542,n21264,n21546);
  xor U22511(n21546,n20635,G36120);
  nand U22512(n21540,n21547,n21548);
  nand U22513(n21548,n21526,n21549);
  nand U22514(n21549,n21523,n21525);
  or U22515(n21547,n21525,n21523);
  and U22516(n21523,n21550,n21551);
  or U22517(n21551,n21544,G36087);
  or U22518(n21550,n21264,G36119);
  nand U22519(n21525,n21552,n21553);
  nand U22520(n21553,n21513,n21554);
  nand U22521(n21554,n21512,n21511);
  or U22522(n21552,n21511,n21512);
  and U22523(n21512,n21555,n21556);
  nand U22524(n21556,n21501,n21557);
  or U22525(n21557,n21500,n21498);
  nand U22526(n21555,n21498,n21500);
  nand U22527(n21500,n21558,n21487);
  nand U22528(n21487,n21559,n21560,n21488);
  or U22529(n21560,n21544,G36084);
  or U22530(n21559,n21264,G36116);
  nand U22531(n21558,n21486,n21485);
  nand U22532(n21485,n21473,n21474);
  nand U22533(n21474,n21470,n21469);
  nand U22534(n21469,n21561,n21562,n21563);
  nand U22535(n21562,n21544,G36115);
  nand U22536(n21561,n21264,G36083);
  and U22537(n21470,n21564,n21565);
  nand U22538(n21565,n21455,n21566);
  or U22539(n21566,n21452,n21454);
  nand U22540(n21564,n21452,n21454);
  nand U22541(n21454,n21567,n21568);
  nand U22542(n21568,n21569,n21570);
  or U22543(n21569,n21440,n21442);
  nand U22544(n21567,n21440,n21442);
  nand U22545(n21442,n21571,n21572);
  nand U22546(n21572,n21573,n21430);
  or U22547(n21573,n21429,n21417);
  nand U22548(n21571,n21417,n21429);
  nand U22549(n21429,n21574,n21575);
  or U22550(n21575,n21544,G36080);
  or U22551(n21574,n21264,G36112);
  and U22552(n21417,n21415,n21416);
  nand U22553(n21416,n21412,n21418);
  nand U22554(n21418,n21576,n21577);
  and U22555(n21412,n21578,n21579);
  nand U22556(n21579,n21580,n21581);
  or U22557(n21580,n21397,n21399);
  nand U22558(n21578,n21397,n21399);
  nand U22559(n21399,n21582,n21583);
  nand U22560(n21583,n21386,n21584);
  or U22561(n21584,n21383,n21385);
  nand U22562(n21582,n21383,n21385);
  nand U22563(n21385,n21585,n21586);
  nand U22564(n21586,n21587,n21372);
  or U22565(n21587,n21371,n21373);
  nand U22566(n21585,n21373,n21371);
  nand U22567(n21371,n21588,n21589);
  or U22568(n21589,n21544,G36076);
  or U22569(n21588,n21264,G36108);
  and U22570(n21373,n21590,n21360);
  nand U22571(n21360,n21591,n21592,n21361);
  or U22572(n21592,n21544,G36075);
  or U22573(n21591,n21264,G36107);
  nand U22574(n21590,n21358,n21359);
  nand U22575(n21359,n21593,n21594,n21595);
  nand U22576(n21594,n21544,G36107);
  nand U22577(n21593,n21264,G36075);
  nand U22578(n21358,n21347,n21596);
  nand U22579(n21596,n21346,n21345);
  nand U22580(n21345,n21331,n21597);
  nand U22581(n21597,n21329,n21332);
  nand U22582(n21332,n21598,n21599,n21336);
  nand U22583(n21599,n21544,G36105);
  nand U22584(n21598,n21264,G36073);
  and U22585(n21329,n21600,n21601);
  nand U22586(n21601,n21602,n21603);
  or U22587(n21602,n21319,n21321);
  nand U22588(n21600,n21319,n21321);
  nand U22589(n21321,n21604,n21605);
  nand U22590(n21605,n21310,n21606);
  or U22591(n21606,n21306,n21307);
  nand U22592(n21604,n21306,n21307);
  nand U22593(n21307,n21607,n21608);
  nand U22594(n21608,n21609,n21610);
  or U22595(n21609,n21289,n21274);
  nand U22596(n21607,n21289,n21274);
  not U22597(n21274,n21291);
  nor U22598(n21291,n21276,n21277);
  nand U22599(n21289,n21611,n21612);
  or U22600(n21612,n21544,G36070);
  nand U22601(n21611,n21544,n19790);
  not U22602(n19790,G36102);
  nand U22603(n21306,n21613,n21614);
  or U22604(n21614,n21544,G36071);
  or U22605(n21613,n21264,G36103);
  nand U22606(n21319,n21615,n21616);
  or U22607(n21616,n21544,G36072);
  or U22608(n21615,n21264,G36104);
  nand U22609(n21331,n21617,n21618,n21619);
  or U22610(n21618,n21544,G36073);
  or U22611(n21617,n21264,G36105);
  nand U22612(n21346,n21620,n21621,n21622);
  not U22613(n21622,n21348);
  nand U22614(n21621,n21544,G36106);
  nand U22615(n21620,n21264,G36074);
  nand U22616(n21347,n21623,n21624,n21348);
  or U22617(n21624,n21544,G36074);
  or U22618(n21623,n21264,G36106);
  nand U22619(n21383,n21625,n21626);
  or U22620(n21626,n21544,G36077);
  or U22621(n21625,n21264,G36109);
  nand U22622(n21397,n21627,n21628);
  or U22623(n21628,n21544,G36078);
  or U22624(n21627,n21264,G36110);
  or U22625(n21415,n21576,n21577);
  nand U22626(n21576,n21629,n21630);
  or U22627(n21630,n21544,G36079);
  or U22628(n21629,n21264,G36111);
  nand U22629(n21440,n21631,n21632);
  or U22630(n21632,n21544,G36081);
  or U22631(n21631,n21264,G36113);
  nand U22632(n21452,n21633,n21634);
  or U22633(n21634,n21544,G36082);
  or U22634(n21633,n21264,G36114);
  nand U22635(n21473,n21635,n21636,n21475);
  or U22636(n21636,n21544,G36083);
  or U22637(n21635,n21264,G36115);
  nand U22638(n21486,n21637,n21638,n21639);
  nand U22639(n21638,n21544,G36116);
  nand U22640(n21637,n21264,G36084);
  and U22641(n21498,n21640,n21641);
  or U22642(n21641,n21544,G36085);
  or U22643(n21640,n21264,G36117);
  nand U22644(n21511,n21642,n21643);
  or U22645(n21643,n21544,G36086);
  or U22646(n21642,n21264,G36118);
  not U22647(n21275,n21304);
  nand U22648(n21304,n21644,n21536);
  nand U22649(n21536,n21544,n20598);
  nand U22650(n21644,n21645,n21646);
  nand U22651(n21646,n21647,n21285,n20282);
  nand U22652(n21647,n20621,n21237,n21263,n20620);
  not U22653(n21645,n21648);
  nand U22654(n21528,n20644,n21278);
  nand U22655(n21278,n21649,n21650);
  nand U22656(n21650,n20282,n21651,n20598,n21285);
  not U22657(n21285,n21271);
  nand U22658(n21651,n21538,n20621,n21652);
  nor U22659(n21652,n21653,n20688,n20612);
  not U22660(n20688,n20620);
  nand U22661(n21649,n21648,n20598);
  nor U22662(n21648,n20602,n21271);
  nor U22663(n21271,n21335,G1341);
  not U22664(n21335,n21260);
  nand U22665(n20602,n20629,G36215);
  nand U22666(G1499,n21654,n21655,n21656);
  nand U22667(n21656,n19794,n19905);
  nand U22668(n21655,G36132,n19783);
  nand U22669(n21654,n19789,n21657);
  nand U22670(n21657,n19900,n21658);
  nand U22671(n21658,n21659,n19902);
  xor U22672(n19902,n21660,n21661);
  xor U22673(n21660,n21662,n21663);
  nand U22674(n21662,n21664,n21665);
  nand U22675(n21665,n21666,n19905);
  nand U22676(n19905,n21667,n21668);
  nand U22677(n21668,n21669,n17853);
  nand U22678(n21667,n21670,G36429);
  nand U22679(G1498,n21671,n21672,n21673);
  nand U22680(n21673,n19794,n19911);
  nand U22681(n21672,G36131,n19783);
  nand U22682(n21671,n19789,n21674);
  nand U22683(n21674,n19900,n21675);
  nand U22684(n21675,n19912,n19913,n21659);
  nand U22685(n19913,n21661,n21676);
  nand U22686(n21676,n21664,n21677);
  nor U22687(n21661,n21678,n21679);
  nand U22688(n19912,n21679,n21678);
  nand U22689(n21678,n21680,n21681);
  nand U22690(n21680,n21682,n21683);
  and U22691(n21679,n21663,n21684);
  nand U22692(n21684,n21664,n21685);
  nand U22693(n21685,n21666,n19911);
  nand U22694(n19911,n21686,n21687);
  nand U22695(n21687,n21669,n17869);
  nand U22696(n21686,n21670,G36428);
  nand U22697(n19900,n19678,n21688);
  nand U22698(n21688,n21689,n21690);
  nand U22699(n21690,n21691,n21692);
  or U22700(n21689,n19936,G36185);
  nand U22701(n19678,n21693,n21694,n21695);
  nand U22702(n21695,G36068,n21696);
  nand U22703(n21694,G36132,n21697);
  nand U22704(n21693,G36100,n21698);
  nand U22705(G1497,n21699,n21700,n21701,n21702);
  nor U22706(n21702,n21703,n21704,n21705);
  nor U22707(n21705,n19783,n19919);
  nand U22708(n19919,n21706,n21707,n21692);
  nand U22709(n21707,n21708,n20598);
  nand U22710(n21708,n19681,n21709);
  nand U22711(n21709,G36185,n21710);
  nand U22712(n19681,n21711,n21712,n21713);
  nand U22713(n21713,G36067,n21696);
  nand U22714(n21712,G36131,n21697);
  nand U22715(n21711,G36099,n21698);
  nand U22716(n21706,n19949,n20596);
  and U22717(n21704,n19783,G36130);
  nor U22718(n21703,n20820,n21714);
  not U22719(n20820,n19920);
  nand U22720(n21701,n21715,n19923);
  xor U22721(n19923,n21246,n21716);
  and U22722(n21716,n21247,n21245);
  nand U22723(n21245,n21717,n21718);
  nand U22724(n21718,n21243,n21719);
  not U22725(n21717,n21241);
  nand U22726(n21247,n21241,n21719,n21243);
  and U22727(n21243,n21720,n21721,n21722,n21723);
  nand U22728(n21723,n21724,n19938);
  nand U22729(n21722,n21725,n19920);
  nand U22730(n21721,n21726,n19684);
  nand U22731(n21719,n20629,n19684);
  xor U22732(n21241,n21727,n21728);
  nand U22733(n21727,n21729,n21730,n21731,n21732);
  nand U22734(n21731,n19920,n21726);
  nand U22735(n21730,n21725,n19684);
  nand U22736(n21729,n21724,n19687);
  nand U22737(n21246,n21733,n21734);
  nand U22738(n21734,n21735,n21736);
  nand U22739(n21700,n21737,n21738);
  nand U22740(n21699,n19792,n19921);
  xnor U22741(n19921,n21682,n21739);
  and U22742(n21739,n21683,n21681);
  nand U22743(n21681,n21740,n21741,n21663);
  nand U22744(n21741,n21664,n21742);
  nand U22745(n21742,n21666,n19920);
  not U22746(n21666,n21743);
  nand U22747(n21683,n21664,n21744);
  nand U22748(n21744,n21663,n21740);
  nand U22749(n21740,n21256,n19684);
  not U22750(n21663,n21677);
  nand U22751(n21677,n21745,n21746);
  or U22752(n21746,n21747,n19949);
  nand U22753(n21745,n21748,n19684);
  and U22754(n21664,n21749,n21750);
  nand U22755(n21750,n21748,n19920);
  nand U22756(n19920,n21751,n21752);
  nand U22757(n21752,n21669,n17943);
  nand U22758(n21751,n21670,G36427);
  not U22759(n21748,n21753);
  nand U22760(n21749,n19938,n21754);
  nand U22761(n21754,n21755,n21747);
  nand U22762(n21682,n21756,n21757);
  nand U22763(n21757,n21758,n21759);
  nand U22764(G1496,n21760,n21761,n21762,n21763);
  nor U22765(n21763,n21764,n21765,n21766,n21767);
  nor U22766(n21767,n20388,n21714);
  and U22767(n21766,n19937,n21715);
  xor U22768(n19937,n21736,n21768);
  and U22769(n21768,n21735,n21733);
  nand U22770(n21733,n21769,n21770);
  or U22771(n21735,n21769,n21770);
  nand U22772(n21770,n21771,n21772,n21720);
  nand U22773(n21772,n19938,n21773);
  nand U22774(n21771,n19687,n21774);
  xor U22775(n21769,n21775,n21776);
  nand U22776(n21775,n21777,n21732,n21778);
  nand U22777(n21778,n21773,n19687);
  nand U22778(n21777,n19938,n21779);
  nand U22779(n21736,n21780,n21781);
  nand U22780(n21781,n21782,n21783);
  nor U22781(n21765,n20703,n21784);
  xor U22782(n20703,n21759,n21785);
  and U22783(n21785,n21786,n21756,n21758);
  nand U22784(n21758,n19687,n21787,n20388);
  not U22785(n20388,n19938);
  nand U22786(n21756,n19938,n21788,n21789);
  nand U22787(n21789,n19687,n21787);
  nand U22788(n19938,n21790,n21791);
  nand U22789(n21791,n21669,n17982);
  nand U22790(n21790,n21670,G36426);
  nand U22791(n21786,n19687,n20819);
  nand U22792(n21759,n21792,n21793);
  nand U22793(n21793,n21794,n21795);
  nor U22794(n21764,n19935,n21796);
  not U22795(n19935,n19684);
  nand U22796(n19684,n21797,n21798,n21799,n21800);
  nand U22797(n21800,n21738,n21801);
  nand U22798(n21799,G36130,n21697);
  nand U22799(n21798,G36098,n21698);
  nand U22800(n21797,G36066,n21696);
  nand U22801(n21762,G36129,n19783);
  nand U22802(n21761,n21737,n20387);
  nand U22803(G1495,n21802,n21803,n21804,n21805);
  nor U22804(n21805,n21806,n21807,n21808,n21809);
  nor U22805(n21809,n20322,n21714);
  and U22806(n21808,n19950,n21715);
  xor U22807(n19950,n21783,n21810);
  and U22808(n21810,n21782,n21780);
  nand U22809(n21780,n21811,n21812);
  or U22810(n21782,n21811,n21812);
  nand U22811(n21812,n21813,n21814,n21720);
  nand U22812(n21814,n19951,n21773);
  nand U22813(n21813,n19690,n21774);
  xor U22814(n21811,n21815,n21776);
  nand U22815(n21815,n21816,n21732,n21817);
  nand U22816(n21817,n21773,n19690);
  nand U22817(n21816,n19951,n21779);
  nand U22818(n21783,n21818,n21819);
  nand U22819(n21819,n21820,n21821);
  nor U22820(n21807,n20707,n21784);
  xor U22821(n20707,n21795,n21822);
  and U22822(n21822,n21823,n21792,n21794);
  nand U22823(n21794,n19690,n21787,n20322);
  not U22824(n20322,n19951);
  nand U22825(n21792,n19951,n21788,n21824);
  nand U22826(n21824,n19690,n21787);
  nand U22827(n19951,n21825,n21826);
  nand U22828(n21826,n21669,n18022);
  nand U22829(n21825,n21670,G36425);
  nand U22830(n21823,n19690,n20819);
  nand U22831(n21795,n21827,n21828);
  nand U22832(n21828,n21829,n21830);
  nor U22833(n21806,n19949,n21796);
  not U22834(n19949,n19687);
  nand U22835(n19687,n21831,n21832,n21833,n21834);
  nand U22836(n21834,n20387,n21801);
  nor U22837(n20387,n21738,n21835);
  and U22838(n21835,n21836,n21837);
  nor U22839(n21738,n21837,n21836);
  not U22840(n21837,G36207);
  nand U22841(n21833,G36129,n21697);
  nand U22842(n21832,G36097,n21698);
  nand U22843(n21831,G36065,n21696);
  nand U22844(n21804,G36128,n19783);
  nand U22845(n21803,n21737,n21838);
  nand U22846(G1494,n21839,n21840,n21841,n21842);
  nor U22847(n21842,n21843,n21844,n21845,n21846);
  nor U22848(n21846,n20586,n21714);
  and U22849(n21845,n19962,n21715);
  xor U22850(n19962,n21821,n21847);
  and U22851(n21847,n21820,n21818);
  nand U22852(n21818,n21848,n21849);
  or U22853(n21820,n21848,n21849);
  nand U22854(n21849,n21850,n21851,n21720);
  nand U22855(n21851,n19963,n21773);
  nand U22856(n21850,n19693,n21774);
  xor U22857(n21848,n21852,n21776);
  nand U22858(n21852,n21853,n21732,n21854);
  nand U22859(n21854,n21773,n19693);
  nand U22860(n21853,n19963,n21779);
  nand U22861(n21821,n21855,n21856);
  nand U22862(n21856,n21857,n21858);
  nor U22863(n21844,n20711,n21784);
  xor U22864(n20711,n21830,n21859);
  and U22865(n21859,n21860,n21827,n21829);
  nand U22866(n21829,n19693,n21787,n20586);
  not U22867(n20586,n19963);
  nand U22868(n21827,n19963,n21788,n21861);
  nand U22869(n21861,n19693,n21787);
  nand U22870(n19963,n21862,n21863);
  nand U22871(n21863,n21669,n18063);
  nand U22872(n21862,n21670,G36424);
  nand U22873(n21860,n19693,n20819);
  nand U22874(n21830,n21864,n21865);
  nand U22875(n21865,n21866,n21867);
  nor U22876(n21843,n19933,n21796);
  not U22877(n19933,n19690);
  nand U22878(n19690,n21868,n21869,n21870,n21871);
  nand U22879(n21871,n21838,n21801);
  not U22880(n21838,n20321);
  nand U22881(n20321,n21872,n21836);
  or U22882(n21836,n21873,n21874);
  nand U22883(n21872,n21873,n21874);
  nand U22884(n21874,G36187,n21875,G36202);
  not U22885(n21873,G36213);
  nand U22886(n21870,G36128,n21697);
  nand U22887(n21869,G36096,n21698);
  nand U22888(n21868,G36064,n21696);
  nand U22889(n21841,G36127,n19783);
  nand U22890(n21840,n21737,n21876);
  nand U22891(G1493,n21877,n21878,n21879,n21880);
  nor U22892(n21880,n21881,n21882,n21883,n21884);
  nor U22893(n21884,n20438,n21714);
  and U22894(n21883,n19974,n21715);
  xor U22895(n19974,n21858,n21885);
  and U22896(n21885,n21857,n21855);
  nand U22897(n21855,n21886,n21887);
  or U22898(n21857,n21886,n21887);
  nand U22899(n21887,n21888,n21889,n21720);
  nand U22900(n21889,n19975,n21773);
  nand U22901(n21888,n19696,n21774);
  xor U22902(n21886,n21890,n21776);
  nand U22903(n21890,n21891,n21732,n21892);
  nand U22904(n21892,n21773,n19696);
  nand U22905(n21891,n19975,n21779);
  nand U22906(n21858,n21893,n21894);
  nand U22907(n21894,n21895,n21896);
  nor U22908(n21882,n20715,n21784);
  xor U22909(n20715,n21867,n21897);
  and U22910(n21897,n21898,n21864,n21866);
  nand U22911(n21866,n19696,n21787,n20438);
  not U22912(n20438,n19975);
  nand U22913(n21864,n19975,n21788,n21899);
  nand U22914(n21899,n19696,n21787);
  nand U22915(n19975,n21900,n21901);
  nand U22916(n21901,n21669,n18105);
  nand U22917(n21900,n21670,G36423);
  nand U22918(n21898,n19696,n20819);
  nand U22919(n21867,n21902,n21903);
  nand U22920(n21903,n21904,n21905);
  nor U22921(n21881,n19948,n21796);
  not U22922(n19948,n19693);
  nand U22923(n19693,n21906,n21907,n21908,n21909);
  nand U22924(n21909,n21876,n21801);
  not U22925(n21876,n20585);
  xnor U22926(n20585,G36187,n21910);
  and U22927(n21910,n21875,G36202);
  nand U22928(n21908,G36127,n21697);
  nand U22929(n21907,G36095,n21698);
  nand U22930(n21906,G36063,n21696);
  nand U22931(n21879,G36126,n19783);
  nand U22932(n21878,n21737,n20437);
  nand U22933(G1492,n21911,n21912,n21913,n21914);
  nor U22934(n21914,n21915,n21916,n21917,n21918);
  nor U22935(n21918,n20478,n21714);
  and U22936(n21917,n19986,n21715);
  xor U22937(n19986,n21896,n21919);
  and U22938(n21919,n21895,n21893);
  nand U22939(n21893,n21920,n21921);
  or U22940(n21895,n21920,n21921);
  nand U22941(n21921,n21922,n21923,n21720);
  nand U22942(n21923,n19987,n21773);
  nand U22943(n21922,n19699,n21774);
  xor U22944(n21920,n21924,n21776);
  nand U22945(n21924,n21925,n21732,n21926);
  nand U22946(n21926,n21773,n19699);
  nand U22947(n21925,n19987,n21779);
  nand U22948(n21896,n21927,n21928);
  nand U22949(n21928,n21929,n21930);
  nor U22950(n21916,n20719,n21784);
  xor U22951(n20719,n21905,n21931);
  and U22952(n21931,n21932,n21902,n21904);
  nand U22953(n21904,n19699,n21787,n20478);
  not U22954(n20478,n19987);
  nand U22955(n21902,n19987,n21788,n21933);
  nand U22956(n21933,n19699,n21787);
  nand U22957(n19987,n21934,n21935);
  nand U22958(n21935,n21669,n18143);
  nand U22959(n21934,n21670,G36422);
  nand U22960(n21932,n19699,n20819);
  nand U22961(n21905,n21936,n21937);
  nand U22962(n21937,n21938,n21939);
  nor U22963(n21915,n19961,n21796);
  not U22964(n19961,n19696);
  nand U22965(n19696,n21940,n21941,n21942,n21943);
  nand U22966(n21943,n20437,n21801);
  xor U22967(n20437,n21875,G36202);
  not U22968(n21875,n21944);
  nand U22969(n21942,G36126,n21697);
  nand U22970(n21941,G36094,n21698);
  nand U22971(n21940,G36062,n21696);
  nand U22972(n21913,G36125,n19783);
  nand U22973(n21912,n21737,n21945);
  nand U22974(G1491,n21946,n21947,n21948,n21949);
  nor U22975(n21949,n21950,n21951,n21952,n21953);
  nor U22976(n21953,n20342,n21714);
  and U22977(n21952,n19998,n21715);
  xor U22978(n19998,n21930,n21954);
  and U22979(n21954,n21929,n21927);
  nand U22980(n21927,n21955,n21956);
  or U22981(n21929,n21955,n21956);
  nand U22982(n21956,n21957,n21958,n21720);
  nand U22983(n21958,n19999,n21773);
  nand U22984(n21957,n19702,n21774);
  xor U22985(n21955,n21959,n21776);
  nand U22986(n21959,n21960,n21732,n21961);
  nand U22987(n21961,n21773,n19702);
  nand U22988(n21960,n19999,n21779);
  nand U22989(n21930,n21962,n21963);
  nand U22990(n21963,n21964,n21965);
  nor U22991(n21951,n20723,n21784);
  xor U22992(n20723,n21939,n21966);
  and U22993(n21966,n21967,n21936,n21938);
  nand U22994(n21938,n19702,n21787,n20342);
  not U22995(n20342,n19999);
  nand U22996(n21936,n19999,n21788,n21968);
  nand U22997(n21968,n19702,n21787);
  nand U22998(n19999,n21969,n21970);
  nand U22999(n21970,n21669,n18182);
  nand U23000(n21969,n21670,G36421);
  nand U23001(n21967,n19702,n20819);
  nand U23002(n21939,n21971,n21972);
  nand U23003(n21972,n21973,n21974);
  nor U23004(n21950,n19973,n21796);
  not U23005(n19973,n19699);
  nand U23006(n19699,n21975,n21976,n21977,n21978);
  nand U23007(n21978,n21945,n21801);
  not U23008(n21945,n20477);
  nand U23009(n20477,n21979,n21944);
  nand U23010(n21944,G36198,n21980,G36211);
  nand U23011(n21979,n21981,n21982);
  nand U23012(n21982,G36211,n21980);
  not U23013(n21980,n21983);
  not U23014(n21981,G36198);
  nand U23015(n21977,G36125,n21697);
  nand U23016(n21976,G36093,n21698);
  nand U23017(n21975,G36061,n21696);
  nand U23018(n21948,G36124,n19783);
  nand U23019(n21947,n21737,n21984);
  nand U23020(G1490,n21985,n21986,n21987,n21988);
  nor U23021(n21988,n21989,n21990,n21991,n21992);
  nor U23022(n21992,n20537,n21714);
  and U23023(n21991,n20010,n21715);
  xor U23024(n20010,n21965,n21993);
  and U23025(n21993,n21964,n21962);
  nand U23026(n21962,n21994,n21995);
  or U23027(n21964,n21994,n21995);
  nand U23028(n21995,n21996,n21997,n21720);
  nand U23029(n21997,n20011,n21773);
  nand U23030(n21996,n19705,n21774);
  xor U23031(n21994,n21998,n21776);
  nand U23032(n21998,n21999,n21732,n22000);
  nand U23033(n22000,n21773,n19705);
  nand U23034(n21999,n20011,n21779);
  nand U23035(n21965,n22001,n22002);
  nand U23036(n22002,n22003,n22004);
  nor U23037(n21990,n20727,n21784);
  xor U23038(n20727,n21974,n22005);
  and U23039(n22005,n22006,n21971,n21973);
  nand U23040(n21973,n19705,n21787,n20537);
  not U23041(n20537,n20011);
  nand U23042(n21971,n20011,n21788,n22007);
  nand U23043(n22007,n19705,n21787);
  nand U23044(n20011,n22008,n22009);
  nand U23045(n22009,n21669,n18224);
  nand U23046(n22008,n21670,G36420);
  nand U23047(n22006,n19705,n20819);
  nand U23048(n21974,n22010,n22011);
  nand U23049(n22011,n22012,n22013);
  nor U23050(n21989,n19985,n21796);
  not U23051(n19985,n19702);
  nand U23052(n19702,n22014,n22015,n22016,n22017);
  nand U23053(n22017,n21984,n21801);
  not U23054(n21984,n20341);
  xor U23055(n20341,n21983,G36211);
  nand U23056(n22016,G36124,n21697);
  nand U23057(n22015,G36092,n21698);
  nand U23058(n22014,G36060,n21696);
  nand U23059(n21987,G36123,n19783);
  nand U23060(n21986,n21737,n22018);
  nand U23061(G1489,n22019,n22020,n22021,n22022);
  nor U23062(n22022,n22023,n22024,n22025,n22026);
  nor U23063(n22026,n20417,n21714);
  and U23064(n22025,n20022,n21715);
  xor U23065(n20022,n22004,n22027);
  and U23066(n22027,n22003,n22001);
  nand U23067(n22001,n22028,n22029);
  or U23068(n22003,n22028,n22029);
  nand U23069(n22029,n22030,n22031,n21720);
  nand U23070(n22031,n20023,n21773);
  nand U23071(n22030,n19708,n21774);
  xor U23072(n22028,n22032,n21776);
  nand U23073(n22032,n22033,n21732,n22034);
  nand U23074(n22034,n21773,n19708);
  nand U23075(n22033,n20023,n21779);
  nand U23076(n22004,n22035,n22036);
  nand U23077(n22036,n22037,n22038);
  nor U23078(n22024,n20731,n21784);
  xor U23079(n20731,n22013,n22039);
  and U23080(n22039,n22040,n22010,n22012);
  nand U23081(n22012,n19708,n21787,n20417);
  not U23082(n20417,n20023);
  nand U23083(n22010,n20023,n21788,n22041);
  nand U23084(n22041,n19708,n21787);
  nand U23085(n20023,n22042,n22043);
  nand U23086(n22043,n21669,n18261);
  nand U23087(n22042,n21670,G36419);
  nand U23088(n22040,n19708,n20819);
  nand U23089(n22013,n22044,n22045);
  nand U23090(n22045,n22046,n22047);
  nor U23091(n22023,n19997,n21796);
  not U23092(n19997,n19705);
  nand U23093(n19705,n22048,n22049,n22050,n22051);
  nand U23094(n22051,n22018,n21801);
  not U23095(n22018,n20536);
  nand U23096(n20536,n22052,n21983);
  nand U23097(n21983,G36192,n22053,G36204);
  nand U23098(n22052,n22054,n22055);
  nand U23099(n22055,G36204,n22053);
  not U23100(n22054,G36192);
  nand U23101(n22050,G36123,n21697);
  nand U23102(n22049,G36091,n21698);
  nand U23103(n22048,G36059,n21696);
  nand U23104(n22021,G36122,n19783);
  nand U23105(n22020,n21737,n22056);
  nand U23106(G1488,n22057,n22058,n22059,n22060);
  nor U23107(n22060,n22061,n22062,n22063,n22064);
  nor U23108(n22064,n20517,n21714);
  and U23109(n22063,n20034,n21715);
  xor U23110(n20034,n22038,n22065);
  and U23111(n22065,n22037,n22035);
  nand U23112(n22035,n22066,n22067);
  or U23113(n22037,n22066,n22067);
  nand U23114(n22067,n22068,n22069,n21720);
  nand U23115(n22069,n20035,n21773);
  nand U23116(n22068,n19711,n21774);
  xor U23117(n22066,n22070,n21776);
  nand U23118(n22070,n22071,n21732,n22072);
  nand U23119(n22072,n21773,n19711);
  nand U23120(n22071,n20035,n21779);
  nand U23121(n22038,n22073,n22074);
  nand U23122(n22074,n22075,n22076);
  nor U23123(n22062,n20735,n21784);
  xor U23124(n20735,n22047,n22077);
  and U23125(n22077,n22078,n22044,n22046);
  nand U23126(n22046,n19711,n21787,n20517);
  not U23127(n20517,n20035);
  nand U23128(n22044,n20035,n21788,n22079);
  nand U23129(n22079,n19711,n21787);
  nand U23130(n20035,n22080,n22081);
  nand U23131(n22081,n21669,n18301);
  nand U23132(n22080,n21670,G36418);
  nand U23133(n22078,n19711,n20819);
  nand U23134(n22047,n22082,n22083);
  nand U23135(n22083,n22084,n22085);
  nor U23136(n22061,n20009,n21796);
  not U23137(n20009,n19708);
  nand U23138(n19708,n22086,n22087,n22088,n22089);
  nand U23139(n22089,n22056,n21801);
  not U23140(n22056,n20416);
  xnor U23141(n20416,n22053,G36204);
  nand U23142(n22088,G36122,n21697);
  nand U23143(n22087,G36090,n21698);
  nand U23144(n22086,G36058,n21696);
  nand U23145(n22059,G36121,n19783);
  nand U23146(n22058,n21737,n20516);
  nand U23147(G1487,n22090,n22091,n22092,n22093);
  nor U23148(n22093,n22094,n22095,n22096,n22097);
  nor U23149(n22097,n20377,n21714);
  and U23150(n22096,n20046,n21715);
  xor U23151(n20046,n22076,n22098);
  and U23152(n22098,n22075,n22073);
  nand U23153(n22073,n22099,n22100);
  or U23154(n22075,n22099,n22100);
  nand U23155(n22100,n22101,n22102,n21720);
  and U23156(n21720,n22103,n22104);
  nand U23157(n22103,n22106,G36120);
  nand U23158(n22102,n20047,n21773);
  nand U23159(n22101,n19714,n21774);
  xor U23160(n22099,n22107,n21776);
  nand U23161(n22107,n22108,n21732,n22109);
  nand U23162(n22109,n21773,n19714);
  nand U23163(n21732,n20644,n22110);
  nand U23164(n22108,n20047,n21779);
  nand U23165(n22076,n22111,n22112);
  nand U23166(n22112,n22113,n22114);
  nor U23167(n22095,n20739,n21784);
  xor U23168(n20739,n22085,n22115);
  and U23169(n22115,n22116,n22082,n22084);
  nand U23170(n22084,n19714,n21787,n20377);
  not U23171(n20377,n20047);
  nand U23172(n22082,n20047,n21788,n22117);
  nand U23173(n22117,n19714,n21787);
  nand U23174(n20047,n22118,n22119,n22120);
  nand U23175(n22120,n21691,n20644);
  nand U23176(n22119,n21669,n18353);
  nand U23177(n22118,n21670,G36417);
  nand U23178(n22116,n19714,n20819);
  nand U23179(n22085,n22121,n22122);
  nand U23180(n22122,n22123,n22124);
  nor U23181(n22094,n20021,n21796);
  not U23182(n20021,n19711);
  nand U23183(n19711,n22125,n22126,n22127,n22128);
  nand U23184(n22128,n20516,n21801);
  nor U23185(n20516,n22129,n22053);
  nor U23186(n22053,n22130,n22131,n21534);
  and U23187(n22129,n22130,n22132);
  or U23188(n22132,n21534,n22131);
  not U23189(n21534,G36208);
  not U23190(n22130,G36194);
  nand U23191(n22127,G36121,n21697);
  nand U23192(n22126,G36089,n21698);
  nand U23193(n22125,G36057,n21696);
  nand U23194(n22092,G36120,n19783);
  nand U23195(n22091,n21737,n22133);
  nand U23196(G1486,n22134,n22135,n22136,n22137);
  nor U23197(n22137,n22138,n22139,n22140,n22141);
  nor U23198(n22141,n20566,n21714);
  and U23199(n22140,n20058,n21715);
  xor U23200(n20058,n22114,n22142);
  and U23201(n22142,n22113,n22111);
  nand U23202(n22111,n22143,n22144);
  or U23203(n22113,n22143,n22144);
  nand U23204(n22144,n22145,n22146,n22147,n22148);
  nand U23205(n22148,n20059,n21773);
  nand U23206(n22147,n19717,n21774);
  nand U23207(n22145,n22106,G36119);
  xor U23208(n22143,n22149,n21776);
  nand U23209(n22149,n22150,n22151,n22152);
  nand U23210(n22152,n21773,n19717);
  nand U23211(n22151,n20059,n21779);
  nand U23212(n22150,n21527,n22110);
  nand U23213(n22114,n22153,n22154);
  nand U23214(n22154,n22155,n22156);
  nor U23215(n22139,n20743,n21784);
  xor U23216(n20743,n22124,n22157);
  and U23217(n22157,n22158,n22121,n22123);
  nand U23218(n22123,n19717,n21787,n20566);
  not U23219(n20566,n20059);
  nand U23220(n22121,n20059,n21788,n22159);
  nand U23221(n22159,n19717,n21787);
  nand U23222(n20059,n22160,n22161,n22162);
  nand U23223(n22162,n21527,n21691);
  not U23224(n21527,n21526);
  nand U23225(n21526,n22163,n22164);
  or U23226(n22164,G35991,G36004);
  nand U23227(n22163,G36004,n22165);
  nand U23228(n22165,n22166,n22167);
  nand U23229(n22161,n21669,n18410);
  nand U23230(n22160,n21670,G36416);
  nand U23231(n22158,n19717,n20819);
  nand U23232(n22124,n22168,n22169);
  nand U23233(n22169,n22170,n22171);
  nor U23234(n22138,n20033,n21796);
  not U23235(n20033,n19714);
  nand U23236(n19714,n22172,n22173,n22174,n22175);
  nand U23237(n22175,n22133,n21801);
  not U23238(n22133,n20376);
  xor U23239(n20376,n22131,G36208);
  nand U23240(n22174,G36120,n21697);
  nand U23241(n22173,G36088,n21698);
  nand U23242(n22172,G36056,n21696);
  nand U23243(n22136,G36119,n19783);
  nand U23244(n22135,n21737,n22176);
  nand U23245(G1485,n22177,n22178,n22179,n22180);
  nor U23246(n22180,n22181,n22182,n22183,n22184);
  nor U23247(n22184,n20468,n21714);
  and U23248(n22183,n20070,n21715);
  xor U23249(n20070,n22156,n22185);
  and U23250(n22185,n22155,n22153);
  nand U23251(n22153,n22186,n22187);
  or U23252(n22155,n22186,n22187);
  nand U23253(n22187,n22188,n22189,n22190,n22191);
  nand U23254(n22191,n20071,n21773);
  nand U23255(n22190,n19720,n21774);
  nand U23256(n22188,n22106,G36118);
  xor U23257(n22186,n22192,n21776);
  nand U23258(n22192,n22193,n22194,n22195);
  nand U23259(n22195,n21773,n19720);
  nand U23260(n22194,n20071,n21779);
  nand U23261(n22193,n21513,n22110);
  nand U23262(n22156,n22196,n22197);
  nand U23263(n22197,n22198,n22199);
  nor U23264(n22182,n20747,n21784);
  xor U23265(n20747,n22171,n22200);
  and U23266(n22200,n22201,n22168,n22170);
  nand U23267(n22170,n19720,n21787,n20468);
  not U23268(n20468,n20071);
  nand U23269(n22168,n20071,n21788,n22202);
  nand U23270(n22202,n19720,n21787);
  nand U23271(n20071,n22203,n22204,n22205);
  nand U23272(n22205,n21513,n21691);
  and U23273(n21513,n22206,n22207);
  nand U23274(n22207,n22208,n22209);
  nand U23275(n22206,G36004,n22210);
  nand U23276(n22210,n22211,n22212);
  nand U23277(n22204,n21669,n18461);
  nand U23278(n22203,n21670,G36415);
  nand U23279(n22201,n19720,n20819);
  nand U23280(n22171,n22213,n22214);
  nand U23281(n22214,n22215,n22216);
  nor U23282(n22181,n20045,n21796);
  not U23283(n20045,n19717);
  nand U23284(n19717,n22217,n22218,n22219,n22220);
  nand U23285(n22220,n22176,n21801);
  not U23286(n22176,n20565);
  nand U23287(n20565,n22221,n22131);
  nand U23288(n22131,G36189,n22222,G36199);
  nand U23289(n22221,n21520,n22223);
  nand U23290(n22223,G36199,n22222);
  not U23291(n22222,n22224);
  not U23292(n21520,G36189);
  nand U23293(n22219,G36119,n21697);
  nand U23294(n22218,G36087,n21698);
  nand U23295(n22217,G36055,n21696);
  nand U23296(n22179,G36118,n19783);
  nand U23297(n22178,n21737,n22225);
  nand U23298(n22177,n19782,n19723);
  nand U23299(G1484,n22226,n22227,n22228,n22229);
  nor U23300(n22229,n22230,n22231,n22232,n22233);
  nor U23301(n22233,n20448,n21714);
  and U23302(n22232,n20082,n21715);
  xor U23303(n20082,n22199,n22234);
  and U23304(n22234,n22198,n22196);
  nand U23305(n22196,n22235,n22236);
  or U23306(n22198,n22235,n22236);
  nand U23307(n22236,n22237,n22238,n22239,n22240);
  nand U23308(n22240,n20083,n21773);
  nand U23309(n22239,n19723,n21774);
  nand U23310(n22237,n22106,G36117);
  xor U23311(n22235,n22241,n21776);
  nand U23312(n22241,n22242,n22243,n22244);
  nand U23313(n22244,n21773,n19723);
  nand U23314(n22243,n20083,n21779);
  nand U23315(n22242,n21501,n22110);
  nand U23316(n22199,n22245,n22246);
  nand U23317(n22246,n22247,n22248);
  nor U23318(n22231,n20751,n21784);
  xor U23319(n20751,n22216,n22249);
  and U23320(n22249,n22250,n22213,n22215);
  nand U23321(n22215,n19723,n21787,n20448);
  not U23322(n20448,n20083);
  nand U23323(n22213,n20083,n21788,n22251);
  nand U23324(n22251,n19723,n21787);
  nand U23325(n20083,n22252,n22253,n22254);
  nand U23326(n22254,n21501,n21691);
  and U23327(n21501,n22255,n22256);
  nand U23328(n22256,n22257,n22209);
  nand U23329(n22255,n22258,G36004);
  nand U23330(n22253,n21669,n18518);
  nand U23331(n22252,n21670,G36414);
  nand U23332(n22250,n19723,n20819);
  nand U23333(n22216,n22259,n22260);
  nand U23334(n22260,n22261,n22262);
  nor U23335(n22230,n20057,n21796);
  not U23336(n20057,n19720);
  nand U23337(n19720,n22263,n22264,n22265,n22266);
  nand U23338(n22266,n22225,n21801);
  not U23339(n22225,n20467);
  xor U23340(n20467,n22224,G36199);
  nand U23341(n22265,G36118,n21697);
  nand U23342(n22264,G36086,n21698);
  nand U23343(n22263,G36054,n21696);
  nand U23344(n22228,G36117,n19783);
  nand U23345(n22227,n21737,n22267);
  nand U23346(n22226,n19782,n19726);
  nand U23347(G1483,n22268,n22269,n22270,n22271);
  nor U23348(n22271,n22272,n22273,n22274,n22275);
  nor U23349(n22275,n20613,n21714);
  and U23350(n22274,n20094,n21715);
  xor U23351(n20094,n22248,n22276);
  and U23352(n22276,n22247,n22245);
  nand U23353(n22245,n22277,n22278);
  or U23354(n22247,n22277,n22278);
  nand U23355(n22278,n22279,n22280,n22281,n22282);
  nand U23356(n22282,n20095,n21773);
  nand U23357(n22281,n19726,n21774);
  nand U23358(n22279,n22106,G36116);
  xor U23359(n22277,n22283,n21776);
  nand U23360(n22283,n22284,n22285,n22286);
  nand U23361(n22286,n21773,n19726);
  nand U23362(n22285,n20095,n21779);
  nand U23363(n22284,n21488,n22110);
  nand U23364(n22248,n22287,n22288);
  nand U23365(n22288,n22289,n22290);
  nor U23366(n22273,n20755,n21784);
  xor U23367(n20755,n22262,n22291);
  and U23368(n22291,n22292,n22259,n22261);
  nand U23369(n22261,n19726,n21787,n20613);
  not U23370(n20613,n20095);
  nand U23371(n22259,n20095,n21788,n22293);
  nand U23372(n22293,n19726,n21787);
  nand U23373(n20095,n22294,n22295,n22296);
  nand U23374(n22296,n21488,n21691);
  not U23375(n21488,n21639);
  nand U23376(n21639,n22297,n22298);
  or U23377(n22298,G35988,G36004);
  nand U23378(n22297,n22299,G36004);
  nand U23379(n22295,n21669,n18568);
  nand U23380(n22294,n21670,G36413);
  nand U23381(n22292,n19726,n20819);
  nand U23382(n22262,n22300,n22301);
  nand U23383(n22301,n22302,n22303);
  nor U23384(n22272,n20069,n21796);
  not U23385(n20069,n19723);
  nand U23386(n19723,n22304,n22305,n22306,n22307);
  nand U23387(n22307,n22267,n21801);
  not U23388(n22267,n20447);
  nand U23389(n20447,n22308,n22224);
  nand U23390(n22224,G36186,n22309,G36201);
  nand U23391(n22308,n21495,n22310);
  nand U23392(n22310,G36186,n22309);
  not U23393(n22309,n22311);
  not U23394(n21495,G36201);
  nand U23395(n22306,G36117,n21697);
  nand U23396(n22305,G36085,n21698);
  nand U23397(n22304,G36053,n21696);
  nand U23398(n22270,G36116,n19783);
  nand U23399(n22269,n21737,n22312);
  nand U23400(n22268,n19782,n19729);
  nand U23401(G1482,n22313,n22314,n22315,n22316);
  nor U23402(n22316,n22317,n22318,n22319,n22320);
  nor U23403(n22320,n20332,n21714);
  and U23404(n22319,n20106,n21715);
  xor U23405(n20106,n22290,n22321);
  and U23406(n22321,n22287,n22289);
  or U23407(n22289,n22322,n22323);
  nand U23408(n22287,n22322,n22323);
  nand U23409(n22323,n22324,n22325,n22326,n22327);
  nand U23410(n22327,n20107,n21773);
  nand U23411(n22326,n19729,n21774);
  nand U23412(n22324,n22106,G36115);
  xor U23413(n22322,n22328,n21776);
  nand U23414(n22328,n22329,n22330,n22331);
  nand U23415(n22331,n21773,n19729);
  nand U23416(n22330,n20107,n21779);
  nand U23417(n22329,n21475,n22110);
  nand U23418(n22290,n22332,n22333);
  nand U23419(n22333,n22334,n22335);
  nor U23420(n22318,n20759,n21784);
  xor U23421(n20759,n22303,n22336);
  and U23422(n22336,n22337,n22300,n22302);
  nand U23423(n22302,n19729,n21787,n20332);
  not U23424(n20332,n20107);
  nand U23425(n22300,n20107,n21788,n22338);
  nand U23426(n22338,n19729,n21787);
  nand U23427(n20107,n22339,n22340,n22341);
  nand U23428(n22341,n21475,n21691);
  not U23429(n21475,n21563);
  nand U23430(n21563,n22342,n22343);
  or U23431(n22343,G35987,G36004);
  nand U23432(n22342,G36004,n22344);
  nand U23433(n22344,n22345,n22346);
  nand U23434(n22340,n21669,n18626);
  nand U23435(n22339,n21670,G36412);
  nand U23436(n22337,n19729,n20819);
  nand U23437(n22303,n22347,n22348);
  nand U23438(n22348,n22349,n22350);
  nor U23439(n22317,n20081,n21796);
  not U23440(n20081,n19726);
  nand U23441(n19726,n22351,n22352,n22353,n22354);
  nand U23442(n22354,n22312,n21801);
  not U23443(n22312,n20599);
  xor U23444(n20599,n22311,G36186);
  nand U23445(n22353,G36116,n21697);
  nand U23446(n22352,G36084,n21698);
  nand U23447(n22351,G36052,n21696);
  nand U23448(n22315,G36115,n19783);
  nand U23449(n22314,n21737,n22355);
  nand U23450(n22313,n19782,n19732);
  nand U23451(G1481,n22356,n22357,n22358,n22359);
  nor U23452(n22359,n22360,n22361,n22362,n22363);
  nor U23453(n22363,n20527,n21714);
  and U23454(n22362,n20118,n21715);
  xor U23455(n20118,n22335,n22364);
  and U23456(n22364,n22334,n22332);
  nand U23457(n22332,n22365,n22366);
  or U23458(n22334,n22365,n22366);
  nand U23459(n22366,n22367,n22368,n22369,n22370);
  nand U23460(n22370,n20119,n21773);
  nand U23461(n22369,n19732,n21774);
  nand U23462(n22367,n22106,G36114);
  xor U23463(n22365,n22371,n21776);
  nand U23464(n22371,n22372,n22373,n22374);
  nand U23465(n22374,n21773,n19732);
  nand U23466(n22373,n20119,n21779);
  nand U23467(n22372,n21456,n22110);
  nand U23468(n22335,n22375,n22376);
  nand U23469(n22376,n22377,n22378);
  nor U23470(n22361,n20763,n21784);
  xor U23471(n20763,n22350,n22379);
  and U23472(n22379,n22380,n22347,n22349);
  nand U23473(n22349,n19732,n21787,n20527);
  not U23474(n20527,n20119);
  nand U23475(n22347,n20119,n21788,n22381);
  nand U23476(n22381,n19732,n21787);
  nand U23477(n20119,n22382,n22383,n22384);
  nand U23478(n22384,n21456,n21691);
  not U23479(n21456,n21455);
  nand U23480(n21455,n22385,n22386);
  or U23481(n22386,G35986,G36004);
  nand U23482(n22385,G36004,n22387);
  nand U23483(n22387,n22388,n22389);
  nand U23484(n22383,n21669,n18678);
  nand U23485(n22382,n21670,G36411);
  nand U23486(n22380,n19732,n20819);
  nand U23487(n22350,n22390,n22391);
  nand U23488(n22391,n22392,n22393);
  or U23489(n22392,n20131,n22394);
  nor U23490(n22360,n20093,n21796);
  not U23491(n20093,n19729);
  nand U23492(n19729,n22395,n22396,n22397,n22398);
  nand U23493(n22398,n22355,n21801);
  not U23494(n22355,n20331);
  nand U23495(n20331,n22399,n22311);
  nand U23496(n22311,G36193,n22400,G36212);
  nand U23497(n22399,n21463,n22401);
  nand U23498(n22401,G36193,n22400);
  not U23499(n22400,n22402);
  not U23500(n21463,G36212);
  nand U23501(n22397,G36115,n21697);
  nand U23502(n22396,G36083,n21698);
  nand U23503(n22395,G36051,n21696);
  nand U23504(n22358,G36114,n19783);
  nand U23505(n22357,n21737,n22403);
  nand U23506(n22356,n19782,n19735);
  nand U23507(G1480,n22404,n22405,n22406,n22407);
  nor U23508(n22407,n22408,n22409,n22410,n22411);
  nor U23509(n22411,n20427,n21714);
  and U23510(n22410,n20130,n21715);
  xor U23511(n20130,n22378,n22412);
  and U23512(n22412,n22377,n22375);
  nand U23513(n22375,n22413,n22414);
  or U23514(n22377,n22413,n22414);
  nand U23515(n22414,n22415,n22416,n22417,n22418);
  nand U23516(n22418,n20131,n21773);
  nand U23517(n22417,n19735,n21774);
  nand U23518(n22416,n22105,G36081);
  nand U23519(n22415,n22106,G36113);
  xor U23520(n22413,n22419,n21776);
  nand U23521(n22419,n22420,n22421,n22422);
  nand U23522(n22422,n21773,n19735);
  nand U23523(n22421,n20131,n21779);
  nand U23524(n22420,n21443,n22110);
  nand U23525(n22378,n22423,n22424);
  nand U23526(n22424,n22425,n22426);
  nor U23527(n22409,n20767,n21784);
  xor U23528(n20767,n22393,n22427);
  nor U23529(n22427,n22428,n22429);
  nor U23530(n22429,n22430,n22394);
  nor U23531(n22430,n22431,n20427);
  not U23532(n20427,n20131);
  not U23533(n22428,n22390);
  nand U23534(n22390,n20131,n21788,n22394);
  nand U23535(n22394,n21787,n19735);
  nand U23536(n20131,n22432,n22433,n22434);
  nand U23537(n22434,n21443,n21691);
  not U23538(n21443,n21570);
  nand U23539(n21570,n22435,n22436,n22437);
  nand U23540(n22436,n22438,n22209);
  nand U23541(n22435,G35985,n22439,G36004);
  nand U23542(n22433,n21669,n18738);
  nand U23543(n22432,n21670,G36410);
  nand U23544(n22393,n22440,n22441);
  nand U23545(n22441,n22442,n22443);
  or U23546(n22442,n20143,n22444);
  nor U23547(n22408,n20105,n21796);
  not U23548(n20105,n19732);
  nand U23549(n19732,n22445,n22446,n22447,n22448);
  nand U23550(n22448,n22403,n21801);
  not U23551(n22403,n20526);
  xor U23552(n20526,n22402,G36193);
  nand U23553(n22447,G36114,n21697);
  nand U23554(n22446,G36082,n21698);
  nand U23555(n22445,G36050,n21696);
  nand U23556(n22406,G36113,n19783);
  nand U23557(n22405,n21737,n22449);
  nand U23558(n22404,n19782,n19738);
  nand U23559(G1479,n22450,n22451,n22452,n22453);
  nor U23560(n22453,n22454,n22455,n22456,n22457);
  nor U23561(n22457,n20547,n21714);
  and U23562(n22456,n20142,n21715);
  xor U23563(n20142,n22426,n22458);
  and U23564(n22458,n22425,n22423);
  nand U23565(n22423,n22459,n22460);
  or U23566(n22425,n22459,n22460);
  nand U23567(n22460,n22461,n22462,n22463,n22464);
  nand U23568(n22464,n20143,n21773);
  nand U23569(n22463,n19738,n21774);
  nand U23570(n22462,n22105,G36080);
  nand U23571(n22461,n22106,G36112);
  xor U23572(n22459,n22465,n21776);
  nand U23573(n22465,n22466,n22467,n22468);
  nand U23574(n22468,n21773,n19738);
  nand U23575(n22467,n20143,n21779);
  nand U23576(n22466,n21431,n22110);
  nand U23577(n22426,n22469,n22470);
  nand U23578(n22470,n22471,n22472);
  nor U23579(n22455,n20771,n21784);
  xor U23580(n20771,n22443,n22473);
  nor U23581(n22473,n22474,n22475);
  nor U23582(n22475,n22476,n22444);
  nor U23583(n22476,n22431,n20547);
  not U23584(n20547,n20143);
  not U23585(n22474,n22440);
  nand U23586(n22440,n20143,n21788,n22444);
  nand U23587(n22444,n21787,n19738);
  nand U23588(n20143,n22477,n22478,n22479);
  nand U23589(n22479,n21431,n21691);
  not U23590(n21431,n21430);
  nand U23591(n21430,n22480,n22481,n22439);
  nand U23592(n22481,n22482,n22209);
  nand U23593(n22480,G35984,n22483,G36004);
  nand U23594(n22478,n21669,n18791);
  nand U23595(n22477,n21670,G36409);
  nand U23596(n22443,n22484,n22485);
  nand U23597(n22485,n22486,n22487);
  nor U23598(n22454,n20117,n21796);
  not U23599(n20117,n19735);
  nand U23600(n19735,n22488,n22489,n22490,n22491);
  nand U23601(n22491,n22449,n21801);
  not U23602(n22449,n20426);
  nand U23603(n20426,n22492,n22402);
  nand U23604(n22402,G36191,n22493,G36203);
  nand U23605(n22492,n21438,n22494);
  nand U23606(n22494,G36191,n22493);
  not U23607(n21438,G36203);
  nand U23608(n22490,G36113,n21697);
  nand U23609(n22489,G36081,n21698);
  nand U23610(n22488,G36049,n21696);
  nand U23611(n22452,G36112,n19783);
  nand U23612(n22451,n21737,n22495);
  nand U23613(n22450,n19782,n19741);
  nand U23614(G1478,n22496,n22497,n22498,n22499);
  nor U23615(n22499,n22500,n22501,n22502,n22503);
  nor U23616(n22503,n20353,n21714);
  and U23617(n22502,n20154,n21715);
  xor U23618(n20154,n22471,n22504);
  and U23619(n22504,n22469,n22472);
  or U23620(n22472,n22505,n22506);
  nand U23621(n22469,n22505,n22506);
  nand U23622(n22506,n22507,n22508,n22509,n22510);
  nand U23623(n22510,n20155,n21773);
  nand U23624(n22509,n19741,n21774);
  nand U23625(n22508,n22105,G36079);
  nand U23626(n22507,n22106,G36111);
  xor U23627(n22505,n22511,n21776);
  nand U23628(n22511,n22512,n22513,n22514);
  nand U23629(n22514,n21773,n19741);
  nand U23630(n22513,n20155,n21779);
  nand U23631(n22512,n21419,n22110);
  nand U23632(n22471,n22515,n22516);
  nand U23633(n22516,n22517,n22518);
  nor U23634(n22501,n20775,n21784);
  xor U23635(n20775,n22487,n22519);
  and U23636(n22519,n22520,n22484,n22486);
  nand U23637(n22486,n19741,n21787,n20353);
  not U23638(n20353,n20155);
  nand U23639(n22484,n20155,n21788,n22521);
  nand U23640(n22521,n19741,n21787);
  nand U23641(n20155,n22522,n22523,n22524);
  nand U23642(n22524,n21419,n21691);
  not U23643(n21419,n21577);
  nand U23644(n21577,n22525,n22526);
  or U23645(n22526,G35983,G36004);
  nand U23646(n22525,G36004,n22527);
  nand U23647(n22523,n21669,n18843);
  nand U23648(n22522,n21670,G36408);
  nand U23649(n22520,n19741,n20819);
  nand U23650(n22487,n22528,n22529);
  nand U23651(n22529,n22530,n22531);
  or U23652(n22530,n20167,n22532);
  nor U23653(n22500,n20129,n21796);
  not U23654(n20129,n19738);
  nand U23655(n19738,n22533,n22534,n22535,n22536);
  nand U23656(n22536,n22495,n21801);
  not U23657(n22495,n20546);
  xnor U23658(n20546,G36191,n22493);
  nand U23659(n22535,G36112,n21697);
  nand U23660(n22534,G36080,n21698);
  nand U23661(n22533,G36048,n21696);
  nand U23662(n22498,G36111,n19783);
  nand U23663(n22497,n21737,n20352);
  nand U23664(n22496,n19782,n19744);
  nand U23665(G1477,n22537,n22538,n22539,n22540);
  nor U23666(n22540,n22541,n22542,n22543,n22544);
  nor U23667(n22544,n20498,n21714);
  and U23668(n22543,n20166,n21715);
  xor U23669(n20166,n22518,n22545);
  and U23670(n22545,n22517,n22515);
  nand U23671(n22515,n22546,n22547);
  or U23672(n22517,n22546,n22547);
  nand U23673(n22547,n22548,n22549,n22550,n22551);
  nand U23674(n22551,n20167,n21773);
  nand U23675(n22550,n19744,n21774);
  nand U23676(n22549,n22105,G36078);
  nand U23677(n22548,n22106,G36110);
  xor U23678(n22546,n21728,n22552);
  and U23679(n22552,n22553,n22554,n22555);
  nand U23680(n22555,n21773,n19744);
  nand U23681(n22554,n20167,n21779);
  nand U23682(n22553,n21400,n22110);
  nand U23683(n22518,n22556,n22557);
  nand U23684(n22557,n22558,n22559);
  nor U23685(n22542,n20779,n21784);
  xor U23686(n20779,n22531,n22560);
  nor U23687(n22560,n22561,n22562);
  nor U23688(n22562,n22563,n22532);
  nor U23689(n22563,n22431,n20498);
  not U23690(n20498,n20167);
  not U23691(n22561,n22528);
  nand U23692(n22528,n20167,n21788,n22532);
  nand U23693(n22532,n21787,n19744);
  nand U23694(n20167,n22564,n22565,n22566);
  nand U23695(n22566,n21400,n21691);
  not U23696(n21400,n21581);
  nand U23697(n21581,n22567,n22568,n22569);
  nand U23698(n22568,n22570,n22209);
  nand U23699(n22567,G35982,n22571,G36004);
  nand U23700(n22565,n21669,n18898);
  nand U23701(n22564,n21670,G36407);
  nand U23702(n22531,n22572,n22573);
  nand U23703(n22573,n22574,n22575);
  or U23704(n22574,n20179,n22576);
  nor U23705(n22541,n20141,n21796);
  not U23706(n20141,n19741);
  nand U23707(n19741,n22577,n22578,n22579,n22580);
  nand U23708(n22580,n20352,n21801);
  nor U23709(n20352,n22493,n22581);
  and U23710(n22581,n22582,n21407);
  nor U23711(n22493,n21407,n22582);
  not U23712(n21407,G36210);
  nand U23713(n22579,G36111,n21697);
  nand U23714(n22578,G36079,n21698);
  nand U23715(n22577,G36047,n21696);
  nand U23716(n22539,G36110,n19783);
  nand U23717(n22538,n21737,n22583);
  nand U23718(n22537,n19782,n19747);
  nand U23719(G1476,n22584,n22585,n22586,n22587);
  nor U23720(n22587,n22588,n22589,n22590,n22591);
  nor U23721(n22591,n20398,n21714);
  and U23722(n22590,n20178,n21715);
  xor U23723(n20178,n22559,n22592);
  and U23724(n22592,n22558,n22556);
  nand U23725(n22556,n22593,n22594);
  or U23726(n22558,n22593,n22594);
  nand U23727(n22594,n22595,n22596,n22597,n22598);
  nand U23728(n22598,n20179,n21773);
  nand U23729(n22597,n19747,n21774);
  nand U23730(n22596,n22105,G36077);
  nand U23731(n22595,n22106,G36109);
  xor U23732(n22593,n21728,n22599);
  and U23733(n22599,n22600,n22601,n22602);
  nand U23734(n22602,n21773,n19747);
  nand U23735(n22601,n20179,n21779);
  nand U23736(n22600,n21387,n22110);
  nand U23737(n22559,n22603,n22604);
  nand U23738(n22604,n22605,n22606);
  nor U23739(n22589,n20783,n21784);
  xor U23740(n20783,n22575,n22607);
  nor U23741(n22607,n22608,n22609);
  nor U23742(n22609,n22610,n22576);
  nor U23743(n22610,n22431,n20398);
  not U23744(n20398,n20179);
  not U23745(n22608,n22572);
  nand U23746(n22572,n20179,n21788,n22576);
  nand U23747(n22576,n21787,n19747);
  nand U23748(n20179,n22611,n22612,n22613);
  nand U23749(n22613,n21387,n21691);
  not U23750(n21387,n21386);
  nand U23751(n21386,n22614,n22615);
  or U23752(n22615,G35981,G36004);
  nand U23753(n22614,G36004,n22616);
  nand U23754(n22612,n21669,n18946);
  nand U23755(n22611,n21670,G36406);
  nand U23756(n22575,n22617,n22618);
  nand U23757(n22618,n22619,n22620);
  or U23758(n22619,n20191,n22621);
  nor U23759(n22588,n20153,n21796);
  not U23760(n20153,n19744);
  nand U23761(n19744,n22622,n22623,n22624,n22625);
  nand U23762(n22625,n22583,n21801);
  not U23763(n22583,n20497);
  nand U23764(n20497,n22626,n22582);
  or U23765(n22582,n21394,n22627);
  nand U23766(n22626,n21394,n22627);
  nand U23767(n22627,G36206,n22628,G36214);
  not U23768(n21394,G36196);
  nand U23769(n22624,G36110,n21697);
  nand U23770(n22623,G36078,n21698);
  nand U23771(n22622,G36046,n21696);
  nand U23772(n22586,G36109,n19783);
  nand U23773(n22585,n21737,n22629);
  nand U23774(n22584,n19782,n19750);
  nand U23775(G1475,n22630,n22631,n22632,n22633);
  nor U23776(n22633,n22634,n22635,n22636,n22637);
  nor U23777(n22637,n20309,n21714);
  and U23778(n22636,n20190,n21715);
  xor U23779(n20190,n22605,n22638);
  and U23780(n22638,n22603,n22606);
  or U23781(n22606,n22639,n22640);
  nand U23782(n22603,n22639,n22640);
  nand U23783(n22640,n22641,n22642,n22643,n22644);
  nand U23784(n22644,n20191,n21773);
  nand U23785(n22643,n19750,n21774);
  nand U23786(n22642,n22105,G36076);
  nand U23787(n22641,n22106,G36108);
  xor U23788(n22639,n21728,n22645);
  and U23789(n22645,n22646,n22647,n22648);
  nand U23790(n22648,n21773,n19750);
  nand U23791(n22647,n20191,n21779);
  nand U23792(n22646,n21374,n22110);
  nand U23793(n22605,n22649,n22650);
  nand U23794(n22650,n22651,n22652);
  nor U23795(n22635,n20787,n21784);
  xor U23796(n20787,n22620,n22653);
  nor U23797(n22653,n22654,n22655);
  nor U23798(n22655,n22656,n22621);
  nor U23799(n22656,n22431,n20309);
  not U23800(n20309,n20191);
  not U23801(n22654,n22617);
  nand U23802(n22617,n20191,n21788,n22621);
  nand U23803(n22621,n21787,n19750);
  nand U23804(n20191,n22657,n22658,n22659);
  nand U23805(n22659,n21374,n21691);
  not U23806(n21374,n21372);
  nand U23807(n21372,n22660,n22661,n22662);
  nand U23808(n22661,n22663,n22209);
  nand U23809(n22660,G35980,n22664,G36004);
  nand U23810(n22658,n21669,n19002);
  nand U23811(n22657,n21670,G36405);
  nand U23812(n22620,n22665,n22666);
  nand U23813(n22666,n22667,n22668);
  or U23814(n22667,n20203,n22669);
  nor U23815(n22634,n20165,n21796);
  not U23816(n20165,n19747);
  nand U23817(n19747,n22670,n22671,n22672,n22673);
  nand U23818(n22673,n22629,n21801);
  not U23819(n22629,n20397);
  xnor U23820(n20397,G36206,n22674);
  nor U23821(n22674,n22675,n21368);
  not U23822(n21368,G36214);
  nand U23823(n22672,G36109,n21697);
  nand U23824(n22671,G36077,n21698);
  nand U23825(n22670,G36045,n21696);
  nand U23826(n22632,G36108,n19783);
  nand U23827(n22631,n21737,n20308);
  nand U23828(n22630,n19782,n19753);
  nand U23829(G1474,n22676,n22677,n22678,n22679);
  nor U23830(n22679,n22680,n22681,n22682,n22683);
  nor U23831(n22683,n20576,n21714);
  and U23832(n22682,n20202,n21715);
  xor U23833(n20202,n22651,n22684);
  and U23834(n22684,n22649,n22652);
  or U23835(n22652,n22685,n22686);
  nand U23836(n22649,n22685,n22686);
  nand U23837(n22686,n22687,n22688,n22689,n22690);
  nand U23838(n22690,n20203,n21773);
  nand U23839(n22689,n19753,n21774);
  nand U23840(n22688,n22105,G36075);
  nand U23841(n22687,n22106,G36107);
  xor U23842(n22685,n21728,n22691);
  and U23843(n22691,n22692,n22693,n22694);
  nand U23844(n22694,n21773,n19753);
  nand U23845(n22693,n20203,n21779);
  nand U23846(n22692,n21361,n22110);
  nand U23847(n22651,n22695,n22696);
  nand U23848(n22696,n22697,n22698);
  nor U23849(n22681,n20791,n21784);
  xor U23850(n20791,n22668,n22699);
  nor U23851(n22699,n22700,n22701);
  nor U23852(n22701,n22702,n22669);
  nor U23853(n22702,n22431,n20576);
  not U23854(n20576,n20203);
  not U23855(n22700,n22665);
  nand U23856(n22669,n21787,n19753);
  nand U23857(n20203,n22703,n22704,n22705);
  nand U23858(n22705,n21361,n21691);
  not U23859(n21361,n21595);
  nand U23860(n21595,n22706,n22707);
  or U23861(n22707,G35979,G36004);
  nand U23862(n22706,G36004,n22708);
  nand U23863(n22708,n22709,n22664);
  nand U23864(n22704,n21669,n19053);
  nand U23865(n22703,n21670,G36404);
  nand U23866(n22668,n22710,n22711);
  nand U23867(n22711,n22712,n22713);
  or U23868(n22712,n20215,n22714);
  nor U23869(n22680,n20177,n21796);
  not U23870(n20177,n19750);
  nand U23871(n19750,n22715,n22716,n22717,n22718);
  nand U23872(n22718,n20308,n21801);
  xnor U23873(n20308,n22675,G36214);
  nand U23874(n22717,G36108,n21697);
  nand U23875(n22716,G36076,n21698);
  nand U23876(n22715,G36044,n21696);
  nand U23877(n22678,G36107,n19783);
  nand U23878(n22677,n21737,n22719);
  nand U23879(n22676,n19782,n19756);
  nand U23880(G1473,n22720,n22721,n22722,n22723);
  nor U23881(n22723,n22724,n22725,n22726,n22727);
  nor U23882(n22727,n20458,n21714);
  and U23883(n22726,n20214,n21715);
  xor U23884(n20214,n22698,n22728);
  and U23885(n22728,n22697,n22695);
  nand U23886(n22695,n22729,n22730);
  or U23887(n22697,n22729,n22730);
  nand U23888(n22730,n22731,n22732,n22733,n22734);
  nand U23889(n22734,n20215,n21773);
  nand U23890(n22733,n19756,n21774);
  nand U23891(n22732,n22105,G36074);
  xor U23892(n22729,n21728,n22735);
  and U23893(n22735,n22736,n22737,n22738);
  nand U23894(n22738,n21773,n19756);
  nand U23895(n22737,n20215,n21779);
  nand U23896(n22736,n21348,n22110);
  nand U23897(n22698,n22739,n22740);
  nand U23898(n22740,n22741,n22742);
  nor U23899(n22725,n20795,n21784);
  xor U23900(n20795,n22713,n22743);
  nor U23901(n22743,n22744,n22745);
  nor U23902(n22745,n22746,n22714);
  nor U23903(n22746,n22431,n20458);
  not U23904(n20458,n20215);
  not U23905(n22744,n22710);
  nand U23906(n22714,n21787,n19756);
  nand U23907(n20215,n22747,n22748,n22749);
  nand U23908(n22749,n21691,n21348);
  nand U23909(n21348,n22750,n22751);
  nand U23910(n22751,G35978,n22209);
  nand U23911(n22750,n22752,n22753,G36004);
  nand U23912(n22748,n21669,n19105);
  nand U23913(n22747,n21670,G36403);
  nand U23914(n22713,n22754,n22755);
  nand U23915(n22755,n22756,n22757);
  or U23916(n22756,n20227,n22758);
  nor U23917(n22724,n20189,n21796);
  not U23918(n20189,n19753);
  nand U23919(n19753,n22759,n22760,n22761,n22762);
  nand U23920(n22762,n22719,n21801);
  not U23921(n22719,n20575);
  nand U23922(n20575,n22675,n22763);
  nand U23923(n22763,n22764,n21355);
  not U23924(n22675,n22628);
  nor U23925(n22628,n21355,n22764);
  nand U23926(n22764,G36200,n22765);
  not U23927(n22765,n22766);
  not U23928(n21355,G36188);
  nand U23929(n22761,G36107,n21697);
  nand U23930(n22760,G36075,n21698);
  nand U23931(n22759,G36043,n21696);
  nand U23932(n22722,G36106,n19783);
  nand U23933(n22721,n21737,n22767);
  nand U23934(n22720,n19782,n19759);
  nand U23935(G1472,n22768,n22769,n22770,n22771);
  nor U23936(n22771,n22772,n22773,n22774,n22775);
  and U23937(n22775,n20226,n21715);
  xor U23938(n20226,n22742,n22776);
  and U23939(n22776,n22741,n22739);
  nand U23940(n22739,n22777,n22778);
  or U23941(n22741,n22777,n22778);
  nand U23942(n22778,n22779,n22780,n22781,n22782);
  nand U23943(n22782,n20227,n21773);
  nand U23944(n22781,n19759,n21774);
  nand U23945(n22780,n22105,G36073);
  xor U23946(n22777,n21728,n22783);
  and U23947(n22783,n22784,n22785,n22786);
  nand U23948(n22786,n21773,n19759);
  nand U23949(n22785,n20227,n21779);
  nand U23950(n22784,n21619,n22110);
  nand U23951(n22742,n22787,n22788);
  nand U23952(n22788,n22789,n22790);
  nor U23953(n22774,n20799,n21784);
  xor U23954(n20799,n22757,n22791);
  nor U23955(n22791,n22792,n22793);
  nor U23956(n22793,n22794,n22758);
  nor U23957(n22794,n22431,n20487);
  not U23958(n20487,n20227);
  not U23959(n22792,n22754);
  nand U23960(n22758,n21787,n19759);
  nand U23961(n22757,n22795,n22796);
  nand U23962(n22796,n22797,n22798);
  or U23963(n22797,n20239,n22799);
  nor U23964(n22773,n20201,n21796);
  not U23965(n20201,n19756);
  nand U23966(n19756,n22800,n22801,n22802,n22803);
  nand U23967(n22803,n22767,n21801);
  not U23968(n22767,n20457);
  xor U23969(n20457,n22766,G36200);
  nand U23970(n22802,G36106,n21697);
  nand U23971(n22801,G36074,n21698);
  nand U23972(n22800,G36042,n21696);
  nor U23973(n22772,n20488,n19781);
  nand U23974(n22770,G36105,n19783);
  nand U23975(n22769,n19794,n20227);
  nand U23976(n20227,n22804,n22805,n22806);
  nand U23977(n22806,n21619,n21691);
  not U23978(n21619,n21336);
  nand U23979(n21336,n22807,n22808,n22809);
  nand U23980(n22808,n22810,n22209);
  nand U23981(n22807,G35977,n22811,G36004);
  nand U23982(n22805,n21669,n19167);
  nand U23983(n22804,n21670,G36402);
  not U23984(n19794,n21714);
  nand U23985(n22768,n19782,n19762);
  nand U23986(G1471,n22812,n22813,n22814,n22815);
  nor U23987(n22815,n22816,n22817,n22818,n22819);
  nor U23988(n22819,n20367,n21714);
  nor U23989(n22818,n20364,n22820);
  not U23990(n20364,n20238);
  xor U23991(n20238,n22789,n22821);
  and U23992(n22821,n22787,n22790);
  or U23993(n22790,n22822,n22823);
  nand U23994(n22787,n22822,n22823);
  nand U23995(n22823,n22824,n22825,n22826,n22827);
  nand U23996(n22827,n20239,n21773);
  nand U23997(n22826,n19762,n21774);
  nand U23998(n22825,n22105,G36072);
  xor U23999(n22822,n21728,n22828);
  and U24000(n22828,n22829,n22830,n22831);
  nand U24001(n22831,n21773,n19762);
  nand U24002(n22830,n20239,n21779);
  nand U24003(n22829,n21322,n22110);
  nand U24004(n22789,n22832,n22833);
  nand U24005(n22833,n22834,n22835);
  nor U24006(n22817,n20362,n21784);
  xor U24007(n20362,n22798,n22836);
  nor U24008(n22836,n22837,n22838);
  nor U24009(n22838,n22839,n22799);
  nor U24010(n22839,n22431,n20367);
  not U24011(n20367,n20239);
  not U24012(n22837,n22795);
  nand U24013(n22799,n21787,n19762);
  nand U24014(n20239,n22840,n22841,n22842);
  nand U24015(n22842,n21322,n21691);
  not U24016(n21322,n21603);
  nand U24017(n21603,n22843,n22844,n22811);
  nand U24018(n22844,n22845,n22209);
  nand U24019(n22843,G35976,n22846,G36004);
  nand U24020(n22841,n21669,n19212);
  nand U24021(n22840,n21670,G36401);
  nand U24022(n22798,n22847,n22848);
  nand U24023(n22848,n22849,n22850);
  or U24024(n22849,n20251,n22851);
  nor U24025(n22816,n20213,n21796);
  not U24026(n20213,n19759);
  nand U24027(n19759,n22852,n22853,n22854,n22855);
  nand U24028(n22855,n22856,n21801);
  not U24029(n22856,n20488);
  nand U24030(n20488,n22857,n22766);
  nand U24031(n22766,G36209,G36197);
  or U24032(n22857,G36209,G36197);
  nand U24033(n22854,G36105,n21697);
  nand U24034(n22853,G36073,n21698);
  nand U24035(n22852,G36041,n21696);
  nand U24036(n22814,G36104,n19783);
  nand U24037(n22813,n19782,n19765);
  nand U24038(n22812,n21737,n21316);
  nand U24039(G1470,n22858,n22859,n22860,n22861);
  nor U24040(n22861,n22862,n22863,n22864,n22865);
  nor U24041(n22865,n20555,n21714);
  and U24042(n22864,n20250,n21715);
  xor U24043(n20250,n22834,n22866);
  and U24044(n22866,n22832,n22835);
  or U24045(n22835,n22867,n22868);
  nand U24046(n22832,n22867,n22868);
  nand U24047(n22868,n22869,n22870,n22871,n22872);
  nand U24048(n22872,n19765,n21774);
  nand U24049(n22871,n20251,n21773);
  nand U24050(n22870,n22105,G36071);
  xor U24051(n22867,n21728,n22873);
  and U24052(n22873,n22874,n22875,n22876);
  nand U24053(n22876,n21308,n22110);
  nand U24054(n22875,n21773,n19765);
  nand U24055(n22874,n20251,n21779);
  nand U24056(n22834,n21294,n22877);
  nand U24057(n22877,n21295,n21292);
  nand U24058(n21292,n22878,n22879);
  nand U24059(n22879,n22880,n21776);
  or U24060(n21295,n22881,n22882);
  nand U24061(n21294,n22881,n22882);
  nand U24062(n22882,n22883,n22884,n22885,n22886);
  nand U24063(n22886,n19795,n21773);
  nand U24064(n22885,n19768,n21774);
  nand U24065(n22884,n22105,G36070);
  xor U24066(n22881,n22887,n21776);
  nand U24067(n22887,n22888,n22889,n22890);
  nand U24068(n22890,n21773,n19768);
  nand U24069(n22889,n19795,n21779);
  nand U24070(n22888,n21287,n22110);
  not U24071(n21287,n21610);
  nor U24072(n22863,n20806,n21784);
  xor U24073(n20806,n22850,n22891);
  nor U24074(n22891,n22892,n22893);
  nor U24075(n22893,n22894,n22851);
  nor U24076(n22894,n22431,n20555);
  not U24077(n20555,n20251);
  not U24078(n22892,n22847);
  nand U24079(n22851,n21787,n19765);
  nand U24080(n19765,n22895,n22896,n22897,n22898);
  nand U24081(n22898,G36103,n21697);
  nand U24082(n22897,G36071,n21698);
  nand U24083(n22896,G36039,n21696);
  nand U24084(n22895,G36190,n21801);
  nand U24085(n20251,n22899,n22900,n22901);
  nand U24086(n22901,n21308,n21691);
  not U24087(n21308,n21310);
  nand U24088(n21310,n22902,n22903);
  or U24089(n22903,G35975,G36004);
  nand U24090(n22902,G36004,n22904);
  nand U24091(n22900,n21669,n19262);
  nand U24092(n22899,n21670,G36400);
  nand U24093(n22850,n20817,n22905);
  nand U24094(n22905,n20815,n20816);
  nand U24095(n20816,n22906,n20406);
  not U24096(n22906,n22907);
  nand U24097(n20817,n22907,n21788,n19795);
  not U24098(n19795,n20406);
  nand U24099(n20406,n22908,n22909,n22910);
  nand U24100(n22910,n21691,n21610);
  nand U24101(n21610,n22911,n22912,n22913);
  nand U24102(n22912,n22914,n22209);
  nand U24103(n22911,G35974,G35973,G36004);
  nand U24104(n22909,n22915,n21669);
  nand U24105(n22908,n21670,n16048);
  nand U24106(n22907,n21787,n19768);
  nor U24107(n22862,n20225,n21796);
  not U24108(n20225,n19762);
  nand U24109(n19762,n22916,n22917,n22918,n22919);
  nand U24110(n22919,G36104,n21697);
  nand U24111(n22918,G36072,n21698);
  nand U24112(n22917,G36040,n21696);
  nand U24113(n22916,n21801,n21316);
  not U24114(n21316,G36209);
  nand U24115(n22860,G36103,n19783);
  nand U24116(n22859,n19782,n19768);
  nor U24117(n19782,n19934,n19783);
  nand U24118(n19934,n20596,n21692);
  not U24119(n20596,n20598);
  nand U24120(n22858,n21737,G36190);
  not U24121(n21737,n19781);
  nand U24122(G1469,n22920,n22921,n22922,n22923);
  nor U24123(n22923,n22924,n22925,n22926);
  nor U24124(n22926,n20506,n19781);
  nand U24125(n19781,n22927,n19789);
  not U24126(n20506,G36195);
  nor U24127(n22925,n20505,n21714);
  nand U24128(n21714,n19789,n20608);
  nor U24129(n22924,n19789,n22928);
  nand U24130(n22922,n19792,n20271);
  nand U24131(n20271,n22929,n22930,n22931);
  nand U24132(n22931,n20819,n19771);
  and U24133(n20819,n22431,n21787);
  not U24134(n22930,n20815);
  nor U24135(n20815,n20505,n22431,n22932);
  not U24136(n22431,n21788);
  nand U24137(n21788,n21755,n21743,n21747,n21753);
  nand U24138(n21743,n20635,n22933);
  nand U24139(n21755,n20622,n20635);
  nand U24140(n22929,n20505,n22932);
  and U24141(n22932,n19771,n21787);
  nand U24142(n21753,n22934,n22933);
  nand U24143(n21747,n20622,n22934);
  or U24144(n22934,n20276,n20643);
  not U24145(n19792,n21784);
  nand U24146(n21784,n19789,n22935);
  nand U24147(n22935,n21198,n20623);
  nand U24148(n22921,n21715,n20273);
  xor U24149(n20273,n22936,n21728);
  nand U24150(n22936,n22878,n22880);
  nand U24151(n22880,n22937,n22938);
  not U24152(n22938,n22939);
  xor U24153(n22937,n21776,n22940);
  not U24154(n21776,n21728);
  nand U24155(n22878,n22941,n22939);
  nand U24156(n22939,n22942,n22943,n22944,n22945);
  nor U24157(n22945,n22946,n22947);
  nor U24158(n22947,n21260,n21277);
  nor U24159(n22946,n20505,n22948);
  not U24160(n20505,n20268);
  nand U24161(n22943,n19771,n21774);
  nand U24162(n21774,n22949,n21202);
  nand U24163(n22942,n22105,G36069);
  xor U24164(n22941,n21728,n22940);
  and U24165(n22940,n22950,n22951,n22952,n22953);
  nand U24166(n22953,n21779,n20268);
  nand U24167(n20268,n22954,n22955,n22956);
  nand U24168(n22956,G35973,n21691);
  nand U24169(n22955,n21669,n19381);
  nand U24170(n22954,n21670,G36398);
  not U24171(n21691,n21710);
  not U24172(n21779,n22949);
  nor U24173(n22949,n21726,n22957);
  and U24174(n22957,n22958,n20622);
  nand U24175(n21726,n22959,n22960);
  or U24176(n22960,n20279,n22961);
  nand U24177(n22959,n22958,n22933);
  nand U24178(n22952,G35973,n22110);
  nor U24179(n22105,n21538,n22962,n21544);
  nor U24180(n22106,n21538,n22962,n21264);
  nor U24181(n21538,n20608,n20272,n21659,n22927);
  not U24182(n22927,n20615);
  not U24183(n21659,n20623);
  nand U24184(n20623,n19903,n20635);
  nor U24185(n19903,n20286,n21251);
  not U24186(n20272,n21198);
  nand U24187(n21198,n20644,n20611);
  nand U24188(n20608,n22963,n20270);
  nand U24189(n20270,n21222,n20625);
  not U24190(n21222,n21197);
  nand U24191(n21197,n20277,n20635,n21251);
  nand U24192(n22963,n21251,n21238);
  nand U24193(n22951,n21773,n19771);
  nand U24194(n19771,n22964,n22965,n22966,n22967);
  nand U24195(n22967,G36101,n21697);
  nand U24196(n22966,G36069,n21698);
  nand U24197(n22965,G36037,n21696);
  nand U24198(n22964,G36195,n21801);
  and U24199(n21724,n20622,n22968);
  nand U24200(n22968,n22961,n22969);
  nand U24201(n22969,n22970,n22971);
  nor U24202(n20622,n22972,n22973);
  nand U24203(n21725,n22974,n22975);
  nand U24204(n22975,n22933,n22971,n22970);
  nand U24205(n22970,n20621,n21263,n22976);
  nand U24206(n22976,n20643,n21653);
  not U24207(n20643,n20284);
  nand U24208(n20284,n21251,n20625);
  not U24209(n21263,n20612);
  nand U24210(n20621,n20276,n21256);
  nor U24211(n20276,n20635,n21251);
  nand U24212(n22933,n19894,n22977,n20279);
  nand U24213(n20279,n22973,n22972);
  not U24214(n22973,n22978);
  nand U24215(n22974,n22979,n22980);
  nand U24216(n22980,n22977,n19894);
  nand U24217(n19894,n22978,n22972);
  not U24218(n22977,n22981);
  not U24219(n22979,n22961);
  nand U24220(n22961,n20641,n22971,n21653);
  or U24221(n22950,n21276,n21260);
  nand U24222(n21260,n22962,n21202);
  nand U24223(n21276,n22982,n22983);
  or U24224(n22983,n21544,G36069);
  nand U24225(n22982,n21544,n22928);
  not U24226(n22928,G36101);
  not U24227(n21544,n21264);
  nor U24228(n21728,n20629,n22958);
  nor U24229(n22958,n20629,n22962,n20620);
  not U24230(n21715,n22820);
  nand U24231(n22820,n19789,n22984);
  nand U24232(n22984,n20274,n22985);
  nand U24233(n22985,n20644,n21256);
  not U24234(n20644,n20635);
  not U24235(n20274,n19788);
  nand U24236(n19788,n20617,n20620);
  nand U24237(n20620,n21251,n21256);
  not U24238(n21251,n20641);
  and U24239(n20617,n22986,n22987);
  nand U24240(n22987,n20612,n20277);
  nor U24241(n20612,n20283,n20625);
  nand U24242(n22986,n21653,n20625);
  not U24243(n21653,n21237);
  nand U24244(n21237,n20611,n20635);
  nand U24245(n22920,n19791,n19768);
  nand U24246(n19768,n22988,n22989,n22990,n22991);
  nand U24247(n22991,G36102,n21697);
  nand U24248(n22993,G36003,n22994,n22209);
  nand U24249(n22992,n22995,n22996,G36004);
  nand U24250(n22990,G36070,n21698);
  nand U24251(n22998,G36002,n22999,n22209);
  nand U24252(n22997,n23000,n23001,G36004);
  nand U24253(n22989,G36038,n21696);
  nand U24254(n23003,n22994,n22999,n22209);
  not U24255(n22994,G36002);
  nand U24256(n23002,n23001,n22996,G36004);
  not U24257(n22996,n23000);
  not U24258(n23001,n22995);
  nand U24259(n22988,G36205,n21801);
  nand U24260(n21801,n23004,n23005);
  nand U24261(n23005,G36003,G36002,n22209);
  nand U24262(n23004,n23000,n22995,G36004);
  not U24263(n19791,n21796);
  nand U24264(n21796,n20278,n19789);
  not U24265(n19789,n19783);
  nand U24266(n23006,n20615,n23007);
  nand U24267(n23007,n20605,n20281,n22981);
  nor U24268(n22981,n22972,n22978);
  nand U24269(n22978,n23008,n23009);
  nand U24270(n23009,G36005,n23010);
  nand U24271(n23008,n20295,n23011);
  nand U24272(n20295,n23012,n23013);
  nand U24273(n22972,n20292,n23014);
  or U24274(n23014,n23011,G36006);
  nand U24275(n20292,n23013,n23015);
  nand U24276(n20281,n23010,n23016);
  nand U24277(n23016,n23017,n23018,n23019,n23020);
  nor U24278(n23020,n23021,n23022,n23023,n23024);
  nand U24279(n23024,n23025,n23026,n23027);
  nand U24280(n23023,n23028,n23029,n23030,n23031);
  nand U24281(n23022,n23032,n23033,n23034,n23035);
  nand U24282(n23021,n23036,n23037,n23038,n23039);
  nor U24283(n23019,n23040,G36007,G36009,G36008);
  nand U24284(n23040,n23041,n23042,n23043,n23044);
  nor U24285(n23018,G36021,G36020,G36019,G36018);
  nor U24286(n23017,G36017,G36016,G36015,G36014);
  nand U24287(n20605,n21692,n20283);
  nand U24288(n20283,n20641,n20635);
  nand U24289(n20615,n21238,n20641);
  nand U24290(n20641,n23045,n23046,n23047);
  nand U24291(n23046,n23048,n22209);
  nand U24292(n23045,G35993,n23049,G36004);
  nor U24293(n21238,n20635,n20286);
  nand U24294(n20286,n20277,n20625);
  nand U24295(n20635,n23050,n23051,n23049);
  nand U24296(n23051,n23052,n22209);
  nand U24297(n23050,G35992,n22166,G36004);
  not U24298(n20278,n19936);
  nand U24299(n19936,n21692,n20598);
  not U24300(n21692,n20287);
  nor U24301(G1468,n20291,n23039);
  not U24302(n23039,G36036);
  nor U24303(G1467,n20291,n23038);
  not U24304(n23038,G36035);
  nor U24305(G1466,n20291,n23037);
  not U24306(n23037,G36034);
  nor U24307(G1465,n20291,n23036);
  not U24308(n23036,G36033);
  nor U24309(G1464,n20291,n23035);
  not U24310(n23035,G36032);
  nor U24311(G1463,n20291,n23034);
  not U24312(n23034,G36031);
  nor U24313(G1462,n20291,n23033);
  not U24314(n23033,G36030);
  nor U24315(G1461,n20291,n23032);
  not U24316(n23032,G36029);
  nor U24317(G1460,n20291,n23031);
  not U24318(n23031,G36028);
  nor U24319(G1459,n20291,n23030);
  not U24320(n23030,G36027);
  nor U24321(G1458,n20291,n23029);
  not U24322(n23029,G36026);
  nor U24323(G1457,n20291,n23028);
  not U24324(n23028,G36025);
  nor U24325(G1456,n20291,n23026);
  not U24326(n23026,G36024);
  nor U24327(G1455,n20291,n23025);
  not U24328(n23025,G36023);
  nor U24329(G1454,n20291,n23027);
  not U24330(n23027,G36022);
  and U24331(G1453,n20290,G36021);
  and U24332(G1452,n20290,G36020);
  and U24333(G1451,n20290,G36019);
  and U24334(G1450,n20290,G36018);
  and U24335(G1449,n20290,G36017);
  and U24336(G1448,n20290,G36016);
  and U24337(G1447,n20290,G36015);
  and U24338(G1446,n20290,G36014);
  nor U24339(G1445,n20291,n23044);
  not U24340(n23044,G36013);
  nor U24341(G1444,n20291,n23043);
  not U24342(n23043,G36012);
  nor U24343(G1443,n20291,n23042);
  not U24344(n23042,G36011);
  nor U24345(G1442,n20291,n23041);
  not U24346(n23041,G36010);
  not U24347(n20291,n20290);
  and U24348(G1441,n20290,G36009);
  and U24349(G1440,n20290,G36008);
  and U24350(G1439,n20290,G36007);
  nand U24351(n20290,n20282,n23011);
  not U24352(n23011,n23010);
  nor U24353(n23010,n23013,n23053);
  and U24354(n23053,n23054,n23015);
  xnor U24355(n23054,n23012,G36185);
  nor U24356(n20282,n22962,G1406,n20629);
  not U24357(n20629,n21202);
  nand U24358(G1438,n23055,n23056,n23057);
  nand U24359(n23057,n23058,G36429);
  nand U24360(n23056,n23059,n22999,n23060);
  nand U24361(n23055,n23061,n17853);
  and U24362(n17853,n23062,n23063);
  nand U24363(n23063,n23064,n23065,n23066);
  not U24364(n23066,n23067);
  nand U24365(n23065,n23068,n23069);
  nand U24366(n23062,n23068,n23070,n23067);
  xor U24367(n23067,n23071,G1);
  nand U24368(n23071,n23072,n23073);
  nand U24369(n23073,n15634,n15644);
  not U24370(n15644,G36429);
  or U24371(n23072,n15634,G36184);
  nand U24372(n23070,G2,n23064);
  nand U24373(n23064,n23074,n23075);
  nand U24374(n23068,n23076,n23077);
  nand U24375(G1437,n23078,n23079,n23080,n23081);
  nand U24376(n23081,n23061,n17869);
  xor U24377(n17869,n23082,n23076);
  not U24378(n23076,n23075);
  nand U24379(n23075,n23083,n23084);
  nand U24380(n23084,n15634,n15645);
  not U24381(n15645,G36428);
  nand U24382(n23083,n15649,n15647);
  not U24383(n15647,G36183);
  xor U24384(n23082,n23069,n23074);
  not U24385(n23074,n23077);
  nand U24386(n23077,n23085,n23086);
  nand U24387(n23086,G3,n23087);
  nand U24388(n23087,n23088,n23089);
  or U24389(n23085,n23089,n23088);
  not U24390(n23069,G2);
  nand U24391(n23080,n23060,n22995);
  xor U24392(n22995,n22999,n23059);
  not U24393(n22999,G36003);
  nand U24394(n23079,n23058,G36428);
  nand U24395(n23078,n23090,G36003);
  nand U24396(G1436,n23091,n23092,n23093,n23094);
  nand U24397(n23094,n23061,n17943);
  xnor U24398(n17943,n23095,n23089);
  nand U24399(n23089,n23096,n23097);
  or U24400(n23097,n15649,G36427);
  nand U24401(n23096,n15649,n15661);
  not U24402(n15661,G36182);
  xnor U24403(n23095,G3,n23088);
  and U24404(n23088,n23098,n23099);
  nand U24405(n23099,G4,n23100);
  nand U24406(n23100,n23101,n23102);
  or U24407(n23098,n23102,n23101);
  nand U24408(n23093,n23060,n23000);
  nor U24409(n23000,n23059,n23103);
  and U24410(n23103,G36002,n23104);
  nor U24411(n23059,n23104,G36002);
  nand U24412(n23092,n23058,G36427);
  nand U24413(n23091,n23090,G36002);
  nand U24414(G1435,n23105,n23106,n23107,n23108);
  nand U24415(n23108,G36001,n23109);
  nand U24416(n23109,n23110,n23111);
  nand U24417(n23111,n23060,n23112);
  nand U24418(n23107,n23060,n23113,n23114);
  nand U24419(n23106,n23061,n17982);
  xnor U24420(n17982,n23115,n23102);
  nand U24421(n23102,n23116,n23117);
  or U24422(n23117,n15649,G36426);
  nand U24423(n23116,n15649,n15676);
  not U24424(n15676,G36181);
  xnor U24425(n23115,G4,n23101);
  nor U24426(n23101,n23118,n23119);
  not U24427(n23119,n23120);
  nand U24428(n23105,n23058,G36426);
  nand U24429(G1434,n23121,n23122,n23123,n23124);
  nand U24430(n23124,n23125,n23113,n23060);
  nand U24431(n23123,n23061,n18022);
  and U24432(n18022,n23126,n23127);
  nand U24433(n23127,n23118,n23120);
  nor U24434(n23118,n23128,n23129);
  not U24435(n23129,n23130);
  nand U24436(n23126,n23128,n23131);
  nand U24437(n23131,n23130,n23120);
  nand U24438(n23120,n23132,n23133,G5);
  or U24439(n23133,n15649,G36425);
  nand U24440(n23132,n15649,n15688);
  not U24441(n15688,G36180);
  nand U24442(n23130,n23134,n23135,n23136);
  not U24443(n23136,G5);
  nand U24444(n23135,n15649,G36180);
  nand U24445(n23134,n15634,G36425);
  nand U24446(n23128,n23137,n23138);
  nand U24447(n23138,n23139,n23140);
  not U24448(n23140,G6);
  or U24449(n23139,n23141,n23142);
  nand U24450(n23137,n23142,n23141);
  nand U24451(n23122,n23058,G36425);
  nand U24452(n23121,n23090,G36000);
  nand U24453(G1433,n23143,n23144,n23145,n23146);
  nand U24454(n23146,n23147,n23148,n23060);
  nand U24455(n23145,n23061,n18063);
  xor U24456(n18063,n23149,n23142);
  nand U24457(n23142,n23150,n23151);
  or U24458(n23151,n15649,G36424);
  nand U24459(n23150,n15649,n15699);
  not U24460(n15699,G36179);
  xor U24461(n23149,n23141,G6);
  nand U24462(n23141,n23152,n23153);
  nand U24463(n23153,n23154,n23155);
  not U24464(n23155,G7);
  or U24465(n23154,n23156,n23157);
  nand U24466(n23152,n23157,n23156);
  nand U24467(n23144,n23058,G36424);
  nand U24468(n23143,n23090,G35999);
  nand U24469(G1432,n23158,n23159,n23160,n23161);
  nand U24470(n23161,G35998,n23162);
  nand U24471(n23162,n23110,n23163);
  nand U24472(n23163,n23060,n23164);
  nand U24473(n23160,n23060,n23165,n23166);
  nand U24474(n23159,n23061,n18105);
  xor U24475(n18105,n23167,n23157);
  nand U24476(n23157,n23168,n23169);
  or U24477(n23169,n15649,G36423);
  nand U24478(n23168,n15649,n15713);
  not U24479(n15713,G36178);
  xor U24480(n23167,n23156,G7);
  nand U24481(n23156,n23170,n23171);
  nand U24482(n23171,n23172,n23173);
  not U24483(n23173,G8);
  or U24484(n23172,n23174,n23175);
  nand U24485(n23170,n23175,n23174);
  nand U24486(n23158,n23058,G36423);
  nand U24487(G1431,n23176,n23177,n23178,n23179);
  nand U24488(n23179,n23180,n23165,n23060);
  nand U24489(n23178,n23061,n18143);
  xor U24490(n18143,n23181,n23175);
  nand U24491(n23175,n23182,n23183);
  or U24492(n23183,n15649,G36422);
  nand U24493(n23182,n15649,n15725);
  not U24494(n15725,G36177);
  xor U24495(n23181,n23174,G8);
  nand U24496(n23174,n23184,n23185);
  nand U24497(n23185,n23186,n23187);
  not U24498(n23187,G9);
  or U24499(n23186,n23188,n23189);
  nand U24500(n23184,n23189,n23188);
  nand U24501(n23177,n23058,G36422);
  nand U24502(n23176,n23090,G35997);
  nand U24503(G1430,n23190,n23191,n23192,n23193);
  nand U24504(n23193,G35996,n23194);
  nand U24505(n23194,n23110,n23195);
  nand U24506(n23195,n23060,n23196);
  nand U24507(n23192,n23060,n23197,n23198);
  nand U24508(n23191,n23061,n18182);
  xor U24509(n18182,n23199,n23189);
  nand U24510(n23189,n23200,n23201);
  or U24511(n23201,n15649,G36421);
  nand U24512(n23200,n15649,n15744);
  not U24513(n15744,G36176);
  xor U24514(n23199,n23188,G9);
  nand U24515(n23188,n23202,n23203);
  nand U24516(n23203,n23204,n23205);
  not U24517(n23205,G10);
  or U24518(n23204,n23206,n23207);
  nand U24519(n23202,n23207,n23206);
  nand U24520(n23190,n23058,G36421);
  nand U24521(G1429,n23208,n23209,n23210,n23211);
  nand U24522(n23211,n23212,n23197,n23060);
  nand U24523(n23210,n23061,n18224);
  xor U24524(n18224,n23213,n23207);
  nand U24525(n23207,n23214,n23215);
  or U24526(n23215,n15649,G36420);
  nand U24527(n23214,n15649,n15756);
  not U24528(n15756,G36175);
  xor U24529(n23213,n23206,G10);
  nand U24530(n23206,n23216,n23217);
  nand U24531(n23217,n23218,n23219);
  not U24532(n23219,G11);
  or U24533(n23218,n23220,n23221);
  nand U24534(n23216,n23221,n23220);
  nand U24535(n23209,n23058,G36420);
  nand U24536(n23208,n23090,G35995);
  nand U24537(G1428,n23222,n23223,n23224,n23225);
  nand U24538(n23225,n23226,n23227,n23060);
  nand U24539(n23224,n23061,n18261);
  xor U24540(n18261,n23228,n23221);
  nand U24541(n23221,n23229,n23230);
  or U24542(n23230,n15649,G36419);
  nand U24543(n23229,n15649,n15774);
  not U24544(n15774,G36174);
  xor U24545(n23228,n23220,G11);
  nand U24546(n23220,n23231,n23232);
  nand U24547(n23232,n23233,n23234);
  not U24548(n23234,G12);
  or U24549(n23233,n23235,n23236);
  nand U24550(n23231,n23236,n23235);
  nand U24551(n23223,n23058,G36419);
  nand U24552(n23222,n23090,G35994);
  nand U24553(G1427,n23237,n23238,n23239,n23240);
  nand U24554(n23240,G35993,n23241);
  nand U24555(n23241,n23110,n23242);
  nand U24556(n23242,n23060,n23243);
  nand U24557(n23239,n23060,n23049,n23048);
  nand U24558(n23238,n23061,n18301);
  xor U24559(n18301,n23244,n23236);
  nand U24560(n23236,n23245,n23246);
  or U24561(n23246,n15649,G36418);
  nand U24562(n23245,n15649,n15788);
  not U24563(n15788,G36173);
  xor U24564(n23244,n23235,G12);
  nand U24565(n23235,n23247,n23248);
  nand U24566(n23248,n23249,n23250);
  not U24567(n23250,G13);
  or U24568(n23249,n23251,n23252);
  nand U24569(n23247,n23252,n23251);
  nand U24570(n23237,n23058,G36418);
  nand U24571(G1426,n23253,n23254,n23255,n23256);
  nand U24572(n23256,G35992,n23257);
  nand U24573(n23257,n23110,n23258);
  nand U24574(n23258,n23060,n23259);
  nand U24575(n23255,n23060,n22166,n23052);
  nand U24576(n23254,n23061,n18353);
  xor U24577(n18353,n23260,n23252);
  nand U24578(n23252,n23261,n23262);
  or U24579(n23262,n15649,G36417);
  nand U24580(n23261,n15649,n15800);
  not U24581(n15800,G36172);
  xor U24582(n23260,n23251,G13);
  nand U24583(n23251,n23263,n23264);
  nand U24584(n23264,n23265,n23266);
  not U24585(n23266,G14);
  or U24586(n23265,n23267,n23268);
  nand U24587(n23263,n23268,n23267);
  nand U24588(n23253,n23058,G36417);
  nand U24589(G1425,n23269,n23270,n23271,n23272);
  nand U24590(n23272,n22167,n22166,n23060);
  not U24591(n22166,n23259);
  nand U24592(n22167,G35991,n22211);
  nand U24593(n23271,n23061,n18410);
  xor U24594(n18410,n23273,n23268);
  nand U24595(n23268,n23274,n23275);
  or U24596(n23275,n15649,G36416);
  nand U24597(n23274,n15649,n15815);
  not U24598(n15815,G36171);
  xor U24599(n23273,n23267,G14);
  nand U24600(n23267,n23276,n23277);
  nand U24601(n23277,n23278,n23279);
  not U24602(n23279,G15);
  or U24603(n23278,n23280,n23281);
  nand U24604(n23276,n23281,n23280);
  nand U24605(n23270,n23058,G36416);
  nand U24606(n23269,n23090,G35991);
  nand U24607(G1424,n23282,n23283,n23284,n23285);
  nand U24608(n23285,n22212,n22211,n23060);
  nand U24609(n22212,G35990,n23286);
  nand U24610(n23286,n23287,n22257);
  nand U24611(n23284,n23061,n18461);
  xor U24612(n18461,n23288,n23281);
  nand U24613(n23281,n23289,n23290);
  or U24614(n23290,n15649,G36415);
  nand U24615(n23289,n15649,n15832);
  not U24616(n15832,G36170);
  xor U24617(n23288,n23280,G15);
  nand U24618(n23280,n23291,n23292);
  nand U24619(n23292,n23293,n23294);
  not U24620(n23294,G16);
  nand U24621(n23293,n23295,n23296);
  or U24622(n23291,n23296,n23295);
  nand U24623(n23283,n23058,G36415);
  nand U24624(n23282,n23090,G35990);
  nand U24625(G1423,n23297,n23298,n23299,n23300);
  or U24626(n23300,n22258,n23301);
  xnor U24627(n22258,n22257,n23287);
  nand U24628(n23299,n23061,n18518);
  xor U24629(n18518,n23302,n23295);
  nand U24630(n23295,n23303,n23304);
  nand U24631(n23304,n15649,G36169);
  nand U24632(n23303,n15634,G36414);
  xor U24633(n23302,n23296,G16);
  nand U24634(n23296,n23305,n23306);
  nand U24635(n23306,G17,n23307);
  or U24636(n23307,n23308,n23309);
  nand U24637(n23305,n23309,n23308);
  nand U24638(n23298,n23058,G36414);
  nand U24639(n23297,n23090,G35989);
  nand U24640(G1422,n23310,n23311,n23312,n23313);
  or U24641(n23313,n22299,n23301);
  xnor U24642(n22299,n22345,G35988);
  nand U24643(n23312,n23061,n18568);
  xor U24644(n18568,n23314,n23309);
  nand U24645(n23309,n23315,n23316);
  nand U24646(n23316,n15649,G36168);
  nand U24647(n23315,n15634,G36413);
  xor U24648(n23314,n23308,G17);
  nand U24649(n23311,n23058,G36413);
  nand U24650(n23310,n23090,G35988);
  nand U24651(G1421,n23317,n23318,n23319,n23320);
  nand U24652(n23320,n22346,n22345,n23060);
  nand U24653(n22346,G35987,n22388);
  nand U24654(n23319,n23061,n18626);
  nand U24655(n18626,n23321,n23322);
  nand U24656(n23322,n23323,n23324);
  not U24657(n23323,n23308);
  nand U24658(n23308,n23325,n23326,n23327);
  nand U24659(n23321,n23328,n23329);
  nand U24660(n23329,n23327,n23326,n23330);
  not U24661(n23330,n23325);
  nand U24662(n23325,n23328,n23324);
  nand U24663(n23324,n23331,n23332,n23333);
  nand U24664(n23332,n15649,G36167);
  nand U24665(n23331,n15634,G36412);
  nand U24666(n23326,G36412,n15634,G18);
  nand U24667(n23327,n15879,G36167);
  nor U24668(n15879,n23333,n15634);
  not U24669(n23333,G18);
  and U24670(n23328,n23334,n23335);
  nand U24671(n23335,n23336,n23337);
  not U24672(n23337,G19);
  or U24673(n23336,n23338,n23339);
  nand U24674(n23334,n23339,n23338);
  nand U24675(n23318,n23058,G36412);
  nand U24676(n23317,n23090,G35987);
  nand U24677(G1420,n23340,n23341,n23342,n23343);
  nand U24678(n23343,n22389,n22388,n23060);
  nand U24679(n22389,G35986,n22437);
  nand U24680(n23342,n23061,n18678);
  xor U24681(n18678,n23344,n23339);
  nand U24682(n23339,n23345,n23346);
  or U24683(n23346,n15649,G36411);
  nand U24684(n23345,n15649,n15885);
  not U24685(n15885,G36166);
  xor U24686(n23344,n23338,G19);
  nand U24687(n23338,n23347,n23348);
  nand U24688(n23348,n23349,n23350);
  not U24689(n23350,G20);
  nand U24690(n23349,n23351,n23352);
  or U24691(n23347,n23352,n23351);
  nand U24692(n23341,n23058,G36411);
  nand U24693(n23340,n23090,G35986);
  nand U24694(G1419,n23353,n23354,n23355,n23356);
  nand U24695(n23356,G35985,n23357);
  nand U24696(n23357,n23110,n23358);
  nand U24697(n23358,n23060,n23359);
  nand U24698(n23355,n23060,n22439,n22438);
  nand U24699(n23354,n23061,n18738);
  xor U24700(n18738,n23360,n23351);
  nand U24701(n23351,n23361,n23362);
  nand U24702(n23362,n15649,G36165);
  nand U24703(n23361,n15634,G36410);
  xor U24704(n23360,n23352,G20);
  nand U24705(n23352,n23363,n23364);
  nand U24706(n23364,G21,n23365);
  or U24707(n23365,n23366,n23367);
  nand U24708(n23363,n23367,n23366);
  nand U24709(n23353,n23058,G36410);
  nand U24710(G1418,n23368,n23369,n23370,n23371);
  nand U24711(n23371,G35984,n23372);
  nand U24712(n23372,n23110,n23373);
  nand U24713(n23373,n23060,n23374);
  nand U24714(n23370,n23060,n22483,n22482);
  nand U24715(n23369,n23061,n18791);
  xor U24716(n18791,n23375,n23367);
  nand U24717(n23367,n23376,n23377);
  nand U24718(n23377,n15649,G36164);
  nand U24719(n23376,n15634,G36409);
  xor U24720(n23375,n23366,G21);
  nand U24721(n23368,n23058,G36409);
  nand U24722(G1417,n23378,n23379,n23380,n23381);
  or U24723(n23381,n22527,n23301);
  nand U24724(n22527,n22483,n23382);
  nand U24725(n23382,G35983,n22569);
  not U24726(n22483,n23374);
  nand U24727(n23380,n23061,n18843);
  nand U24728(n18843,n23383,n23384);
  nand U24729(n23384,n23385,n23386);
  not U24730(n23385,n23366);
  nand U24731(n23366,n23387,n23388,n23389);
  nand U24732(n23383,n23390,n23391);
  nand U24733(n23391,n23389,n23388,n23392);
  not U24734(n23392,n23387);
  nand U24735(n23387,n23390,n23386);
  nand U24736(n23386,n23393,n23394,n23395);
  nand U24737(n23394,n15649,G36163);
  nand U24738(n23393,n15634,G36408);
  nand U24739(n23388,G36408,n15634,G22);
  nand U24740(n23389,n15932,G36163);
  nor U24741(n15932,n23395,n15634);
  not U24742(n23395,G22);
  and U24743(n23390,n23396,n23397);
  nand U24744(n23397,n23398,n23399);
  not U24745(n23399,G23);
  or U24746(n23398,n23400,n23401);
  nand U24747(n23396,n23401,n23400);
  nand U24748(n23379,n23058,G36408);
  nand U24749(n23378,n23090,G35983);
  nand U24750(G1416,n23402,n23403,n23404,n23405);
  nand U24751(n23405,G35982,n23406);
  nand U24752(n23406,n23110,n23407);
  nand U24753(n23407,n23060,n23408);
  nand U24754(n23404,n23060,n22571,n22570);
  nand U24755(n23403,n23061,n18898);
  xor U24756(n18898,n23409,n23401);
  nand U24757(n23401,n23410,n23411);
  or U24758(n23411,n15649,G36407);
  nand U24759(n23410,n15649,n15938);
  not U24760(n15938,G36162);
  xor U24761(n23409,n23400,G23);
  nand U24762(n23400,n23412,n23413);
  nand U24763(n23413,n23414,n23415);
  not U24764(n23415,G24);
  or U24765(n23414,n23416,n23417);
  nand U24766(n23412,n23417,n23416);
  nand U24767(n23402,n23058,G36407);
  nand U24768(G1415,n23418,n23419,n23420,n23421);
  or U24769(n23421,n22616,n23301);
  nand U24770(n22616,n22571,n23422);
  nand U24771(n23422,G35981,n22662);
  not U24772(n22571,n23408);
  nand U24773(n23420,n23061,n18946);
  xor U24774(n18946,n23423,n23417);
  nand U24775(n23417,n23424,n23425);
  or U24776(n23425,n15649,G36406);
  nand U24777(n23424,n15649,n15950);
  not U24778(n15950,G36161);
  xor U24779(n23423,n23416,G24);
  nand U24780(n23416,n23426,n23427);
  nand U24781(n23427,n23428,n23429);
  or U24782(n23428,n23430,n23431);
  nand U24783(n23426,n23431,n23430);
  nand U24784(n23419,n23058,G36406);
  nand U24785(n23418,n23090,G35981);
  nand U24786(G1414,n23432,n23433,n23434,n23435);
  nand U24787(n23435,G35980,n23436);
  nand U24788(n23436,n23110,n23437);
  nand U24789(n23437,n23060,n23438);
  nand U24790(n23434,n23060,n22664,n22663);
  nand U24791(n23433,n23061,n19002);
  xnor U24792(n19002,n23439,n23430);
  and U24793(n23430,n23440,n23441);
  nand U24794(n23441,n15649,G36160);
  nand U24795(n23440,n15634,G36405);
  xor U24796(n23439,n23431,n23429);
  not U24797(n23429,G25);
  nor U24798(n23431,n23442,n23443);
  and U24799(n23443,n23444,n23445);
  nand U24800(n23432,n23058,G36405);
  nand U24801(G1413,n23446,n23447,n23448,n23449);
  nand U24802(n23449,n22709,n22664,n23060);
  not U24803(n22664,n23438);
  nand U24804(n22709,G35979,n22753);
  nand U24805(n23448,n23061,n19053);
  xor U24806(n19053,n23445,n23450);
  nor U24807(n23450,n23451,n23442);
  nand U24808(n23442,n23452,n23453);
  nand U24809(n23453,G36404,n15634,G26);
  nand U24810(n23452,n15986,G36159);
  nor U24811(n15986,n23454,n15634);
  not U24812(n23451,n23444);
  nand U24813(n23444,n23455,n23456,n23454);
  not U24814(n23454,G26);
  nand U24815(n23456,n15649,G36159);
  nand U24816(n23455,n15634,G36404);
  nand U24817(n23445,n23457,n23458);
  nand U24818(n23458,n23459,n23460);
  nand U24819(n23447,n23058,G36404);
  nand U24820(n23446,n23090,G35979);
  nand U24821(G1412,n23461,n23462,n23463,n23464);
  nand U24822(n23464,n22752,n22753,n23060);
  nand U24823(n22752,G35978,n22809);
  nand U24824(n23463,n23061,n19105);
  xor U24825(n19105,n23460,n23465);
  and U24826(n23465,n23459,n23457);
  and U24827(n23457,n23466,n23467);
  nand U24828(n23467,G36403,n15634,G27);
  nand U24829(n23466,n15997,G36158);
  nor U24830(n15997,n23468,n15634);
  nand U24831(n23459,n23469,n23470,n23468);
  not U24832(n23468,G27);
  nand U24833(n23470,n15649,G36158);
  nand U24834(n23469,n15634,G36403);
  nand U24835(n23460,n23471,n23472);
  or U24836(n23472,n23473,n23474);
  not U24837(n23471,n23475);
  nand U24838(n23462,n23058,G36403);
  nand U24839(n23461,n23090,G35978);
  nand U24840(G1411,n23476,n23477,n23478,n23479);
  nand U24841(n23479,G35977,n23480);
  nand U24842(n23480,n23110,n23481);
  nand U24843(n23481,n23060,n23482);
  nand U24844(n23478,n23060,n22811,n22810);
  nand U24845(n23477,n23061,n19167);
  xnor U24846(n19167,n23473,n23483);
  nor U24847(n23483,n23474,n23475);
  nand U24848(n23475,n23484,n23485);
  nand U24849(n23485,G36402,n15634,G28);
  nand U24850(n23484,n16012,G36157);
  nor U24851(n16012,n23486,n15634);
  and U24852(n23474,n23487,n23488,n23486);
  not U24853(n23486,G28);
  nand U24854(n23488,n15649,G36157);
  nand U24855(n23487,n15634,G36402);
  nand U24856(n23473,n23489,n23490);
  nand U24857(n23490,n23491,n23492);
  not U24858(n23492,G29);
  or U24859(n23491,n23493,n23494);
  nand U24860(n23489,n23494,n23493);
  nand U24861(n23476,n23058,G36402);
  nand U24862(G1410,n23495,n23496,n23497,n23498);
  nand U24863(n23498,G35976,n23499);
  nand U24864(n23499,n23110,n23500);
  nand U24865(n23500,n23060,n23501);
  nand U24866(n23497,n23060,n22846,n22845);
  nand U24867(n23496,n23061,n19212);
  xor U24868(n19212,n23502,n23494);
  nand U24869(n23494,n23503,n23504);
  or U24870(n23504,n15649,G36401);
  nand U24871(n23503,n15649,n16018);
  not U24872(n16018,G36156);
  xor U24873(n23502,n23493,G29);
  nand U24874(n23493,n23505,n23506);
  nand U24875(n23506,n23507,n23508);
  not U24876(n23508,G30);
  nand U24877(n23507,n23509,n23510);
  or U24878(n23505,n23510,n23509);
  nand U24879(n23495,n23058,G36401);
  nand U24880(G1409,n23511,n23512,n23513,n23514);
  or U24881(n23514,n22904,n23301);
  nand U24882(n22904,n22846,n23515);
  nand U24883(n23515,G35975,n22913);
  not U24884(n22846,n23501);
  nand U24885(n23513,n23061,n19262);
  xor U24886(n19262,n23516,n23509);
  nand U24887(n23509,n23517,n23518);
  nand U24888(n23518,n15649,G36155);
  nand U24889(n23517,n15634,G36400);
  xor U24890(n23516,n23510,G30);
  nand U24891(n23510,n23519,n23520);
  nand U24892(n23520,G31,n23521);
  nand U24893(n23512,n23058,G36400);
  nand U24894(n23511,n23090,G35975);
  not U24895(n23090,n23110);
  nand U24896(G1408,n23522,n23523,n23524,n23525);
  nand U24897(n23525,G35974,n23526);
  nand U24898(n23526,n23110,n23527);
  nand U24899(n23527,n23060,n21277);
  nand U24900(n23524,n23060,G35973,n22914);
  nand U24901(n23523,n23061,n19320);
  not U24902(n19320,n22915);
  xor U24903(n22915,n23528,G31);
  nand U24904(n23528,n23521,n23519);
  nand U24905(n23519,n23529,n23530,n23531);
  nand U24906(n23530,n15634,n16048);
  not U24907(n16048,G36399);
  nand U24908(n23529,n15649,n16050);
  not U24909(n16050,G36154);
  nand U24910(n23521,n23532,n23533,n23534);
  nand U24911(n23533,n15649,G36154);
  nand U24912(n23532,n15634,G36399);
  nand U24913(n23522,n23058,G36399);
  nand U24914(G1407,n23535,n23536,n23537);
  nand U24915(n23537,n23061,n19381);
  and U24916(n19381,n23534,n23538);
  nand U24917(n23538,n23539,n23540);
  not U24918(n23534,n23531);
  nor U24919(n23531,n23539,n23540);
  not U24920(n23540,G32);
  nand U24921(n23539,n23541,n23542);
  nand U24922(n23542,n15634,n16066);
  not U24923(n16066,G36398);
  or U24924(n23541,n15634,G36153);
  nand U24925(n23536,G35973,n23543);
  nand U24926(n23543,n23110,n23301);
  nand U24927(n23301,n23110,G36215);
  nand U24928(n23110,G36215,n22209);
  nand U24929(n23535,n23058,G36398);
  or U24930(n23545,n21535,G36461,n17712,G36623);
  not U24931(n17712,G36378);
  or U24932(n23544,G36216,G36378,G36133,n14016);
  not U24933(G1406,G36215);
  nand U24934(G1341,n23546,G36215);
  nand U24935(n23546,n23547,n21710);
  nand U24936(n21710,n21264,n20598);
  nand U24937(n20598,n23548,n23549,n23104);
  nand U24938(n23104,n23112,n23114);
  nand U24939(n23549,n23114,n22209);
  not U24940(n23114,G36001);
  nand U24941(n23548,G36001,n23113,G36004);
  nand U24942(n21264,n23550,n23551);
  or U24943(n23551,G36000,G36004);
  nand U24944(n23550,G36004,n23552);
  nand U24945(n23552,n23113,n23125);
  nand U24946(n23125,G36000,n23148);
  not U24947(n23113,n23112);
  nor U24948(n23112,n23148,G36000);
  nand U24949(n23547,n21202,n23553);
  nand U24950(n23553,n20287,n22971);
  not U24951(n22971,n22962);
  nor U24952(n22962,n23013,n23012,n23015);
  nand U24953(n23015,n23554,n23555,n23556);
  nand U24954(n23555,n23166,n22209);
  nand U24955(n23554,G35998,n23165,G36004);
  and U24956(n23012,n23557,n23558);
  nand U24957(n23558,G35997,n22209);
  nand U24958(n23557,n23180,n23165,G36004);
  not U24959(n23165,n23164);
  nand U24960(n23180,G35997,n23559);
  nand U24961(n23559,n23196,n23198);
  nand U24962(n23013,n23560,n23561);
  or U24963(n23561,G35999,G36004);
  nand U24964(n23560,G36004,n23562);
  nand U24965(n23562,n23148,n23147);
  nand U24966(n23147,G35999,n23556);
  or U24967(n23148,n23556,G35999);
  nand U24968(n23556,n23164,n23166);
  not U24969(n23166,G35998);
  nor U24970(n23164,G35996,G35997,n23197);
  nand U24971(n20287,n21256,n20611);
  not U24972(n20611,n20277);
  nand U24973(n20277,n23563,n23564);
  or U24974(n23564,G35995,G36004);
  nand U24975(n23563,G36004,n23565);
  nand U24976(n23565,n23197,n23212);
  nand U24977(n23212,G35995,n23227);
  not U24978(n23197,n23196);
  not U24979(n21256,n20625);
  nand U24980(n20625,n23566,n23567);
  or U24981(n23567,G35994,G36004);
  nand U24982(n23566,G36004,n23568);
  nand U24983(n23568,n23227,n23226);
  nand U24984(n23226,G35994,n23047);
  xor U24985(n21202,n23198,n23569);
  nor U24986(n23569,n23196,n22209);
  not U24987(n22209,G36004);
  nor U24988(n23196,n23227,G35995);
  or U24989(n23227,n23047,G35994);
  nand U24990(n23047,n23243,n23048);
  not U24991(n23048,G35993);
  not U24992(n23243,n23049);
  nand U24993(n23049,n23259,n23052);
  not U24994(n23052,G35992);
  nor U24995(n23259,n22211,G35991);
  nand U24996(n22211,n22257,n22208,n23287);
  nor U24997(n23287,n22345,G35988);
  or U24998(n22345,n22388,G35987);
  or U24999(n22388,n22437,G35986);
  nand U25000(n22437,n23359,n22438);
  not U25001(n22438,G35985);
  not U25002(n23359,n22439);
  nand U25003(n22439,n23374,n22482);
  not U25004(n22482,G35984);
  nor U25005(n23374,n22569,G35983);
  nand U25006(n22569,n23408,n22570);
  not U25007(n22570,G35982);
  nor U25008(n23408,n22662,G35981);
  nand U25009(n22662,n23438,n22663);
  not U25010(n22663,G35980);
  nor U25011(n23438,n22753,G35979);
  or U25012(n22753,n22809,G35978);
  nand U25013(n22809,n23482,n22810);
  not U25014(n22810,G35977);
  not U25015(n23482,n22811);
  nand U25016(n22811,n23501,n22845);
  not U25017(n22845,G35976);
  nor U25018(n23501,n22913,G35975);
  nand U25019(n22913,n21277,n22914);
  not U25020(n22914,G35974);
  not U25021(n21277,G35973);
  not U25022(n22208,G35990);
  not U25023(n22257,G35989);
  not U25024(n23198,G35996);
  nand U25025(G10242,n23570,n23571);
  nand U25026(n23571,n23572,n23573);
  nand U25027(n23573,n23574,n23575);
  not U25028(n23572,n23576);
  nand U25029(n23570,n23574,n23575,n23576);
  nand U25030(G10240,n23577,n23578);
  nand U25031(n23578,n23579,n23580);
  nand U25032(n23580,n23581,n23582);
  not U25033(n23579,n23583);
  nand U25034(n23577,n23581,n23582,n23583);
  nand U25035(G10238,n23584,n23585);
  nand U25036(n23585,n23586,n23587);
  nand U25037(n23587,n23588,n23589);
  not U25038(n23586,n23590);
  nand U25039(n23584,n23588,n23589,n23590);
  nand U25040(G10236,n23591,n23592);
  nand U25041(n23592,n23593,n23594);
  nand U25042(n23594,n23595,n23596);
  not U25043(n23593,n23597);
  nand U25044(n23591,n23595,n23596,n23597);
  nand U25045(G10234,n23598,n23599);
  nand U25046(n23599,n23600,n23601);
  nand U25047(n23601,n23602,n23603);
  not U25048(n23600,n23604);
  nand U25049(n23598,n23602,n23603,n23604);
  nand U25050(G10232,n23605,n23606);
  nand U25051(n23606,n23607,n23608);
  nand U25052(n23608,n23609,n23610);
  not U25053(n23607,n23611);
  nand U25054(n23605,n23609,n23610,n23611);
  nand U25055(G10230,n23612,n23613);
  nand U25056(n23613,n23614,n23615);
  nand U25057(n23615,n23616,n23617);
  not U25058(n23614,n23618);
  nand U25059(n23612,n23616,n23617,n23618);
  nand U25060(G10228,n23619,n23620);
  nand U25061(n23620,n23621,n23622);
  nand U25062(n23622,n23623,n23624);
  not U25063(n23621,n23625);
  nand U25064(n23619,n23623,n23624,n23625);
  nand U25065(G10226,n23626,n23627);
  nand U25066(n23627,n23628,n23629);
  nand U25067(n23629,n23630,n23631);
  nand U25068(n23626,n23630,n23631,n23632);
  nand U25069(G10222,n23633,n23634);
  nand U25070(n23634,n23635,n23636);
  nand U25071(n23635,n23637,n23638);
  nand U25072(n23633,n23637,n23638,n23639);
  nand U25073(G10220,n23640,n23641);
  nand U25074(n23641,n23642,n23643);
  nand U25075(n23643,n23644,n23645);
  not U25076(n23642,n23646);
  nand U25077(n23640,n23644,n23645,n23646);
  nand U25078(G10218,n23647,n23648);
  nand U25079(n23648,n23649,n23650);
  nand U25080(n23650,n23651,n23652);
  not U25081(n23649,n23653);
  nand U25082(n23647,n23651,n23652,n23653);
  nand U25083(G10216,n23654,n23655);
  nand U25084(n23655,n23656,n23657);
  nand U25085(n23657,n23658,n23659);
  not U25086(n23656,n23660);
  nand U25087(n23654,n23658,n23659,n23660);
  nand U25088(G10214,n23661,n23662);
  nand U25089(n23662,n23663,n23664);
  nand U25090(n23664,n23665,n23666);
  not U25091(n23663,n23667);
  nand U25092(n23661,n23665,n23666,n23667);
  nand U25093(G10212,n23668,n23669);
  nand U25094(n23669,n23670,n23671);
  nand U25095(n23671,n23672,n23673);
  not U25096(n23670,n23674);
  nand U25097(n23668,n23672,n23673,n23674);
  nand U25098(G10210,n23675,n23676);
  nand U25099(n23676,n23677,n23678);
  nand U25100(n23678,n23679,n23680);
  not U25101(n23677,n23681);
  nand U25102(n23675,n23679,n23680,n23681);
  nand U25103(G10208,n23682,n23683);
  nand U25104(n23683,n23684,n23685);
  nand U25105(n23685,n23686,n23687);
  not U25106(n23684,n23688);
  nand U25107(n23682,n23686,n23687,n23688);
  xor U25108(G10188,n23689,n23690);
  xor U25109(n23690,G36641,n23691);
  nand U25110(G10149,n23692,n23693);
  nand U25111(n23693,n23694,n13676);
  nand U25112(G10148,n23695,n23696);
  nand U25113(n23696,n23697,n23631,n23698);
  xor U25114(n23698,n23699,G36623);
  nand U25115(n23697,n23628,n23630);
  not U25116(n23628,n23632);
  nand U25117(n23695,n23700,n23630,n23701);
  xor U25118(n23701,n14016,n23699);
  nand U25119(n23699,n23702,n23703);
  nand U25120(n23703,n23704,n23705,n23706);
  xor U25121(n23706,G36378,G36133);
  nand U25122(n23705,n23707,n17696);
  nand U25123(n23702,n23707,n23708,n23709);
  xor U25124(n23709,n21535,G36378);
  not U25125(n21535,G36133);
  nand U25126(n23708,G36379,n23704);
  nand U25127(n23704,n23710,n21521);
  not U25128(n21521,G36134);
  nand U25129(n23707,G36134,n23711);
  not U25130(n14016,G36623);
  nand U25131(n23630,G36624,n23712);
  nand U25132(n23700,n23631,n23632);
  nand U25133(n23632,n23713,n23624);
  or U25134(n23624,n23714,n13879);
  nand U25135(n23713,n23625,n23623);
  nand U25136(n23623,n23714,n13879);
  not U25137(n13879,G36625);
  xnor U25138(n23714,n23715,n23716);
  xor U25139(n23716,G36380,G36135);
  nand U25140(n23625,n23717,n23617);
  or U25141(n23617,n23718,n13867);
  nand U25142(n23717,n23618,n23616);
  nand U25143(n23616,n13867,n23718);
  nand U25144(n23718,n23719,n23720,n23721);
  or U25145(n23721,n23722,n21496);
  nand U25146(n23720,n23723,n21496,n17671);
  nand U25147(n23719,G36381,n23724);
  nand U25148(n23724,n23725,n23726);
  nand U25149(n23726,G36136,n23723);
  not U25150(n23723,n23727);
  not U25151(n13867,G36626);
  nand U25152(n23618,n23728,n23610);
  nand U25153(n23610,G36627,n23729);
  nand U25154(n23728,n23611,n23609);
  or U25155(n23609,n23729,G36627);
  nand U25156(n23729,n23730,n23731);
  nand U25157(n23731,n23732,n23733);
  nand U25158(n23733,n23734,n23735);
  nand U25159(n23735,n21482,n17657);
  nand U25160(n23730,n23736,n23734);
  not U25161(n23734,n23737);
  nand U25162(n23611,n23738,n23603);
  or U25163(n23603,n23739,n13844);
  nand U25164(n23738,n23604,n23602);
  nand U25165(n23602,n23739,n13844);
  not U25166(n13844,G36628);
  xnor U25167(n23739,n23740,n23741);
  nor U25168(n23741,n23742,n23743);
  nand U25169(n23604,n23744,n23596);
  or U25170(n23596,n23745,n13832);
  nand U25171(n23744,n23597,n23595);
  nand U25172(n23595,n23745,n13832);
  not U25173(n13832,G36629);
  xnor U25174(n23745,n23746,n23747);
  xor U25175(n23747,G36384,G36139);
  nand U25176(n23597,n23748,n23589);
  nand U25177(n23589,G36630,n23749);
  nand U25178(n23748,n23590,n23588);
  or U25179(n23588,n23749,G36630);
  xnor U25180(n23749,n23750,n23751);
  xor U25181(n23751,G36385,G36140);
  nand U25182(n23590,n23752,n23582);
  nand U25183(n23582,G36631,n23753);
  nand U25184(n23752,n23583,n23581);
  or U25185(n23581,n23753,G36631);
  nand U25186(n23753,n23754,n23755);
  nand U25187(n23755,n23756,n23757);
  not U25188(n23756,n23758);
  nand U25189(n23754,n23759,n23760,n23761);
  xor U25190(n23761,n21426,G36386);
  nand U25191(n23760,G36387,n23762);
  nand U25192(n23583,n23763,n23575);
  nand U25193(n23575,n23764,G36632);
  nand U25194(n23763,n23576,n23574);
  or U25195(n23574,n23764,G36632);
  xnor U25196(n23764,n23765,n23766);
  xor U25197(n23766,G36387,G36142);
  nand U25198(n23576,n23767,n23687);
  or U25199(n23687,n23768,n13785);
  nand U25200(n23767,n23688,n23686);
  nand U25201(n23686,n23768,n13785);
  not U25202(n13785,G36633);
  xnor U25203(n23768,n23769,n23770);
  xor U25204(n23770,G36388,G36143);
  nand U25205(n23688,n23771,n23680);
  or U25206(n23680,n23772,n13773);
  nand U25207(n23771,n23681,n23679);
  nand U25208(n23679,n23772,n13773);
  not U25209(n13773,G36634);
  xor U25210(n23772,n23773,n23774);
  xor U25211(n23773,n17560,G36144);
  nand U25212(n23681,n23672,n23775);
  nand U25213(n23775,n23673,n23674);
  nand U25214(n23674,n23776,n23666);
  nand U25215(n23666,G36636,n23777);
  nand U25216(n23776,n23667,n23665);
  or U25217(n23665,n23777,G36636);
  xnor U25218(n23777,n23778,n23779);
  xor U25219(n23779,G36391,G36146);
  nand U25220(n23667,n23780,n23659);
  nand U25221(n23659,G36637,n23781);
  nand U25222(n23780,n23660,n23658);
  or U25223(n23658,n23781,G36637);
  xnor U25224(n23781,n23782,n23783);
  xor U25225(n23783,G36392,G36147);
  nand U25226(n23660,n23784,n23652);
  or U25227(n23652,n23785,n13728);
  nand U25228(n23784,n23653,n23651);
  nand U25229(n23651,n23785,n13728);
  not U25230(n13728,G36638);
  xnor U25231(n23785,n23786,n23787);
  xnor U25232(n23786,G36393,G36148);
  nand U25233(n23653,n23788,n23645);
  or U25234(n23645,n23789,n13716);
  nand U25235(n23788,n23646,n23644);
  nand U25236(n23644,n23789,n13716);
  not U25237(n13716,G36639);
  xnor U25238(n23789,n23790,n23791);
  xor U25239(n23791,G36394,G36149);
  nand U25240(n23646,n23637,n23792);
  nand U25241(n23792,n23639,n23638);
  or U25242(n23638,n23793,G36640);
  not U25243(n23639,n23636);
  nand U25244(n23636,n23794,n23795);
  nand U25245(n23795,n23796,n23797);
  not U25246(n23797,G36641);
  or U25247(n23796,n23692,n23689);
  nand U25248(n23794,n23689,n23692);
  not U25249(n23692,n23691);
  nor U25250(n23691,n23694,n13676);
  not U25251(n13676,G36642);
  xor U25252(n23694,G36152,G36397);
  xnor U25253(n23689,n23798,G36396);
  nand U25254(n23798,n23799,n23800);
  nand U25255(n23637,G36640,n23793);
  xnor U25256(n23793,n23801,n23802);
  xor U25257(n23802,G36395,G36150);
  or U25258(n23673,n23803,G36635);
  nand U25259(n23672,G36635,n23803);
  xnor U25260(n23803,n23804,n23805);
  xor U25261(n23805,G36390,G36145);
  or U25262(n23631,n23712,G36624);
  xnor U25263(n23712,n23806,n23710);
  not U25264(n23710,n23711);
  nand U25265(n23711,n23807,n23808);
  nand U25266(n23808,G36380,n23809);
  nand U25267(n23809,n21508,n23715);
  or U25268(n23807,n23715,n21508);
  not U25269(n21508,G36135);
  nand U25270(n23715,n23722,n23725,n23810);
  nand U25271(n23810,n21496,n17671);
  nand U25272(n23725,n23727,n21496);
  not U25273(n21496,G36136);
  nand U25274(n23722,n23727,n17671);
  not U25275(n17671,G36381);
  nor U25276(n23727,n23737,n23736);
  nor U25277(n23736,n23811,n23732);
  nor U25278(n23732,n23812,n23743);
  nor U25279(n23743,n21464,n17645);
  not U25280(n17645,G36383);
  not U25281(n21464,G36138);
  nor U25282(n23812,n23740,n23742);
  nor U25283(n23742,G36383,G36138);
  nand U25284(n23740,n23813,n23814);
  nand U25285(n23814,n23815,n17632);
  not U25286(n17632,G36384);
  or U25287(n23815,n23746,n21450);
  nand U25288(n23813,n23746,n21450);
  not U25289(n21450,G36139);
  nand U25290(n23746,n23816,n23817);
  nand U25291(n23817,n23818,n17619);
  not U25292(n17619,G36385);
  nand U25293(n23818,G36140,n23750);
  or U25294(n23816,n23750,G36140);
  nand U25295(n23750,n23758,n23757);
  nand U25296(n23757,G36141,G36386);
  nand U25297(n23758,n23762,n23819,n23820);
  nand U25298(n23820,n21426,n17601);
  not U25299(n17601,G36386);
  not U25300(n21426,G36141);
  nand U25301(n23819,n23759,n17587);
  not U25302(n17587,G36387);
  nand U25303(n23759,n23765,G36142);
  not U25304(n23765,n23821);
  nand U25305(n23762,n23821,n21408);
  not U25306(n21408,G36142);
  nand U25307(n23821,n23822,n23823);
  nand U25308(n23823,n23824,n17574);
  not U25309(n17574,G36388);
  or U25310(n23824,n23769,n21395);
  nand U25311(n23822,n23769,n21395);
  not U25312(n21395,G36143);
  nand U25313(n23769,n23825,n23826);
  nand U25314(n23826,n23827,n17560);
  not U25315(n17560,G36389);
  or U25316(n23827,n23774,n21381);
  nand U25317(n23825,n23774,n21381);
  not U25318(n21381,G36144);
  nand U25319(n23774,n23828,n23829);
  nand U25320(n23829,n23830,n17548);
  not U25321(n17548,G36390);
  nand U25322(n23830,G36145,n23804);
  or U25323(n23828,n23804,G36145);
  nand U25324(n23804,n23831,n23832);
  nand U25325(n23832,G36391,n23833);
  or U25326(n23833,n23778,G36146);
  nand U25327(n23831,G36146,n23778);
  nand U25328(n23778,n23834,n23835);
  nand U25329(n23835,G36392,n23836);
  or U25330(n23836,n23782,G36147);
  nand U25331(n23834,G36147,n23782);
  nand U25332(n23782,n23837,n23838);
  nand U25333(n23838,G36393,n23839);
  or U25334(n23839,G36148,n23787);
  nand U25335(n23837,n23787,G36148);
  and U25336(n23787,n23840,n23841);
  nand U25337(n23841,n23842,n17497);
  not U25338(n17497,G36394);
  or U25339(n23842,n23790,n21317);
  nand U25340(n23840,n23790,n21317);
  not U25341(n21317,G36149);
  nand U25342(n23790,n23843,n23844);
  nand U25343(n23844,n23845,n17484);
  not U25344(n17484,G36395);
  nand U25345(n23845,G36150,n23801);
  or U25346(n23843,n23801,G36150);
  nand U25347(n23801,n23800,n23846);
  nand U25348(n23846,G36396,n23799);
  nand U25349(n23799,n21286,n23847);
  nand U25350(n23847,G36152,G36397);
  not U25351(n21286,G36151);
  nand U25352(n23800,G36152,G36397,G36151);
  nor U25353(n23811,G36382,G36137);
  nor U25354(n23737,n21482,n17657);
  not U25355(n17657,G36382);
  not U25356(n21482,G36137);
  xor U25357(n23806,n17696,G36134);
  not U25358(n17696,G36379);
endmodule

