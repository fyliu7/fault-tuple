
module b17s_1 ( G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, 
        G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, 
        G29, G30, G31, G32, G33, G34, G35, G36, G37, G58839, G58840, G58841, 
        G58842, G58843, G58844, G58845, G58846, G58847, G58848, G58849, G58850, 
        G58851, G58852, G58853, G58854, G58855, G58856, G58857, G58858, G58859, 
        G58860, G58861, G58862, G58863, G58864, G58865, G58866, G58867, G58868, 
        G58869, G58870, G58871, G58872, G58873, G58874, G58875, G58876, G58877, 
        G58878, G58879, G58880, G58881, G58882, G58883, G58884, G58885, G58886, 
        G58887, G58888, G58889, G58890, G58891, G58892, G58893, G58894, G58895, 
        G58896, G58897, G58898, G58899, G58900, G58901, G58902, G58903, G58904, 
        G58905, G58906, G58907, G58908, G58909, G58910, G58911, G58912, G58913, 
        G58914, G58915, G58916, G58917, G58918, G58919, G58920, G58921, G58922, 
        G58923, G58924, G58925, G58926, G58927, G58928, G58929, G58930, G58931, 
        G58932, G58933, G58934, G58935, G58936, G58937, G58938, G58939, G58940, 
        G58941, G58942, G58943, G58944, G58945, G58946, G58947, G58948, G58949, 
        G58950, G58951, G58952, G58953, G58954, G58955, G58956, G58957, G58958, 
        G58959, G58960, G58961, G58962, G58963, G58964, G58965, G58966, G58967, 
        G58968, G58969, G58970, G58971, G58972, G58973, G58974, G58975, G58976, 
        G58977, G58978, G58979, G58980, G58981, G58982, G58983, G58984, G58985, 
        G58986, G58987, G58988, G58989, G58990, G58991, G58992, G58993, G58994, 
        G58995, G58996, G58997, G58998, G58999, G59000, G59001, G59002, G59003, 
        G59004, G59005, G59006, G59007, G59008, G59009, G59010, G59011, G59012, 
        G59013, G59014, G59015, G59016, G59017, G59018, G59019, G59020, G59021, 
        G59022, G59023, G59024, G59025, G59026, G59027, G59028, G59029, G59030, 
        G59031, G59032, G59033, G59034, G59035, G59036, G59037, G59038, G59039, 
        G59040, G59041, G59042, G59043, G59044, G59045, G59046, G59047, G59048, 
        G59049, G59050, G59051, G59052, G59053, G59054, G59055, G59056, G59057, 
        G59058, G59059, G59060, G59061, G59062, G59063, G59064, G59065, G59066, 
        G59067, G59068, G59069, G59070, G59071, G59072, G59073, G59074, G59075, 
        G59076, G59077, G59078, G59079, G59080, G59081, G59082, G59083, G59084, 
        G59085, G59086, G59087, G59088, G59089, G59090, G59091, G59092, G59093, 
        G59094, G59095, G59096, G59097, G59098, G59099, G59100, G59101, G59102, 
        G59103, G59104, G59105, G59106, G59107, G59108, G59109, G59110, G59111, 
        G59112, G59113, G59114, G59115, G59116, G59117, G59118, G59119, G59120, 
        G59121, G59122, G59123, G59124, G59125, G59126, G59127, G59128, G59129, 
        G59130, G59131, G59132, G59133, G59134, G59135, G59136, G59137, G59138, 
        G59139, G59140, G59141, G59142, G59143, G59144, G59145, G59146, G59147, 
        G59148, G59149, G59150, G59151, G59152, G59153, G59154, G59155, G59156, 
        G59157, G59158, G59159, G59160, G59161, G59162, G59163, G59164, G59165, 
        G59166, G59167, G59168, G59169, G59170, G59171, G59172, G59173, G59174, 
        G59175, G59176, G59177, G59178, G59179, G59180, G59181, G59182, G59183, 
        G59184, G59185, G59186, G59187, G59188, G59189, G59190, G59191, G59192, 
        G59193, G59194, G59195, G59196, G59197, G59198, G59199, G59200, G59201, 
        G59202, G59203, G59204, G59205, G59206, G59207, G59208, G59209, G59210, 
        G59211, G59212, G59213, G59214, G59215, G59216, G59217, G59218, G59219, 
        G59220, G59221, G59222, G59223, G59224, G59225, G59226, G59227, G59228, 
        G59229, G59230, G59231, G59232, G59233, G59234, G59235, G59236, G59237, 
        G59238, G59239, G59240, G59241, G59242, G59243, G59244, G59245, G59246, 
        G59247, G59248, G59249, G59250, G59251, G59252, G59253, G59254, G59255, 
        G59256, G59257, G59258, G59259, G59260, G59261, G59262, G59263, G59264, 
        G59265, G59266, G59267, G59268, G59269, G59270, G59271, G59272, G59273, 
        G59274, G59275, G59276, G59277, G59278, G59279, G59280, G59281, G59282, 
        G59283, G59284, G59285, G59286, G59287, G59288, G59289, G59290, G59291, 
        G59292, G59293, G59294, G59295, G59296, G59297, G59298, G59299, G59300, 
        G59301, G59302, G59303, G59304, G59305, G59306, G59307, G59308, G59309, 
        G59310, G59311, G59312, G59313, G59314, G59315, G59316, G59317, G59318, 
        G59319, G59320, G59321, G59322, G59323, G59324, G59325, G59326, G59327, 
        G59328, G59329, G59330, G59331, G59332, G59333, G59334, G59335, G59336, 
        G59337, G59338, G59339, G59340, G59341, G59342, G59343, G59344, G59345, 
        G59346, G59347, G59348, G59349, G59350, G59351, G59352, G59353, G59354, 
        G59355, G59356, G59357, G59358, G59359, G59360, G59361, G59362, G59363, 
        G59364, G59365, G59366, G59367, G59368, G59369, G59370, G59371, G59372, 
        G59373, G59374, G59375, G59376, G59377, G59378, G59379, G59380, G59381, 
        G59382, G59383, G59384, G59385, G59386, G59387, G59388, G59389, G59390, 
        G59391, G59392, G59393, G59394, G59395, G59396, G59397, G59398, G59399, 
        G59400, G59401, G59402, G59403, G59404, G59405, G59406, G59407, G59408, 
        G59409, G59410, G59411, G59412, G59413, G59414, G59415, G59416, G59417, 
        G59418, G59419, G59420, G59421, G59422, G59423, G59424, G59425, G59426, 
        G59427, G59428, G59429, G59430, G59431, G59432, G59433, G59434, G59435, 
        G59436, G59437, G59438, G59439, G59440, G59441, G59442, G59443, G59444, 
        G59445, G59446, G59447, G59448, G59449, G59450, G59451, G59452, G59453, 
        G59454, G59455, G59456, G59457, G59458, G59459, G59460, G59461, G59462, 
        G59463, G59464, G59465, G59466, G59467, G59468, G59469, G59470, G59471, 
        G59472, G59473, G59474, G59475, G59476, G59477, G59478, G59479, G59480, 
        G59481, G59482, G59483, G59484, G59485, G59486, G59487, G59488, G59489, 
        G59490, G59491, G59492, G59493, G59494, G59495, G59496, G59497, G59498, 
        G59499, G59500, G59501, G59502, G59503, G59504, G59505, G59506, G59507, 
        G59508, G59509, G59510, G59511, G59512, G59513, G59514, G59515, G59516, 
        G59517, G59518, G59519, G59520, G59521, G59522, G59523, G59524, G59525, 
        G59526, G59527, G59528, G59529, G59530, G59531, G59532, G59533, G59534, 
        G59535, G59536, G59537, G59538, G59539, G59540, G59541, G59542, G59543, 
        G59544, G59545, G59546, G59547, G59548, G59549, G59550, G59551, G59552, 
        G59553, G59554, G59555, G59556, G59557, G59558, G59559, G59560, G59561, 
        G59562, G59563, G59564, G59565, G59566, G59567, G59568, G59569, G59570, 
        G59571, G59572, G59573, G59574, G59575, G59576, G59577, G59578, G59579, 
        G59580, G59581, G59582, G59583, G59584, G59585, G59586, G59587, G59588, 
        G59589, G59590, G59591, G59592, G59593, G59594, G59595, G59596, G59597, 
        G59598, G59599, G59600, G59601, G59602, G59603, G59604, G59605, G59606, 
        G59607, G59608, G59609, G59610, G59611, G59612, G59613, G59614, G59615, 
        G59616, G59617, G59618, G59619, G59620, G59621, G59622, G59623, G59624, 
        G59625, G59626, G59627, G59628, G59629, G59630, G59631, G59632, G59633, 
        G59634, G59635, G59636, G59637, G59638, G59639, G59640, G59641, G59642, 
        G59643, G59644, G59645, G59646, G59647, G59648, G59649, G59650, G59651, 
        G59652, G59653, G59654, G59655, G59656, G59657, G59658, G59659, G59660, 
        G59661, G59662, G59663, G59664, G59665, G59666, G59667, G59668, G59669, 
        G59670, G59671, G59672, G59673, G59674, G59675, G59676, G59677, G59678, 
        G59679, G59680, G59681, G59682, G59683, G59684, G59685, G59686, G59687, 
        G59688, G59689, G59690, G59691, G59692, G59693, G59694, G59695, G59696, 
        G59697, G59698, G59699, G59700, G59701, G59702, G59703, G59704, G59705, 
        G59706, G59707, G59708, G59709, G59710, G59711, G59712, G59713, G59714, 
        G59715, G59716, G59717, G59718, G59719, G59720, G59721, G59722, G59723, 
        G59724, G59725, G59726, G59727, G59728, G59729, G59730, G59731, G59732, 
        G59733, G59734, G59735, G59736, G59737, G59738, G59739, G59740, G59741, 
        G59742, G59743, G59744, G59745, G59746, G59747, G59748, G59749, G59750, 
        G59751, G59752, G59753, G59754, G59755, G59756, G59757, G59758, G59759, 
        G59760, G59761, G59762, G59763, G59764, G59765, G59766, G59767, G59768, 
        G59769, G59770, G59771, G59772, G59773, G59774, G59775, G59776, G59777, 
        G59778, G59779, G59780, G59781, G59782, G59783, G59784, G59785, G59786, 
        G59787, G59788, G59789, G59790, G59791, G59792, G59793, G59794, G59795, 
        G59796, G59797, G59798, G59799, G59800, G59801, G59802, G59803, G59804, 
        G59805, G59806, G59807, G59808, G59809, G59810, G59811, G59812, G59813, 
        G59814, G59815, G59816, G59817, G59818, G59819, G59820, G59821, G59822, 
        G59823, G59824, G59825, G59826, G59827, G59828, G59829, G59830, G59831, 
        G59832, G59833, G59834, G59835, G59836, G59837, G59838, G59839, G59840, 
        G59841, G59842, G59843, G59844, G59845, G59846, G59847, G59848, G59849, 
        G59850, G59851, G59852, G59853, G59854, G59855, G59856, G59857, G59858, 
        G59859, G59860, G59861, G59862, G59863, G59864, G59865, G59866, G59867, 
        G59868, G59869, G59870, G59871, G59872, G59873, G59874, G59875, G59876, 
        G59877, G59878, G59879, G59880, G59881, G59882, G59883, G59884, G59885, 
        G59886, G59887, G59888, G59889, G59890, G59891, G59892, G59893, G59894, 
        G59895, G59896, G59897, G59898, G59899, G59900, G59901, G59902, G59903, 
        G59904, G59905, G59906, G59907, G59908, G59909, G59910, G59911, G59912, 
        G59913, G59914, G59915, G59916, G59917, G59918, G59919, G59920, G59921, 
        G59922, G59923, G59924, G59925, G59926, G59927, G59928, G59929, G59930, 
        G59931, G59932, G59933, G59934, G59935, G59936, G59937, G59938, G59939, 
        G59940, G59941, G59942, G59943, G59944, G59945, G59946, G59947, G59948, 
        G59949, G59950, G59951, G59952, G59953, G59954, G59955, G59956, G59957, 
        G59958, G59959, G59960, G59961, G59962, G59963, G59964, G59965, G59966, 
        G59967, G59968, G59969, G59970, G59971, G59972, G59973, G59974, G59975, 
        G59976, G59977, G59978, G59979, G59980, G59981, G59982, G59983, G59984, 
        G59985, G59986, G59987, G59988, G59989, G59990, G59991, G59992, G59993, 
        G59994, G59995, G59996, G59997, G59998, G59999, G60000, G60001, G60002, 
        G60003, G60004, G60005, G60006, G60007, G60008, G60009, G60010, G60011, 
        G60012, G60013, G60014, G60015, G60016, G60017, G60018, G60019, G60020, 
        G60021, G60022, G60023, G60024, G60025, G60026, G60027, G60028, G60029, 
        G60030, G60031, G60032, G60033, G60034, G60035, G60036, G60037, G60038, 
        G60039, G60040, G60041, G60042, G60043, G60044, G60045, G60046, G60047, 
        G60048, G60049, G60050, G60051, G60052, G60053, G60054, G60055, G60056, 
        G60057, G60058, G60059, G60060, G60061, G60062, G60063, G60064, G60065, 
        G60066, G60067, G60068, G60069, G60070, G60071, G60072, G60073, G60074, 
        G60075, G60076, G60077, G60078, G60079, G60080, G60081, G60082, G60083, 
        G60084, G60085, G60086, G60087, G60088, G60089, G60090, G60091, G60092, 
        G60093, G60094, G60095, G60096, G60097, G60098, G60099, G60100, G60101, 
        G60102, G60103, G60104, G60105, G60106, G60107, G60108, G60109, G60110, 
        G60111, G60112, G60113, G60114, G60115, G60116, G60117, G60118, G60119, 
        G60120, G60121, G60122, G60123, G60124, G60125, G60126, G60127, G60128, 
        G60129, G60130, G60131, G60132, G60133, G60134, G60135, G60136, G60137, 
        G60138, G60139, G60140, G60141, G60142, G60143, G60144, G60145, G60146, 
        G60147, G60148, G60149, G60150, G60151, G60152, G60153, G60154, G60155, 
        G60156, G60157, G60158, G60159, G60160, G60161, G60162, G60163, G60164, 
        G60165, G60166, G60167, G60168, G60169, G60170, G60171, G60172, G60173, 
        G60174, G60175, G60176, G60177, G60178, G60179, G60180, G60181, G60182, 
        G60183, G60184, G60185, G60186, G60187, G60188, G60189, G60190, G60191, 
        G60192, G60193, G60194, G60195, G60196, G60197, G60198, G60199, G60200, 
        G60201, G60202, G60203, G60204, G60205, G60206, G60207, G60208, G60209, 
        G60210, G60211, G60212, G60213, G60214, G60215, G60216, G60217, G60218, 
        G60219, G60220, G60221, G60222, G60223, G60224, G60225, G60226, G60227, 
        G60228, G60229, G60230, G60231, G60232, G60233, G60234, G60235, G60236, 
        G60237, G60238, G60239, G60240, G60241, G60242, G60243, G60244, G60245, 
        G60246, G60247, G60248, G60249, G60250, G60251, G60252, G60253, G1700, 
        G1701, G1702, G1703, G1704, G1705, G1706, G1707, G1708, G1709, G1711, 
        G1712, G1713, G1714, G1715, G1716, G1717, G1718, G1719, G1720, G1692, 
        G1693, G1694, G1695, G1696, G1697, G1698, G1699, G1710, G1721, G1556, 
        G1557, G1558, G1559, G1560, G1561, G1562, G1563, G1564, G1565, G1566, 
        G1567, G1568, G1569, G1570, G1571, G1572, G1573, G1574, G1575, G1576, 
        G1577, G1578, G1579, G1580, G1581, G1582, G1583, G1584, G1585, G1586, 
        G1587, G1596, G1597, G1598, G1599, G1600, G1601, G1602, G1603, G1604, 
        G1605, G1606, G1607, G1608, G1609, G1610, G1611, G1612, G1613, G1614, 
        G1615, G1616, G1617, G1618, G1619, G1620, G1621, G1622, G1623, G1624, 
        G1625, G1626, G1627, G1552, G1731, G1553, G1730, G3276, G3275, G3274, 
        G3273, G2314, G2315, G2316, G2317, G2318, G2319, G2320, G2321, G2322, 
        G2323, G2324, G2325, G2326, G2327, G2328, G2329, G2330, G2331, G2332, 
        G2333, G2334, G2335, G2336, G2337, G2338, G2339, G2340, G2341, G2342, 
        G2343, G2344, G2345, G2346, G3272, G3271, G2347, G2348, G2349, G2350, 
        G2351, G2352, G2353, G2354, G2355, G2356, G2357, G2358, G2359, G2360, 
        G2361, G2362, G2363, G2364, G2365, G2366, G2367, G2368, G2369, G2370, 
        G2371, G2372, G2373, G2374, G2375, G2376, G2377, G2378, G2379, G2380, 
        G2381, G2382, G2383, G2384, G2385, G2386, G2387, G2388, G2389, G2390, 
        G2391, G2392, G2393, G2394, G2395, G2396, G2397, G2398, G2399, G2400, 
        G2401, G2402, G2403, G2404, G2405, G2406, G2407, G2408, G2409, G2410, 
        G2411, G2412, G2413, G2414, G2415, G2416, G2417, G2418, G2419, G2420, 
        G2421, G2422, G2423, G2424, G2425, G2426, G2427, G2428, G2429, G2430, 
        G2431, G2432, G2433, G2434, G2435, G2436, G2437, G2438, G2439, G2440, 
        G2441, G2442, G2443, G2444, G2445, G2446, G2447, G2448, G2449, G2450, 
        G2451, G2452, G2453, G2454, G2455, G2456, G2457, G2458, G2459, G2460, 
        G2461, G2462, G2463, G2464, G2465, G2466, G2467, G2468, G2469, G2470, 
        G2471, G2472, G2473, G2474, G2475, G2476, G2477, G2478, G2479, G2480, 
        G2481, G2482, G2483, G2484, G2485, G2486, G2487, G2488, G2489, G2490, 
        G2491, G2492, G2493, G2494, G2495, G2496, G2497, G2498, G2499, G2500, 
        G2501, G2502, G2503, G2504, G2505, G2506, G2507, G2508, G3270, G3269, 
        G3268, G3266, G3265, G2509, G2510, G2511, G2512, G2747, G2513, G2514, 
        G2515, G2516, G2517, G2518, G2519, G2520, G2521, G2522, G2523, G2524, 
        G2525, G2526, G2527, G2528, G2529, G2530, G2531, G2532, G2533, G2534, 
        G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, 
        G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, 
        G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, 
        G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, 
        G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, 
        G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594, 
        G2595, G2596, G2597, G2598, G2599, G2600, G2601, G2602, G2603, G2604, 
        G2605, G2606, G2607, G2608, G2609, G2610, G2611, G2612, G2613, G2614, 
        G2615, G2616, G2617, G2618, G2619, G2620, G2621, G2622, G2623, G2624, 
        G2625, G2626, G2627, G2628, G2629, G2630, G2631, G2632, G2633, G2634, 
        G2635, G2636, G2637, G2638, G2639, G2640, G2641, G2642, G2643, G2644, 
        G2645, G2646, G2647, G2648, G2649, G2650, G2651, G2652, G2653, G2654, 
        G2655, G2656, G2657, G2658, G2659, G2660, G2661, G2662, G2663, G2664, 
        G2665, G2666, G2667, G2668, G2669, G2670, G2671, G2672, G2673, G2674, 
        G2675, G2676, G2677, G2678, G2679, G2680, G2681, G2682, G2683, G2684, 
        G2685, G2686, G2687, G2688, G2689, G2690, G2691, G2692, G2693, G2694, 
        G2695, G2696, G2697, G2698, G2699, G2700, G2701, G2702, G2703, G2704, 
        G2705, G2706, G2707, G2708, G2709, G2710, G2711, G2712, G2713, G2714, 
        G2715, G2716, G2717, G2718, G2719, G2720, G2721, G2722, G2723, G2724, 
        G2725, G2726, G2727, G2728, G2729, G2730, G2731, G2732, G2733, G2734, 
        G2735, G2736, G2737, G2738, G2739, G3264, G2740, G2741, G2742, G3263, 
        G2743, G3262, G2744, G2745, G3261, G3260, G9273, G9272, G9271, G9270, 
        G8311, G8312, G8313, G8314, G8315, G8316, G8317, G8318, G8319, G8320, 
        G8321, G8322, G8323, G8324, G8325, G8326, G8327, G8328, G8329, G8330, 
        G8331, G8332, G8333, G8334, G8335, G8336, G8337, G8338, G8339, G8340, 
        G8341, G8342, G8343, G9269, G9268, G8344, G8345, G8346, G8347, G8348, 
        G8349, G8350, G8351, G8352, G8353, G8354, G8355, G8356, G8357, G8358, 
        G8359, G8360, G8361, G8362, G8363, G8364, G8365, G8366, G8367, G8368, 
        G8369, G8370, G8371, G8372, G8373, G8374, G8375, G8376, G8377, G8378, 
        G8379, G8380, G8381, G8382, G8383, G8384, G8385, G8386, G8387, G8388, 
        G8389, G8390, G8391, G8392, G8393, G8394, G8395, G8396, G8397, G8398, 
        G8399, G8400, G8401, G8402, G8403, G8404, G8405, G8406, G8407, G8408, 
        G8409, G8410, G8411, G8412, G8413, G8414, G8415, G8416, G8417, G8418, 
        G8419, G8420, G8421, G8422, G8423, G8424, G8425, G8426, G8427, G8428, 
        G8429, G8430, G8431, G8432, G8433, G8434, G8435, G8436, G8437, G8438, 
        G8439, G8440, G8441, G8442, G8443, G8444, G8445, G8446, G8447, G8448, 
        G8449, G8450, G8451, G8452, G8453, G8454, G8455, G8456, G8457, G8458, 
        G8459, G8460, G8461, G8462, G8463, G8464, G8465, G8466, G8467, G8468, 
        G8469, G8470, G8471, G8472, G8473, G8474, G8475, G8476, G8477, G8478, 
        G8479, G8480, G8481, G8482, G8483, G8484, G8485, G8486, G8487, G8488, 
        G8489, G8490, G8491, G8492, G8493, G8494, G8495, G8496, G8497, G8498, 
        G8499, G8500, G8501, G8502, G8503, G8504, G8505, G9267, G9266, G9265, 
        G9263, G9262, G8506, G8507, G8508, G8509, G8744, G8510, G8511, G8512, 
        G8513, G8514, G8515, G8516, G8517, G8518, G8519, G8520, G8521, G8522, 
        G8523, G8524, G8525, G8526, G8527, G8528, G8529, G8530, G8531, G8532, 
        G8533, G8534, G8535, G8536, G8537, G8538, G8539, G8540, G8541, G8542, 
        G8543, G8544, G8545, G8546, G8547, G8548, G8549, G8550, G8551, G8552, 
        G8553, G8554, G8555, G8556, G8557, G8558, G8559, G8560, G8561, G8562, 
        G8563, G8564, G8565, G8566, G8567, G8568, G8569, G8570, G8571, G8572, 
        G8573, G8574, G8575, G8576, G8577, G8578, G8579, G8580, G8581, G8582, 
        G8583, G8584, G8585, G8586, G8587, G8588, G8589, G8590, G8591, G8592, 
        G8593, G8594, G8595, G8596, G8597, G8598, G8599, G8600, G8601, G8602, 
        G8603, G8604, G8605, G8606, G8607, G8608, G8609, G8610, G8611, G8612, 
        G8613, G8614, G8615, G8616, G8617, G8618, G8619, G8620, G8621, G8622, 
        G8623, G8624, G8625, G8626, G8627, G8628, G8629, G8630, G8631, G8632, 
        G8633, G8634, G8635, G8636, G8637, G8638, G8639, G8640, G8641, G8642, 
        G8643, G8644, G8645, G8646, G8647, G8648, G8649, G8650, G8651, G8652, 
        G8653, G8654, G8655, G8656, G8657, G8658, G8659, G8660, G8661, G8662, 
        G8663, G8664, G8665, G8666, G8667, G8668, G8669, G8670, G8671, G8672, 
        G8673, G8674, G8675, G8676, G8677, G8678, G8679, G8680, G8681, G8682, 
        G8683, G8684, G8685, G8686, G8687, G8688, G8689, G8690, G8691, G8692, 
        G8693, G8694, G8695, G8696, G8697, G8698, G8699, G8700, G8701, G8702, 
        G8703, G8704, G8705, G8706, G8707, G8708, G8709, G8710, G8711, G8712, 
        G8713, G8714, G8715, G8716, G8717, G8718, G8719, G8720, G8721, G8722, 
        G8723, G8724, G8725, G8726, G8727, G8728, G8729, G8730, G8731, G8732, 
        G8733, G8734, G8735, G8736, G9261, G8737, G8738, G8739, G9260, G8740, 
        G9259, G8741, G8742, G9258, G9257, G15270, G15269, G15268, G15267, 
        G14308, G14309, G14310, G14311, G14312, G14313, G14314, G14315, G14316, 
        G14317, G14318, G14319, G14320, G14321, G14322, G14323, G14324, G14325, 
        G14326, G14327, G14328, G14329, G14330, G14331, G14332, G14333, G14334, 
        G14335, G14336, G14337, G14338, G14339, G14340, G15266, G15265, G14341, 
        G14342, G14343, G14344, G14345, G14346, G14347, G14348, G14349, G14350, 
        G14351, G14352, G14353, G14354, G14355, G14356, G14357, G14358, G14359, 
        G14360, G14361, G14362, G14363, G14364, G14365, G14366, G14367, G14368, 
        G14369, G14370, G14371, G14372, G14373, G14374, G14375, G14376, G14377, 
        G14378, G14379, G14380, G14381, G14382, G14383, G14384, G14385, G14386, 
        G14387, G14388, G14389, G14390, G14391, G14392, G14393, G14394, G14395, 
        G14396, G14397, G14398, G14399, G14400, G14401, G14402, G14403, G14404, 
        G14405, G14406, G14407, G14408, G14409, G14410, G14411, G14412, G14413, 
        G14414, G14415, G14416, G14417, G14418, G14419, G14420, G14421, G14422, 
        G14423, G14424, G14425, G14426, G14427, G14428, G14429, G14430, G14431, 
        G14432, G14433, G14434, G14435, G14436, G14437, G14438, G14439, G14440, 
        G14441, G14442, G14443, G14444, G14445, G14446, G14447, G14448, G14449, 
        G14450, G14451, G14452, G14453, G14454, G14455, G14456, G14457, G14458, 
        G14459, G14460, G14461, G14462, G14463, G14464, G14465, G14466, G14467, 
        G14468, G14469, G14470, G14471, G14472, G14473, G14474, G14475, G14476, 
        G14477, G14478, G14479, G14480, G14481, G14482, G14483, G14484, G14485, 
        G14486, G14487, G14488, G14489, G14490, G14491, G14492, G14493, G14494, 
        G14495, G14496, G14497, G14498, G14499, G14500, G14501, G14502, G15264, 
        G15263, G15262, G15260, G15259, G14503, G14504, G14505, G14506, G14741, 
        G14507, G14508, G14509, G14510, G14511, G14512, G14513, G14514, G14515, 
        G14516, G14517, G14518, G14519, G14520, G14521, G14522, G14523, G14524, 
        G14525, G14526, G14527, G14528, G14529, G14530, G14531, G14532, G14533, 
        G14534, G14535, G14536, G14537, G14538, G14539, G14540, G14541, G14542, 
        G14543, G14544, G14545, G14546, G14547, G14548, G14549, G14550, G14551, 
        G14552, G14553, G14554, G14555, G14556, G14557, G14558, G14559, G14560, 
        G14561, G14562, G14563, G14564, G14565, G14566, G14567, G14568, G14569, 
        G14570, G14571, G14572, G14573, G14574, G14575, G14576, G14577, G14578, 
        G14579, G14580, G14581, G14582, G14583, G14584, G14585, G14586, G14587, 
        G14588, G14589, G14590, G14591, G14592, G14593, G14594, G14595, G14596, 
        G14597, G14598, G14599, G14600, G14601, G14602, G14603, G14604, G14605, 
        G14606, G14607, G14608, G14609, G14610, G14611, G14612, G14613, G14614, 
        G14615, G14616, G14617, G14618, G14619, G14620, G14621, G14622, G14623, 
        G14624, G14625, G14626, G14627, G14628, G14629, G14630, G14631, G14632, 
        G14633, G14634, G14635, G14636, G14637, G14638, G14639, G14640, G14641, 
        G14642, G14643, G14644, G14645, G14646, G14647, G14648, G14649, G14650, 
        G14651, G14652, G14653, G14654, G14655, G14656, G14657, G14658, G14659, 
        G14660, G14661, G14662, G14663, G14664, G14665, G14666, G14667, G14668, 
        G14669, G14670, G14671, G14672, G14673, G14674, G14675, G14676, G14677, 
        G14678, G14679, G14680, G14681, G14682, G14683, G14684, G14685, G14686, 
        G14687, G14688, G14689, G14690, G14691, G14692, G14693, G14694, G14695, 
        G14696, G14697, G14698, G14699, G14700, G14701, G14702, G14703, G14704, 
        G14705, G14706, G14707, G14708, G14709, G14710, G14711, G14712, G14713, 
        G14714, G14715, G14716, G14717, G14718, G14719, G14720, G14721, G14722, 
        G14723, G14724, G14725, G14726, G14727, G14728, G14729, G14730, G14731, 
        G14732, G14733, G15258, G14734, G14735, G14736, G15257, G14737, G15256, 
        G14738, G14739, G15255, G15254 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
         G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
         G31, G32, G33, G34, G35, G36, G37, G58839, G58840, G58841, G58842,
         G58843, G58844, G58845, G58846, G58847, G58848, G58849, G58850,
         G58851, G58852, G58853, G58854, G58855, G58856, G58857, G58858,
         G58859, G58860, G58861, G58862, G58863, G58864, G58865, G58866,
         G58867, G58868, G58869, G58870, G58871, G58872, G58873, G58874,
         G58875, G58876, G58877, G58878, G58879, G58880, G58881, G58882,
         G58883, G58884, G58885, G58886, G58887, G58888, G58889, G58890,
         G58891, G58892, G58893, G58894, G58895, G58896, G58897, G58898,
         G58899, G58900, G58901, G58902, G58903, G58904, G58905, G58906,
         G58907, G58908, G58909, G58910, G58911, G58912, G58913, G58914,
         G58915, G58916, G58917, G58918, G58919, G58920, G58921, G58922,
         G58923, G58924, G58925, G58926, G58927, G58928, G58929, G58930,
         G58931, G58932, G58933, G58934, G58935, G58936, G58937, G58938,
         G58939, G58940, G58941, G58942, G58943, G58944, G58945, G58946,
         G58947, G58948, G58949, G58950, G58951, G58952, G58953, G58954,
         G58955, G58956, G58957, G58958, G58959, G58960, G58961, G58962,
         G58963, G58964, G58965, G58966, G58967, G58968, G58969, G58970,
         G58971, G58972, G58973, G58974, G58975, G58976, G58977, G58978,
         G58979, G58980, G58981, G58982, G58983, G58984, G58985, G58986,
         G58987, G58988, G58989, G58990, G58991, G58992, G58993, G58994,
         G58995, G58996, G58997, G58998, G58999, G59000, G59001, G59002,
         G59003, G59004, G59005, G59006, G59007, G59008, G59009, G59010,
         G59011, G59012, G59013, G59014, G59015, G59016, G59017, G59018,
         G59019, G59020, G59021, G59022, G59023, G59024, G59025, G59026,
         G59027, G59028, G59029, G59030, G59031, G59032, G59033, G59034,
         G59035, G59036, G59037, G59038, G59039, G59040, G59041, G59042,
         G59043, G59044, G59045, G59046, G59047, G59048, G59049, G59050,
         G59051, G59052, G59053, G59054, G59055, G59056, G59057, G59058,
         G59059, G59060, G59061, G59062, G59063, G59064, G59065, G59066,
         G59067, G59068, G59069, G59070, G59071, G59072, G59073, G59074,
         G59075, G59076, G59077, G59078, G59079, G59080, G59081, G59082,
         G59083, G59084, G59085, G59086, G59087, G59088, G59089, G59090,
         G59091, G59092, G59093, G59094, G59095, G59096, G59097, G59098,
         G59099, G59100, G59101, G59102, G59103, G59104, G59105, G59106,
         G59107, G59108, G59109, G59110, G59111, G59112, G59113, G59114,
         G59115, G59116, G59117, G59118, G59119, G59120, G59121, G59122,
         G59123, G59124, G59125, G59126, G59127, G59128, G59129, G59130,
         G59131, G59132, G59133, G59134, G59135, G59136, G59137, G59138,
         G59139, G59140, G59141, G59142, G59143, G59144, G59145, G59146,
         G59147, G59148, G59149, G59150, G59151, G59152, G59153, G59154,
         G59155, G59156, G59157, G59158, G59159, G59160, G59161, G59162,
         G59163, G59164, G59165, G59166, G59167, G59168, G59169, G59170,
         G59171, G59172, G59173, G59174, G59175, G59176, G59177, G59178,
         G59179, G59180, G59181, G59182, G59183, G59184, G59185, G59186,
         G59187, G59188, G59189, G59190, G59191, G59192, G59193, G59194,
         G59195, G59196, G59197, G59198, G59199, G59200, G59201, G59202,
         G59203, G59204, G59205, G59206, G59207, G59208, G59209, G59210,
         G59211, G59212, G59245, G59246, G59247, G59248, G59249, G59250,
         G59251, G59252, G59253, G59254, G59255, G59256, G59257, G59258,
         G59259, G59260, G59261, G59262, G59263, G59264, G59265, G59266,
         G59267, G59268, G59269, G59270, G59271, G59272, G59273, G59274,
         G59275, G59276, G59277, G59278, G59279, G59280, G59281, G59282,
         G59283, G59284, G59285, G59286, G59287, G59288, G59289, G59290,
         G59291, G59292, G59293, G59294, G59295, G59296, G59297, G59298,
         G59299, G59300, G59301, G59302, G59303, G59304, G59305, G59306,
         G59307, G59308, G59309, G59310, G59311, G59312, G59313, G59314,
         G59315, G59316, G59317, G59318, G59319, G59320, G59321, G59322,
         G59323, G59324, G59325, G59326, G59327, G59328, G59329, G59330,
         G59331, G59332, G59333, G59334, G59335, G59336, G59337, G59338,
         G59339, G59340, G59341, G59342, G59343, G59344, G59346, G59347,
         G59348, G59349, G59352, G59354, G59355, G59356, G59357, G59358,
         G59359, G59360, G59361, G59362, G59363, G59364, G59365, G59366,
         G59367, G59368, G59369, G59370, G59371, G59372, G59373, G59374,
         G59375, G59376, G59377, G59378, G59379, G59380, G59381, G59382,
         G59383, G59384, G59385, G59386, G59387, G59388, G59389, G59390,
         G59391, G59392, G59393, G59394, G59395, G59396, G59397, G59398,
         G59399, G59400, G59401, G59402, G59403, G59404, G59405, G59406,
         G59407, G59408, G59409, G59410, G59411, G59412, G59413, G59414,
         G59415, G59416, G59417, G59418, G59419, G59420, G59421, G59422,
         G59423, G59424, G59425, G59426, G59427, G59428, G59429, G59430,
         G59431, G59432, G59433, G59434, G59435, G59436, G59437, G59438,
         G59439, G59440, G59441, G59442, G59443, G59444, G59445, G59446,
         G59447, G59448, G59449, G59450, G59451, G59452, G59453, G59454,
         G59455, G59456, G59457, G59458, G59459, G59460, G59461, G59462,
         G59463, G59464, G59465, G59466, G59467, G59468, G59469, G59470,
         G59471, G59472, G59473, G59474, G59475, G59476, G59477, G59478,
         G59479, G59480, G59481, G59482, G59483, G59484, G59485, G59486,
         G59487, G59488, G59489, G59490, G59491, G59492, G59493, G59494,
         G59495, G59496, G59497, G59498, G59499, G59500, G59501, G59502,
         G59503, G59504, G59505, G59506, G59507, G59508, G59509, G59510,
         G59511, G59512, G59513, G59514, G59515, G59516, G59517, G59518,
         G59519, G59520, G59521, G59522, G59523, G59524, G59525, G59526,
         G59527, G59528, G59529, G59530, G59531, G59532, G59533, G59534,
         G59535, G59536, G59537, G59538, G59539, G59540, G59541, G59542,
         G59543, G59544, G59545, G59546, G59547, G59548, G59549, G59550,
         G59551, G59552, G59553, G59554, G59555, G59556, G59557, G59558,
         G59559, G59560, G59561, G59562, G59563, G59564, G59565, G59566,
         G59567, G59568, G59569, G59570, G59571, G59572, G59573, G59574,
         G59575, G59576, G59577, G59578, G59579, G59580, G59581, G59582,
         G59583, G59584, G59585, G59586, G59587, G59588, G59589, G59590,
         G59591, G59592, G59593, G59594, G59595, G59596, G59597, G59598,
         G59599, G59600, G59601, G59602, G59603, G59604, G59605, G59606,
         G59607, G59608, G59609, G59610, G59611, G59612, G59613, G59614,
         G59615, G59616, G59617, G59618, G59619, G59620, G59621, G59622,
         G59623, G59624, G59625, G59626, G59627, G59628, G59629, G59630,
         G59631, G59632, G59633, G59634, G59635, G59636, G59637, G59638,
         G59639, G59640, G59641, G59642, G59643, G59644, G59645, G59646,
         G59647, G59648, G59649, G59650, G59651, G59652, G59653, G59654,
         G59655, G59656, G59657, G59658, G59659, G59660, G59661, G59662,
         G59663, G59664, G59665, G59666, G59667, G59668, G59669, G59670,
         G59671, G59672, G59673, G59674, G59675, G59676, G59677, G59678,
         G59679, G59680, G59681, G59682, G59683, G59684, G59685, G59686,
         G59687, G59688, G59689, G59690, G59691, G59692, G59693, G59694,
         G59695, G59696, G59697, G59698, G59699, G59700, G59701, G59702,
         G59703, G59704, G59705, G59706, G59707, G59708, G59709, G59710,
         G59711, G59712, G59713, G59714, G59715, G59716, G59717, G59718,
         G59719, G59720, G59721, G59722, G59723, G59724, G59725, G59726,
         G59727, G59728, G59729, G59730, G59731, G59732, G59733, G59734,
         G59735, G59736, G59737, G59738, G59739, G59740, G59741, G59742,
         G59743, G59744, G59745, G59746, G59747, G59748, G59749, G59750,
         G59751, G59752, G59753, G59754, G59755, G59756, G59757, G59758,
         G59759, G59760, G59761, G59762, G59763, G59764, G59765, G59766,
         G59767, G59768, G59769, G59770, G59771, G59772, G59773, G59774,
         G59775, G59776, G59777, G59778, G59779, G59780, G59781, G59782,
         G59783, G59784, G59785, G59786, G59787, G59788, G59789, G59790,
         G59791, G59792, G59793, G59794, G59795, G59796, G59797, G59798,
         G59799, G59800, G59801, G59802, G59803, G59804, G59805, G59806,
         G59807, G59808, G59839, G59840, G59841, G59842, G59843, G59844,
         G59845, G59846, G59847, G59848, G59849, G59850, G59851, G59852,
         G59853, G59854, G59855, G59856, G59857, G59858, G59859, G59860,
         G59861, G59862, G59863, G59864, G59865, G59866, G59867, G59868,
         G59869, G59870, G59871, G59872, G59873, G59874, G59875, G59876,
         G59877, G59878, G59879, G59880, G59881, G59882, G59883, G59884,
         G59885, G59886, G59887, G59888, G59889, G59890, G59891, G59892,
         G59893, G59894, G59895, G59896, G59897, G59898, G59899, G59900,
         G59901, G59902, G59903, G59904, G59905, G59906, G59907, G59908,
         G59909, G59910, G59911, G59912, G59913, G59914, G59915, G59916,
         G59917, G59918, G59919, G59920, G59921, G59922, G59923, G59924,
         G59925, G59926, G59927, G59928, G59929, G59930, G59931, G59932,
         G59933, G59934, G59935, G59936, G59937, G59938, G59939, G59940,
         G59941, G59942, G59943, G59944, G59945, G59946, G59947, G59948,
         G59949, G59950, G59951, G59952, G59953, G59954, G59955, G59956,
         G59957, G59958, G59959, G59960, G59961, G59962, G59963, G59964,
         G59965, G59966, G59967, G59968, G59969, G59970, G59971, G59972,
         G59973, G59974, G59975, G59976, G59977, G59978, G59979, G59980,
         G59981, G59982, G59983, G59984, G59985, G59986, G59987, G59988,
         G59989, G59990, G59991, G59992, G59993, G59994, G59995, G59996,
         G59997, G59998, G59999, G60000, G60001, G60002, G60003, G60004,
         G60005, G60006, G60007, G60008, G60009, G60010, G60011, G60012,
         G60013, G60014, G60015, G60016, G60017, G60018, G60019, G60020,
         G60021, G60022, G60023, G60024, G60025, G60026, G60027, G60028,
         G60029, G60030, G60031, G60032, G60033, G60034, G60035, G60036,
         G60037, G60038, G60039, G60040, G60041, G60042, G60043, G60044,
         G60045, G60046, G60047, G60048, G60049, G60050, G60051, G60052,
         G60053, G60054, G60055, G60056, G60057, G60058, G60059, G60060,
         G60061, G60062, G60063, G60064, G60065, G60066, G60067, G60068,
         G60069, G60070, G60071, G60072, G60073, G60074, G60075, G60076,
         G60077, G60078, G60079, G60080, G60081, G60082, G60083, G60084,
         G60085, G60086, G60087, G60088, G60089, G60090, G60091, G60092,
         G60093, G60094, G60095, G60096, G60097, G60098, G60099, G60100,
         G60101, G60102, G60103, G60104, G60105, G60106, G60107, G60108,
         G60109, G60110, G60111, G60112, G60113, G60114, G60115, G60116,
         G60117, G60118, G60119, G60120, G60121, G60122, G60123, G60124,
         G60125, G60126, G60127, G60128, G60129, G60130, G60131, G60132,
         G60133, G60134, G60135, G60136, G60137, G60138, G60139, G60140,
         G60141, G60142, G60143, G60144, G60145, G60146, G60147, G60148,
         G60149, G60150, G60151, G60152, G60153, G60154, G60155, G60156,
         G60157, G60158, G60159, G60160, G60161, G60162, G60163, G60164,
         G60165, G60166, G60167, G60168, G60169, G60170, G60171, G60172,
         G60173, G60174, G60175, G60176, G60177, G60178, G60179, G60180,
         G60181, G60182, G60183, G60184, G60185, G60186, G60187, G60188,
         G60189, G60190, G60191, G60192, G60193, G60194, G60195, G60196,
         G60197, G60198, G60199, G60200, G60201, G60202, G60203, G60204,
         G60205, G60206, G60207, G60208, G60209, G60210, G60211, G60212,
         G60213, G60214, G60215, G60216, G60217, G60218, G60219, G60220,
         G60221, G60222, G60223, G60224, G60225, G60226, G60227, G60228,
         G60229, G60230, G60231, G60232, G60233, G60234, G60235, G60236,
         G60237, G60238, G60239, G60240, G60241, G60242, G60243, G60244,
         G60245, G60246, G60247, G60248, G60249, G60250, G60252, G60253,
		 
G59213,  G59214,  G59215,  G59216,  G59217,  G59218,  G59219,  G59220, 
     G59221,  G59222,  G59223,  G59224,  G59225,  G59226,  G59227,  G59228, 
     G59229,  G59230,  G59231,  G59232,  G59233,  G59234,  G59235,  G59236, 
     G59237,  G59238,  G59239,  G59240,  G59241,  G59242,  G59243,  G59244, 
     G59345,  G59350,  G59351,  G59353,  G59809,  G59810,  G59811,  G59812, 
     G59813,  G59814,  G59815,  G59816,  G59817,  G59818,  G59819,  G59820, 
     G59821,  G59822,  G59823,  G59824,  G59825,  G59826,  G59827,  G59828, 
     G59829,  G59830,  G59831,  G59832,  G59833,  G59834,  G59835,  G59836, 
     G59837,  G59838,  G60251;
	 
  output G1700, G1701, G1702, G1703, G1704, G1705, G1706, G1707, G1708, G1709,
         G1711, G1712, G1713, G1714, G1715, G1716, G1717, G1718, G1719, G1720,
         G1692, G1693, G1694, G1695, G1696, G1697, G1698, G1699, G1710, G1721,
         G1556, G1557, G1558, G1559, G1560, G1561, G1562, G1563, G1564, G1565,
         G1566, G1567, G1568, G1569, G1570, G1571, G1572, G1573, G1574, G1575,
         G1576, G1577, G1578, G1579, G1580, G1581, G1582, G1583, G1584, G1585,
         G1586, G1587, G1596, G1597, G1598, G1599, G1600, G1601, G1602, G1603,
         G1604, G1605, G1606, G1607, G1608, G1609, G1610, G1611, G1612, G1613,
         G1614, G1615, G1616, G1617, G1618, G1619, G1620, G1621, G1622, G1623,
         G1624, G1625, G1626, G1627, G1552, G1731, G1553, G1730, G3276, G3275,
         G3274, G3273, G2314, G2315, G2316, G2317, G2318, G2319, G2320, G2321,
         G2322, G2323, G2324, G2325, G2326, G2327, G2328, G2329, G2330, G2331,
         G2332, G2333, G2334, G2335, G2336, G2337, G2338, G2339, G2340, G2341,
         G2342, G2343, G2344, G2345, G2346, G3272, G3271, G2347, G2348, G2349,
         G2350, G2351, G2352, G2353, G2354, G2355, G2356, G2357, G2358, G2359,
         G2360, G2361, G2362, G2363, G2364, G2365, G2366, G2367, G2368, G2369,
         G2370, G2371, G2372, G2373, G2374, G2375, G2376, G2377, G2378, G2379,
         G2380, G2381, G2382, G2383, G2384, G2385, G2386, G2387, G2388, G2389,
         G2390, G2391, G2392, G2393, G2394, G2395, G2396, G2397, G2398, G2399,
         G2400, G2401, G2402, G2403, G2404, G2405, G2406, G2407, G2408, G2409,
         G2410, G2411, G2412, G2413, G2414, G2415, G2416, G2417, G2418, G2419,
         G2420, G2421, G2422, G2423, G2424, G2425, G2426, G2427, G2428, G2429,
         G2430, G2431, G2432, G2433, G2434, G2435, G2436, G2437, G2438, G2439,
         G2440, G2441, G2442, G2443, G2444, G2445, G2446, G2447, G2448, G2449,
         G2450, G2451, G2452, G2453, G2454, G2455, G2456, G2457, G2458, G2459,
         G2460, G2461, G2462, G2463, G2464, G2465, G2466, G2467, G2468, G2469,
         G2470, G2471, G2472, G2473, G2474, G2475, G2476, G2477, G2478, G2479,
         G2480, G2481, G2482, G2483, G2484, G2485, G2486, G2487, G2488, G2489,
         G2490, G2491, G2492, G2493, G2494, G2495, G2496, G2497, G2498, G2499,
         G2500, G2501, G2502, G2503, G2504, G2505, G2506, G2507, G2508, G3270,
         G3269, G3268, G3266, G3265, G2509, G2510, G2511, G2512, G2747, G2513,
         G2514, G2515, G2516, G2517, G2518, G2519, G2520, G2521, G2522, G2523,
         G2524, G2525, G2526, G2527, G2528, G2529, G2530, G2531, G2532, G2533,
         G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543,
         G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553,
         G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563,
         G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573,
         G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583,
         G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593,
         G2594, G2595, G2596, G2597, G2598, G2599, G2600, G2601, G2602, G2603,
         G2604, G2605, G2606, G2607, G2608, G2609, G2610, G2611, G2612, G2613,
         G2614, G2615, G2616, G2617, G2618, G2619, G2620, G2621, G2622, G2623,
         G2624, G2625, G2626, G2627, G2628, G2629, G2630, G2631, G2632, G2633,
         G2634, G2635, G2636, G2637, G2638, G2639, G2640, G2641, G2642, G2643,
         G2644, G2645, G2646, G2647, G2648, G2649, G2650, G2651, G2652, G2653,
         G2654, G2655, G2656, G2657, G2658, G2659, G2660, G2661, G2662, G2663,
         G2664, G2665, G2666, G2667, G2668, G2669, G2670, G2671, G2672, G2673,
         G2674, G2675, G2676, G2677, G2678, G2679, G2680, G2681, G2682, G2683,
         G2684, G2685, G2686, G2687, G2688, G2689, G2690, G2691, G2692, G2693,
         G2694, G2695, G2696, G2697, G2698, G2699, G2700, G2701, G2702, G2703,
         G2704, G2705, G2706, G2707, G2708, G2709, G2710, G2711, G2712, G2713,
         G2714, G2715, G2716, G2717, G2718, G2719, G2720, G2721, G2722, G2723,
         G2724, G2725, G2726, G2727, G2728, G2729, G2730, G2731, G2732, G2733,
         G2734, G2735, G2736, G2737, G2738, G2739, G3264, G2740, G2741, G2742,
         G3263, G2743, G3262, G2744, G2745, G3261, G3260, G9273, G9272, G9271,
         G9270, G8311, G8312, G8313, G8314, G8315, G8316, G8317, G8318, G8319,
         G8320, G8321, G8322, G8323, G8324, G8325, G8326, G8327, G8328, G8329,
         G8330, G8331, G8332, G8333, G8334, G8335, G8336, G8337, G8338, G8339,
         G8340, G8341, G8342, G8343, G9269, G9268, G8344, G8345, G8346, G8347,
         G8348, G8349, G8350, G8351, G8352, G8353, G8354, G8355, G8356, G8357,
         G8358, G8359, G8360, G8361, G8362, G8363, G8364, G8365, G8366, G8367,
         G8368, G8369, G8370, G8371, G8372, G8373, G8374, G8375, G8376, G8377,
         G8378, G8379, G8380, G8381, G8382, G8383, G8384, G8385, G8386, G8387,
         G8388, G8389, G8390, G8391, G8392, G8393, G8394, G8395, G8396, G8397,
         G8398, G8399, G8400, G8401, G8402, G8403, G8404, G8405, G8406, G8407,
         G8408, G8409, G8410, G8411, G8412, G8413, G8414, G8415, G8416, G8417,
         G8418, G8419, G8420, G8421, G8422, G8423, G8424, G8425, G8426, G8427,
         G8428, G8429, G8430, G8431, G8432, G8433, G8434, G8435, G8436, G8437,
         G8438, G8439, G8440, G8441, G8442, G8443, G8444, G8445, G8446, G8447,
         G8448, G8449, G8450, G8451, G8452, G8453, G8454, G8455, G8456, G8457,
         G8458, G8459, G8460, G8461, G8462, G8463, G8464, G8465, G8466, G8467,
         G8468, G8469, G8470, G8471, G8472, G8473, G8474, G8475, G8476, G8477,
         G8478, G8479, G8480, G8481, G8482, G8483, G8484, G8485, G8486, G8487,
         G8488, G8489, G8490, G8491, G8492, G8493, G8494, G8495, G8496, G8497,
         G8498, G8499, G8500, G8501, G8502, G8503, G8504, G8505, G9267, G9266,
         G9265, G9263, G9262, G8506, G8507, G8508, G8509, G8744, G8510, G8511,
         G8512, G8513, G8514, G8515, G8516, G8517, G8518, G8519, G8520, G8521,
         G8522, G8523, G8524, G8525, G8526, G8527, G8528, G8529, G8530, G8531,
         G8532, G8533, G8534, G8535, G8536, G8537, G8538, G8539, G8540, G8541,
         G8542, G8543, G8544, G8545, G8546, G8547, G8548, G8549, G8550, G8551,
         G8552, G8553, G8554, G8555, G8556, G8557, G8558, G8559, G8560, G8561,
         G8562, G8563, G8564, G8565, G8566, G8567, G8568, G8569, G8570, G8571,
         G8572, G8573, G8574, G8575, G8576, G8577, G8578, G8579, G8580, G8581,
         G8582, G8583, G8584, G8585, G8586, G8587, G8588, G8589, G8590, G8591,
         G8592, G8593, G8594, G8595, G8596, G8597, G8598, G8599, G8600, G8601,
         G8602, G8603, G8604, G8605, G8606, G8607, G8608, G8609, G8610, G8611,
         G8612, G8613, G8614, G8615, G8616, G8617, G8618, G8619, G8620, G8621,
         G8622, G8623, G8624, G8625, G8626, G8627, G8628, G8629, G8630, G8631,
         G8632, G8633, G8634, G8635, G8636, G8637, G8638, G8639, G8640, G8641,
         G8642, G8643, G8644, G8645, G8646, G8647, G8648, G8649, G8650, G8651,
         G8652, G8653, G8654, G8655, G8656, G8657, G8658, G8659, G8660, G8661,
         G8662, G8663, G8664, G8665, G8666, G8667, G8668, G8669, G8670, G8671,
         G8672, G8673, G8674, G8675, G8676, G8677, G8678, G8679, G8680, G8681,
         G8682, G8683, G8684, G8685, G8686, G8687, G8688, G8689, G8690, G8691,
         G8692, G8693, G8694, G8695, G8696, G8697, G8698, G8699, G8700, G8701,
         G8702, G8703, G8704, G8705, G8706, G8707, G8708, G8709, G8710, G8711,
         G8712, G8713, G8714, G8715, G8716, G8717, G8718, G8719, G8720, G8721,
         G8722, G8723, G8724, G8725, G8726, G8727, G8728, G8729, G8730, G8731,
         G8732, G8733, G8734, G8735, G8736, G9261, G8737, G8738, G8739, G9260,
         G8740, G9259, G8741, G8742, G9258, G9257, G15270, G15269, G15268,
         G15267, G14308, G14309, G14310, G14311, G14312, G14313, G14314,
         G14315, G14316, G14317, G14318, G14319, G14320, G14321, G14322,
         G14323, G14324, G14325, G14326, G14327, G14328, G14329, G14330,
         G14331, G14332, G14333, G14334, G14335, G14336, G14337, G14338,
         G14339, G14340, G15266, G15265, G14341, G14342, G14343, G14344,
         G14345, G14346, G14347, G14348, G14349, G14350, G14351, G14352,
         G14353, G14354, G14355, G14356, G14357, G14358, G14359, G14360,
         G14361, G14362, G14363, G14364, G14365, G14366, G14367, G14368,
         G14369, G14370, G14371, G14372, G14373, G14374, G14375, G14376,
         G14377, G14378, G14379, G14380, G14381, G14382, G14383, G14384,
         G14385, G14386, G14387, G14388, G14389, G14390, G14391, G14392,
         G14393, G14394, G14395, G14396, G14397, G14398, G14399, G14400,
         G14401, G14402, G14403, G14404, G14405, G14406, G14407, G14408,
         G14409, G14410, G14411, G14412, G14413, G14414, G14415, G14416,
         G14417, G14418, G14419, G14420, G14421, G14422, G14423, G14424,
         G14425, G14426, G14427, G14428, G14429, G14430, G14431, G14432,
         G14433, G14434, G14435, G14436, G14437, G14438, G14439, G14440,
         G14441, G14442, G14443, G14444, G14445, G14446, G14447, G14448,
         G14449, G14450, G14451, G14452, G14453, G14454, G14455, G14456,
         G14457, G14458, G14459, G14460, G14461, G14462, G14463, G14464,
         G14465, G14466, G14467, G14468, G14469, G14470, G14471, G14472,
         G14473, G14474, G14475, G14476, G14477, G14478, G14479, G14480,
         G14481, G14482, G14483, G14484, G14485, G14486, G14487, G14488,
         G14489, G14490, G14491, G14492, G14493, G14494, G14495, G14496,
         G14497, G14498, G14499, G14500, G14501, G14502, G15264, G15263,
         G15262, G15260, G15259, G14503, G14504, G14505, G14506, G14741,
         G14507, G14508, G14509, G14510, G14511, G14512, G14513, G14514,
         G14515, G14516, G14517, G14518, G14519, G14520, G14521, G14522,
         G14523, G14524, G14525, G14526, G14527, G14528, G14529, G14530,
         G14531, G14532, G14533, G14534, G14535, G14536, G14537, G14538,
         G14539, G14540, G14541, G14542, G14543, G14544, G14545, G14546,
         G14547, G14548, G14549, G14550, G14551, G14552, G14553, G14554,
         G14555, G14556, G14557, G14558, G14559, G14560, G14561, G14562,
         G14563, G14564, G14565, G14566, G14567, G14568, G14569, G14570,
         G14571, G14572, G14573, G14574, G14575, G14576, G14577, G14578,
         G14579, G14580, G14581, G14582, G14583, G14584, G14585, G14586,
         G14587, G14588, G14589, G14590, G14591, G14592, G14593, G14594,
         G14595, G14596, G14597, G14598, G14599, G14600, G14601, G14602,
         G14603, G14604, G14605, G14606, G14607, G14608, G14609, G14610,
         G14611, G14612, G14613, G14614, G14615, G14616, G14617, G14618,
         G14619, G14620, G14621, G14622, G14623, G14624, G14625, G14626,
         G14627, G14628, G14629, G14630, G14631, G14632, G14633, G14634,
         G14635, G14636, G14637, G14638, G14639, G14640, G14641, G14642,
         G14643, G14644, G14645, G14646, G14647, G14648, G14649, G14650,
         G14651, G14652, G14653, G14654, G14655, G14656, G14657, G14658,
         G14659, G14660, G14661, G14662, G14663, G14664, G14665, G14666,
         G14667, G14668, G14669, G14670, G14671, G14672, G14673, G14674,
         G14675, G14676, G14677, G14678, G14679, G14680, G14681, G14682,
         G14683, G14684, G14685, G14686, G14687, G14688, G14689, G14690,
         G14691, G14692, G14693, G14694, G14695, G14696, G14697, G14698,
         G14699, G14700, G14701, G14702, G14703, G14704, G14705, G14706,
         G14707, G14708, G14709, G14710, G14711, G14712, G14713, G14714,
         G14715, G14716, G14717, G14718, G14719, G14720, G14721, G14722,
         G14723, G14724, G14725, G14726, G14727, G14728, G14729, G14730,
         G14731, G14732, G14733, G15258, G14734, G14735, G14736, G15257,
         G14737, G15256, G14738, G14739, G15255, G15254;

  wire   n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
         n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
         n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135,
         n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
         n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151,
         n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159,
         n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167,
         n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
         n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183,
         n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
         n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
         n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207,
         n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
         n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223,
         n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231,
         n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
         n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247,
         n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255,
         n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
         n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
         n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279,
         n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
         n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295,
         n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
         n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311,
         n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319,
         n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327,
         n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
         n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
         n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351,
         n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
         n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
         n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847,
         n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855,
         n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863,
         n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
         n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879,
         n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
         n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895,
         n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903,
         n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
         n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919,
         n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927,
         n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935,
         n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
         n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951,
         n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
         n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967,
         n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975,
         n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
         n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991,
         n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999,
         n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007,
         n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
         n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023,
         n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
         n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039,
         n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047,
         n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
         n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063,
         n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071,
         n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079,
         n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
         n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095,
         n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
         n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111,
         n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119,
         n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
         n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135,
         n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143,
         n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151,
         n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
         n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167,
         n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
         n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183,
         n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191,
         n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
         n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207,
         n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215,
         n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223,
         n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
         n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239,
         n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247,
         n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255,
         n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263,
         n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
         n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279,
         n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287,
         n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295,
         n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
         n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
         n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319,
         n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327,
         n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335,
         n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
         n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351,
         n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359,
         n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367,
         n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
         n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
         n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391,
         n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399,
         n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407,
         n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
         n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423,
         n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431,
         n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439,
         n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
         n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
         n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463,
         n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471,
         n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479,
         n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
         n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495,
         n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503,
         n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511,
         n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
         n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
         n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535,
         n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543,
         n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551,
         n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
         n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567,
         n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575,
         n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583,
         n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
         n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
         n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607,
         n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615,
         n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
         n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631,
         n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639,
         n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647,
         n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655,
         n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
         n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
         n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679,
         n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687,
         n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
         n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703,
         n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
         n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719,
         n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727,
         n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
         n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743,
         n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751,
         n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759,
         n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
         n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
         n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783,
         n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791,
         n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799,
         n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
         n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815,
         n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823,
         n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831,
         n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
         n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
         n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855,
         n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863,
         n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871,
         n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
         n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887,
         n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895,
         n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903,
         n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
         n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919,
         n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927,
         n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935,
         n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943,
         n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
         n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959,
         n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967,
         n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975,
         n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
         n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991,
         n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999,
         n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
         n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015,
         n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
         n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031,
         n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039,
         n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047,
         n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
         n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063,
         n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071,
         n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
         n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087,
         n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
         n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103,
         n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111,
         n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119,
         n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
         n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135,
         n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143,
         n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
         n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159,
         n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
         n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175,
         n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183,
         n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191,
         n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
         n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207,
         n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
         n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223,
         n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231,
         n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
         n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247,
         n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255,
         n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263,
         n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
         n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279,
         n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
         n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295,
         n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303,
         n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311,
         n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319,
         n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327,
         n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335,
         n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
         n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351,
         n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359,
         n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367,
         n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375,
         n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383,
         n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391,
         n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399,
         n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
         n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
         n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423,
         n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431,
         n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439,
         n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447,
         n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455,
         n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
         n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471,
         n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479,
         n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
         n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495,
         n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503,
         n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511,
         n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519,
         n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527,
         n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535,
         n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543,
         n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
         n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
         n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567,
         n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
         n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583,
         n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591,
         n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599,
         n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607,
         n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615,
         n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
         n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
         n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639,
         n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
         n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655,
         n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663,
         n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671,
         n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679,
         n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687,
         n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
         n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
         n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711,
         n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
         n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727,
         n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735,
         n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743,
         n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751,
         n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
         n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767,
         n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
         n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783,
         n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791,
         n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799,
         n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807,
         n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815,
         n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823,
         n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
         n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839,
         n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
         n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855,
         n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863,
         n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871,
         n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879,
         n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887,
         n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895,
         n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
         n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911,
         n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
         n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927,
         n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935,
         n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943,
         n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951,
         n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959,
         n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
         n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
         n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983,
         n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
         n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999,
         n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007,
         n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015,
         n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023,
         n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031,
         n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
         n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
         n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055,
         n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
         n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071,
         n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079,
         n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087,
         n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095,
         n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103,
         n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111,
         n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
         n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127,
         n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
         n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143,
         n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151,
         n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159,
         n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167,
         n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
         n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183,
         n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
         n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199,
         n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
         n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215,
         n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223,
         n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231,
         n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239,
         n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
         n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255,
         n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
         n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271,
         n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
         n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287,
         n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295,
         n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303,
         n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
         n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319,
         n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327,
         n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
         n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343,
         n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
         n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359,
         n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367,
         n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375,
         n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
         n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391,
         n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399,
         n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
         n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
         n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423,
         n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431,
         n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439,
         n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447,
         n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455,
         n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463,
         n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471,
         n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
         n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
         n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495,
         n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503,
         n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511,
         n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
         n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527,
         n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535,
         n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543,
         n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
         n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
         n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567,
         n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575,
         n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583,
         n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
         n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599,
         n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607,
         n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615,
         n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623,
         n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
         n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639,
         n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647,
         n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655,
         n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663,
         n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671,
         n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679,
         n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687,
         n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695,
         n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
         n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711,
         n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719,
         n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
         n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735,
         n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743,
         n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751,
         n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759,
         n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767,
         n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
         n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783,
         n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791,
         n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
         n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807,
         n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815,
         n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
         n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831,
         n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839,
         n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
         n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855,
         n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
         n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871,
         n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879,
         n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887,
         n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
         n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903,
         n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911,
         n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
         n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927,
         n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
         n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943,
         n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951,
         n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959,
         n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
         n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975,
         n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983,
         n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
         n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
         n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007,
         n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015,
         n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
         n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031,
         n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039,
         n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047,
         n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055,
         n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
         n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
         n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079,
         n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087,
         n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095,
         n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103,
         n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111,
         n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119,
         n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
         n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
         n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143,
         n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151,
         n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159,
         n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167,
         n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175,
         n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183,
         n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191,
         n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
         n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
         n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215,
         n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223,
         n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231,
         n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239,
         n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247,
         n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255,
         n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263,
         n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
         n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
         n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287,
         n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295,
         n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303,
         n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311,
         n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319,
         n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327,
         n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335,
         n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
         n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
         n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359,
         n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367,
         n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375,
         n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383,
         n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391,
         n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399,
         n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
         n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415,
         n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
         n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431,
         n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439,
         n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447,
         n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455,
         n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463,
         n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
         n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
         n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487,
         n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
         n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503,
         n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511,
         n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519,
         n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527,
         n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535,
         n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
         n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551,
         n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559,
         n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
         n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575,
         n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583,
         n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591,
         n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599,
         n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607,
         n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
         n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623,
         n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631,
         n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
         n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647,
         n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655,
         n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663,
         n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671,
         n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
         n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
         n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695,
         n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703,
         n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
         n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719,
         n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727,
         n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735,
         n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743,
         n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
         n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759,
         n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767,
         n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775,
         n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
         n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791,
         n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799,
         n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807,
         n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
         n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
         n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831,
         n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839,
         n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847,
         n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
         n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863,
         n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871,
         n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879,
         n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887,
         n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
         n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903,
         n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911,
         n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919,
         n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
         n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935,
         n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943,
         n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
         n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
         n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967,
         n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975,
         n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983,
         n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991,
         n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
         n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007,
         n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
         n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023,
         n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
         n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039,
         n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047,
         n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055,
         n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063,
         n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
         n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079,
         n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087,
         n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095,
         n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
         n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111,
         n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119,
         n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
         n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135,
         n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
         n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151,
         n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159,
         n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167,
         n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
         n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183,
         n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191,
         n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
         n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
         n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215,
         n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223,
         n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231,
         n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
         n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247,
         n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255,
         n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
         n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271,
         n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
         n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287,
         n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295,
         n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303,
         n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
         n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319,
         n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
         n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335,
         n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343,
         n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
         n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359,
         n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367,
         n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375,
         n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
         n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391,
         n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399,
         n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407,
         n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415,
         n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
         n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431,
         n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439,
         n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447,
         n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
         n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463,
         n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471,
         n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479,
         n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
         n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495,
         n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503,
         n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511,
         n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519,
         n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527,
         n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535,
         n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543,
         n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
         n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559,
         n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567,
         n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575,
         n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
         n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591,
         n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
         n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607,
         n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615,
         n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623,
         n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631,
         n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639,
         n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647,
         n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655,
         n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663,
         n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
         n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679,
         n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687,
         n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695,
         n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703,
         n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711,
         n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719,
         n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727,
         n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735,
         n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
         n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751,
         n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759,
         n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767,
         n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775,
         n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783,
         n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791,
         n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799,
         n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807,
         n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
         n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823,
         n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831,
         n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839,
         n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847,
         n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
         n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863,
         n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871,
         n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879,
         n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
         n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895,
         n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903,
         n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911,
         n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919,
         n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
         n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935,
         n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943,
         n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951,
         n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
         n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967,
         n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975,
         n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983,
         n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991,
         n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
         n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007,
         n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015,
         n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023,
         n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
         n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039,
         n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047,
         n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055,
         n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063,
         n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
         n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079,
         n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087,
         n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095,
         n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103,
         n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111,
         n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119,
         n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127,
         n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135,
         n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
         n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151,
         n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159,
         n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
         n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175,
         n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183,
         n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191,
         n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199,
         n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207,
         n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
         n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223,
         n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231,
         n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
         n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247,
         n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255,
         n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263,
         n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271,
         n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279,
         n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287,
         n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295,
         n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
         n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311,
         n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319,
         n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327,
         n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335,
         n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343,
         n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351,
         n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359,
         n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367,
         n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
         n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383,
         n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391,
         n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399,
         n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407,
         n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415,
         n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423,
         n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431,
         n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439,
         n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
         n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455,
         n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463,
         n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471,
         n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479,
         n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487,
         n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495,
         n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
         n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511,
         n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
         n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527,
         n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535,
         n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543,
         n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551,
         n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559,
         n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567,
         n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
         n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
         n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591,
         n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599,
         n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607,
         n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615,
         n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623,
         n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631,
         n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639,
         n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
         n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
         n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663,
         n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671,
         n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679,
         n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687,
         n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695,
         n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703,
         n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711,
         n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
         n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
         n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735,
         n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743,
         n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751,
         n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759,
         n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767,
         n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775,
         n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783,
         n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
         n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799,
         n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807,
         n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815,
         n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823,
         n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831,
         n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839,
         n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847,
         n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855,
         n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
         n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871,
         n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879,
         n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887,
         n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895,
         n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903,
         n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911,
         n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919,
         n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927,
         n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
         n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943,
         n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951,
         n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959,
         n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967,
         n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975,
         n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983,
         n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991,
         n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999,
         n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
         n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015,
         n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023,
         n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031,
         n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039,
         n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047,
         n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055,
         n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063,
         n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
         n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079,
         n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087,
         n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095,
         n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103,
         n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111,
         n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119,
         n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127,
         n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135,
         n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
         n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151,
         n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159,
         n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167,
         n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175,
         n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183,
         n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191,
         n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199,
         n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207,
         n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
         n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223,
         n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231,
         n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239,
         n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247,
         n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255,
         n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263,
         n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271,
         n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279,
         n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
         n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295,
         n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303,
         n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311,
         n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319,
         n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327,
         n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335,
         n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343,
         n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
         n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
         n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367,
         n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375,
         n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383,
         n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391,
         n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399,
         n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407,
         n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415,
         n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
         n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
         n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439,
         n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447,
         n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455,
         n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463,
         n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471,
         n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479,
         n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487,
         n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
         n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
         n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511,
         n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519,
         n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527,
         n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535,
         n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543,
         n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551,
         n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
         n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567,
         n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
         n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583,
         n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591,
         n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599,
         n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607,
         n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615,
         n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623,
         n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
         n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639,
         n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
         n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655,
         n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663,
         n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671,
         n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679,
         n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687,
         n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695,
         n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703,
         n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711,
         n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
         n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727,
         n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735,
         n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743,
         n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751,
         n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759,
         n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767,
         n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775,
         n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783,
         n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
         n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799,
         n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807,
         n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815,
         n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823,
         n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831,
         n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
         n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847,
         n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855,
         n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
         n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871,
         n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879,
         n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887,
         n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895,
         n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903,
         n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
         n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919,
         n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927,
         n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
         n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943,
         n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951,
         n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959,
         n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967,
         n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975,
         n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
         n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991,
         n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999,
         n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
         n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015,
         n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023,
         n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031,
         n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039,
         n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
         n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055,
         n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063,
         n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071,
         n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
         n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087,
         n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095,
         n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103,
         n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111,
         n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
         n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127,
         n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135,
         n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143,
         n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
         n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159,
         n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167,
         n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175,
         n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183,
         n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
         n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199,
         n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207,
         n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215,
         n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
         n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231,
         n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239,
         n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247,
         n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255,
         n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263,
         n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271,
         n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279,
         n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287,
         n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
         n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303,
         n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311,
         n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319,
         n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327,
         n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335,
         n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343,
         n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351,
         n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359,
         n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
         n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375,
         n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383,
         n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391,
         n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399,
         n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407,
         n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415,
         n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423,
         n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431,
         n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
         n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447,
         n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455,
         n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463,
         n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471,
         n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479,
         n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487,
         n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495,
         n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503,
         n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
         n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519,
         n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527,
         n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535,
         n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543,
         n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551,
         n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559,
         n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567,
         n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575,
         n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
         n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591,
         n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599,
         n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607,
         n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615,
         n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623,
         n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631,
         n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
         n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647,
         n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
         n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663,
         n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671,
         n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679,
         n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687,
         n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695,
         n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703,
         n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711,
         n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719,
         n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
         n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735,
         n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743,
         n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
         n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759,
         n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767,
         n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775,
         n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783,
         n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791,
         n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
         n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807,
         n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815,
         n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823,
         n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831,
         n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839,
         n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847,
         n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855,
         n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863,
         n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
         n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879,
         n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887,
         n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895,
         n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903,
         n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911,
         n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919,
         n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927,
         n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935,
         n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
         n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951,
         n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959,
         n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967,
         n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975,
         n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983,
         n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991,
         n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999,
         n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007,
         n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015,
         n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023,
         n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031,
         n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039,
         n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047,
         n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055,
         n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063,
         n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
         n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
         n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087,
         n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095,
         n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103,
         n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111,
         n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119,
         n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127,
         n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135,
         n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
         n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
         n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159,
         n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167,
         n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175,
         n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183,
         n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191,
         n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199,
         n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207,
         n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
         n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
         n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231,
         n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239,
         n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247,
         n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255,
         n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263,
         n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271,
         n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279,
         n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
         n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
         n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303,
         n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311,
         n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319,
         n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327,
         n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335,
         n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343,
         n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351,
         n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359,
         n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
         n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375,
         n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383,
         n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391,
         n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399,
         n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407,
         n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415,
         n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423,
         n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431,
         n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
         n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447,
         n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455,
         n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463,
         n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471,
         n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479,
         n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487,
         n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
         n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503,
         n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
         n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519,
         n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527,
         n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535,
         n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543,
         n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551,
         n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559,
         n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
         n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575,
         n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
         n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591,
         n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599,
         n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607,
         n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615,
         n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623,
         n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631,
         n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639,
         n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647,
         n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
         n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663,
         n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671,
         n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679,
         n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687,
         n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695,
         n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703,
         n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711,
         n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
         n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
         n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735,
         n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743,
         n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751,
         n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759,
         n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767,
         n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775,
         n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783,
         n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791,
         n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
         n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807,
         n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815,
         n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823,
         n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831,
         n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839,
         n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847,
         n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855,
         n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863,
         n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
         n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879,
         n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887,
         n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895,
         n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903,
         n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911,
         n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919,
         n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927,
         n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935,
         n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
         n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951,
         n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959,
         n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999,
         n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007,
         n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015,
         n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023,
         n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031,
         n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039,
         n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047,
         n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055,
         n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063,
         n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071,
         n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079,
         n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
         n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095,
         n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103,
         n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111,
         n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119,
         n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127,
         n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135,
         n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143,
         n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151,
         n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159,
         n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167,
         n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175,
         n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183,
         n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191,
         n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199,
         n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207,
         n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215,
         n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223,
         n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231,
         n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239,
         n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247,
         n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255,
         n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263,
         n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271,
         n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279,
         n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287,
         n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295,
         n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303,
         n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311,
         n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319,
         n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327,
         n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335,
         n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343,
         n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351,
         n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359,
         n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367,
         n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
         n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383,
         n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391,
         n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399,
         n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407,
         n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415,
         n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423,
         n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431,
         n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439,
         n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
         n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455,
         n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463,
         n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471,
         n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479,
         n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487,
         n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495,
         n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503,
         n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511,
         n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519,
         n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527,
         n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535,
         n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543,
         n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551,
         n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559,
         n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567,
         n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575,
         n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583,
         n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591,
         n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599,
         n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607,
         n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615,
         n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623,
         n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631,
         n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639,
         n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647,
         n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655,
         n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
         n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671,
         n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679,
         n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687,
         n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695,
         n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703,
         n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711,
         n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719,
         n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727,
         n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
         n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743,
         n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751,
         n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759,
         n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767,
         n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775,
         n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783,
         n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791,
         n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799,
         n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807,
         n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815,
         n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823,
         n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831,
         n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839,
         n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847,
         n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
         n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863,
         n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871,
         n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879,
         n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887,
         n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895,
         n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903,
         n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
         n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919,
         n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927,
         n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935,
         n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943,
         n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951,
         n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959,
         n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967,
         n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975,
         n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983,
         n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991,
         n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999,
         n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007,
         n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015,
         n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
         n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031,
         n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039,
         n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047,
         n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055,
         n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063,
         n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071,
         n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
         n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087,
         n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095,
         n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103,
         n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111,
         n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119,
         n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127,
         n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
         n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143,
         n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151,
         n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159,
         n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167,
         n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175,
         n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183,
         n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
         n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199,
         n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207,
         n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215,
         n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223,
         n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231,
         n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239,
         n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
         n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255,
         n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263,
         n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271,
         n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279,
         n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287,
         n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295,
         n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303,
         n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311,
         n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319,
         n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327,
         n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
         n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343,
         n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351,
         n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359,
         n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367,
         n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375,
         n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383,
         n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
         n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399,
         n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407,
         n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415,
         n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423,
         n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431,
         n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439,
         n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447,
         n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455,
         n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463,
         n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471,
         n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479,
         n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487,
         n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495,
         n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503,
         n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511,
         n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519,
         n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527,
         n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535,
         n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543,
         n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551,
         n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559,
         n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567,
         n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575,
         n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583,
         n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591,
         n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599,
         n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
         n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615,
         n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623,
         n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631,
         n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639,
         n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647,
         n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655,
         n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663,
         n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671,
         n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679,
         n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687,
         n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695,
         n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703,
         n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711,
         n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719,
         n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727,
         n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735,
         n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743,
         n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751,
         n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759,
         n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767,
         n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775,
         n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783,
         n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791,
         n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799,
         n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807,
         n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815,
         n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823,
         n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831,
         n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839,
         n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847,
         n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855,
         n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
         n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871,
         n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879,
         n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887,
         n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895,
         n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903,
         n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911,
         n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919,
         n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927,
         n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
         n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943,
         n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951,
         n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959,
         n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967,
         n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975,
         n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983,
         n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991,
         n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999,
         n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
         n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
         n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023,
         n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031,
         n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039,
         n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047,
         n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055,
         n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063,
         n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071,
         n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
         n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087,
         n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095,
         n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103,
         n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111,
         n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119,
         n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127,
         n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135,
         n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143,
         n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
         n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159,
         n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167,
         n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175,
         n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183,
         n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191,
         n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199,
         n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207,
         n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215,
         n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
         n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231,
         n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239,
         n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247,
         n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255,
         n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263,
         n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271,
         n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279,
         n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287,
         n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
         n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303,
         n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311,
         n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319,
         n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327,
         n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335,
         n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343,
         n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351,
         n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359,
         n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
         n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375,
         n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383,
         n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391,
         n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399,
         n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407,
         n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415,
         n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423,
         n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431,
         n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
         n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447,
         n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455,
         n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463,
         n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471,
         n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479,
         n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487,
         n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495,
         n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503,
         n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511,
         n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519,
         n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527,
         n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535,
         n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543,
         n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551,
         n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559,
         n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567,
         n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575,
         n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583,
         n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591,
         n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599,
         n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607,
         n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615,
         n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623,
         n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631,
         n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639,
         n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647,
         n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655,
         n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663,
         n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671,
         n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679,
         n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687,
         n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695,
         n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703,
         n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711,
         n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719,
         n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727,
         n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735,
         n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743,
         n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751,
         n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759,
         n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767,
         n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775,
         n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783,
         n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791,
         n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
         n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807,
         n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815,
         n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823,
         n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831,
         n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839,
         n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847,
         n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855,
         n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863,
         n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871,
         n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879,
         n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887,
         n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895,
         n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903,
         n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911,
         n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919,
         n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927,
         n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935,
         n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943,
         n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951,
         n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959,
         n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967,
         n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975,
         n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983,
         n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991,
         n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999,
         n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007,
         n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
         n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023,
         n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031,
         n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039,
         n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047,
         n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055,
         n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063,
         n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071,
         n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079,
         n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
         n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095,
         n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103,
         n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111,
         n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119,
         n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127,
         n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135,
         n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143,
         n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151,
         n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
         n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167,
         n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175,
         n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183,
         n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191,
         n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199,
         n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207,
         n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215,
         n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223,
         n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
         n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239,
         n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247,
         n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255,
         n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263,
         n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271,
         n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279,
         n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287,
         n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295,
         n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303,
         n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311,
         n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319,
         n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327,
         n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335,
         n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343,
         n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351,
         n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359,
         n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367,
         n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375,
         n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383,
         n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391,
         n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399,
         n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407,
         n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415,
         n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423,
         n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431,
         n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439,
         n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447,
         n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455,
         n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463,
         n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471,
         n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479,
         n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487,
         n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
         n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503,
         n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511,
         n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519,
         n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527,
         n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535,
         n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543,
         n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551,
         n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559,
         n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567,
         n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575,
         n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583,
         n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591,
         n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599,
         n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607,
         n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615,
         n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623,
         n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631,
         n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639,
         n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647,
         n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655,
         n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663,
         n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671,
         n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679,
         n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687,
         n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695,
         n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703,
         n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711,
         n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719,
         n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727,
         n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735,
         n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743,
         n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751,
         n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759,
         n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767,
         n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775,
         n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783,
         n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791,
         n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799,
         n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807,
         n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815,
         n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823,
         n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831,
         n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839,
         n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847,
         n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
         n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863,
         n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871,
         n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879,
         n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887,
         n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895,
         n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903,
         n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911,
         n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919,
         n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927,
         n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935,
         n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943,
         n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951,
         n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959,
         n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967,
         n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975,
         n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983,
         n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991,
         n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999,
         n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007,
         n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015,
         n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023,
         n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031,
         n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039,
         n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047,
         n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055,
         n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063,
         n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071,
         n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
         n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087,
         n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095,
         n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103,
         n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111,
         n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119,
         n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127,
         n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135,
         n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143,
         n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151,
         n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159,
         n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167,
         n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175,
         n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183,
         n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191,
         n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199,
         n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207,
         n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215,
         n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223,
         n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231,
         n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239,
         n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247,
         n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255,
         n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263,
         n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271,
         n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279,
         n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287,
         n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295,
         n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303,
         n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311,
         n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319,
         n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327,
         n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335,
         n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343,
         n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351,
         n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359,
         n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367,
         n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375,
         n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383,
         n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391,
         n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399,
         n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407,
         n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415,
         n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423,
         n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431,
         n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439,
         n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447,
         n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455,
         n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463,
         n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471,
         n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479,
         n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487,
         n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495,
         n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503,
         n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511,
         n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519,
         n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527,
         n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535,
         n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543,
         n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551,
         n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559,
         n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567,
         n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575,
         n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583,
         n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591,
         n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599,
         n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607,
         n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615,
         n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623,
         n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631,
         n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639,
         n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647,
         n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655,
         n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663,
         n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671,
         n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679,
         n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687,
         n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695,
         n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703,
         n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711,
         n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719,
         n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727,
         n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735,
         n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743,
         n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751,
         n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759,
         n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767,
         n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775,
         n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783,
         n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791,
         n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799,
         n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807,
         n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815,
         n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823,
         n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831,
         n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839,
         n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847,
         n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855,
         n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863,
         n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871,
         n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879,
         n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887,
         n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895,
         n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903,
         n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911,
         n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919,
         n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927,
         n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935,
         n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943,
         n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951,
         n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959,
         n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967,
         n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975,
         n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983,
         n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991,
         n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999,
         n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007,
         n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015,
         n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023,
         n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031,
         n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039,
         n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047,
         n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055,
         n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063,
         n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071,
         n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079,
         n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087,
         n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095,
         n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103,
         n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111,
         n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119,
         n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127,
         n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135,
         n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143,
         n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151,
         n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159,
         n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167,
         n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175,
         n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183,
         n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191,
         n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199,
         n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207,
         n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215,
         n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223,
         n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231,
         n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239,
         n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247,
         n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255,
         n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263,
         n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271,
         n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
         n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287,
         n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295,
         n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303,
         n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311,
         n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319,
         n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327,
         n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335,
         n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343,
         n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351,
         n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359,
         n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367,
         n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375,
         n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383,
         n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391,
         n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399,
         n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407,
         n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415,
         n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423,
         n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431,
         n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439,
         n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447,
         n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455,
         n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463,
         n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471,
         n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479,
         n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487,
         n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495,
         n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503,
         n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511,
         n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519,
         n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527,
         n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535,
         n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543,
         n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551,
         n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559,
         n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567,
         n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575,
         n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583,
         n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591,
         n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599,
         n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607,
         n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615,
         n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623,
         n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631,
         n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639,
         n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647,
         n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655,
         n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663,
         n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671,
         n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679,
         n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687,
         n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695,
         n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703,
         n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711,
         n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719,
         n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727,
         n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735,
         n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743,
         n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751,
         n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759,
         n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767,
         n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775,
         n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783,
         n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791,
         n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799,
         n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807,
         n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815,
         n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823,
         n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831,
         n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839,
         n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847,
         n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855,
         n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863,
         n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871,
         n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879,
         n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887,
         n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895,
         n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903,
         n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911,
         n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919,
         n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927,
         n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935,
         n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
         n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951,
         n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959,
         n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967,
         n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975,
         n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983,
         n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
         n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999,
         n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007,
         n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015,
         n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023,
         n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031,
         n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039,
         n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047,
         n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055,
         n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063,
         n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071,
         n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079,
         n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087,
         n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095,
         n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103,
         n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111,
         n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119,
         n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127,
         n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135,
         n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143,
         n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151,
         n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159,
         n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167,
         n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175,
         n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
         n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191,
         n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199,
         n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207,
         n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215,
         n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223,
         n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
         n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239,
         n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247,
         n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255,
         n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263,
         n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271,
         n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279,
         n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287,
         n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295,
         n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303,
         n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311,
         n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319,
         n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327,
         n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335,
         n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343,
         n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351,
         n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359,
         n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367,
         n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375,
         n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383,
         n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391,
         n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399,
         n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407,
         n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415,
         n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423,
         n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431,
         n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439,
         n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
         n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455,
         n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463,
         n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471,
         n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479,
         n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487,
         n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495,
         n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503,
         n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511,
         n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519,
         n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527,
         n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535,
         n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543,
         n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551,
         n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559,
         n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567,
         n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575,
         n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583,
         n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591,
         n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599,
         n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607,
         n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615,
         n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623,
         n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631,
         n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639,
         n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647,
         n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655,
         n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663,
         n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671,
         n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679,
         n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687,
         n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695,
         n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703,
         n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711,
         n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719,
         n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727,
         n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735,
         n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743,
         n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751,
         n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759,
         n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767,
         n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775,
         n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783,
         n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791,
         n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799,
         n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807,
         n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815,
         n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823,
         n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831,
         n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839,
         n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847,
         n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855,
         n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863,
         n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871,
         n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879,
         n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887,
         n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895,
         n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903,
         n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911,
         n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919,
         n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927,
         n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935,
         n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943,
         n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951,
         n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959,
         n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967,
         n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975,
         n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983,
         n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991,
         n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
         n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007,
         n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015,
         n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023,
         n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031,
         n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039,
         n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
         n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055,
         n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063,
         n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071,
         n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079,
         n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087,
         n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095,
         n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103,
         n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111,
         n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119,
         n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127,
         n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135,
         n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143,
         n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151,
         n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159,
         n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167,
         n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175,
         n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183,
         n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191,
         n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199,
         n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207,
         n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215,
         n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223,
         n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231,
         n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239,
         n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247,
         n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255,
         n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263,
         n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271,
         n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279,
         n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287,
         n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
         n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303,
         n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311,
         n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319,
         n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327,
         n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335,
         n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343,
         n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351,
         n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359,
         n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367,
         n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375,
         n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383,
         n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391,
         n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399,
         n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407,
         n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415,
         n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423,
         n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431,
         n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439,
         n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447,
         n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455,
         n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463,
         n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471,
         n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479,
         n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487,
         n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495,
         n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503,
         n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511,
         n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519,
         n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527,
         n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
         n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543,
         n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551,
         n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559,
         n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567,
         n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575,
         n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583,
         n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591,
         n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599,
         n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607,
         n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615,
         n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623,
         n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631,
         n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639,
         n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647,
         n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655,
         n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663,
         n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671,
         n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679,
         n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687,
         n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695,
         n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703,
         n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711,
         n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719,
         n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727,
         n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735,
         n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743,
         n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
         n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759,
         n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767,
         n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775,
         n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783,
         n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791,
         n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799,
         n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807,
         n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815,
         n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823,
         n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831,
         n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839,
         n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847,
         n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855,
         n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863,
         n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871,
         n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879,
         n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887,
         n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895,
         n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903,
         n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911,
         n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919,
         n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927,
         n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935,
         n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943,
         n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951,
         n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959,
         n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967,
         n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975,
         n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983,
         n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991,
         n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999,
         n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007,
         n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015,
         n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023,
         n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031,
         n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039,
         n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047,
         n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055,
         n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063,
         n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071,
         n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079,
         n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087,
         n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095,
         n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103,
         n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111,
         n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119,
         n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127,
         n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135,
         n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143,
         n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151,
         n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159,
         n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167,
         n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175,
         n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183,
         n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191,
         n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199,
         n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207,
         n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215,
         n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223,
         n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231,
         n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239,
         n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247,
         n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255,
         n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263,
         n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271,
         n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279,
         n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287,
         n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295,
         n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303,
         n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311,
         n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319,
         n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327,
         n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335,
         n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343,
         n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351,
         n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359,
         n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367,
         n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375,
         n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383,
         n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391,
         n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399,
         n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407,
         n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415,
         n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423,
         n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431,
         n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439,
         n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447,
         n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455,
         n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463,
         n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471,
         n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479,
         n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487,
         n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495,
         n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503,
         n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511,
         n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519,
         n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527,
         n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535,
         n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543,
         n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551,
         n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559,
         n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567,
         n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575,
         n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583,
         n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591,
         n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599,
         n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607,
         n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615,
         n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623,
         n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631,
         n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639,
         n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647,
         n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655,
         n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663,
         n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671,
         n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679,
         n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687,
         n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695,
         n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703,
         n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711,
         n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719,
         n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727,
         n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
         n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743,
         n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751,
         n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759,
         n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767,
         n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775,
         n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783,
         n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791,
         n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799,
         n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807,
         n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815,
         n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823,
         n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831,
         n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839,
         n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847,
         n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855,
         n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863,
         n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871,
         n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879,
         n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887,
         n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895,
         n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903,
         n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911,
         n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919,
         n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927,
         n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935,
         n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943,
         n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951,
         n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959,
         n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967,
         n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975,
         n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983,
         n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991,
         n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999,
         n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007,
         n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015,
         n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023,
         n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031,
         n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039,
         n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047,
         n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055,
         n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063,
         n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071,
         n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079,
         n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087,
         n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095,
         n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103,
         n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111,
         n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119,
         n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127,
         n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135,
         n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143,
         n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151,
         n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159,
         n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167,
         n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175,
         n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183,
         n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191,
         n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199,
         n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207,
         n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215,
         n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223,
         n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231,
         n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239,
         n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247,
         n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255,
         n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263,
         n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271,
         n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279,
         n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287,
         n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295,
         n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303,
         n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311,
         n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319,
         n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327,
         n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335,
         n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343,
         n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351,
         n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359,
         n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367,
         n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375,
         n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383,
         n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391,
         n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399,
         n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407,
         n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415,
         n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423,
         n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431,
         n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439,
         n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447,
         n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455,
         n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463,
         n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471,
         n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479,
         n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487,
         n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495,
         n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503,
         n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511,
         n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519,
         n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527,
         n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535,
         n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543,
         n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551,
         n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559,
         n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567,
         n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575,
         n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583,
         n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591,
         n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
         n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607,
         n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615,
         n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623,
         n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631,
         n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639,
         n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647,
         n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655,
         n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663,
         n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671,
         n41672;
  or U22375(G1730,G59806,G59807,n34802,n34803);
  or U22376(n20960,n34701,n20962);
  nor U22377(n21952,n21950,G59428);
  nor U22378(n28778,n28776,G58979);
  nor U22379(n35797,n35795,G59877);
  nand U22380(n22401,n21044,n22456);
  nand U22381(n29192,n27929,n29247);
  nand U22382(n36233,n34898,n36288);
  nor U22383(n34701,n34795,n20962);
  nor U22384(n22056,n21057,n22055);
  nor U22385(n28882,n27942,n28881);
  nor U22386(n35901,n34911,n35900);
  nor U22387(n27745,n20965,G59390);
  nor U22388(n34464,n27851,G58941);
  nor U22389(n41570,n34820,G59839);
  not U22390(n20961,n20960);
  not U22391(n20962,G1730);
  not U22392(n22414,n22406);
  nor U22393(n22406,n25487,n22163,n21080);
  not U22394(n29205,n29197);
  nor U22395(n29197,n32281,n28959,n27965);
  not U22396(n36246,n36238);
  nor U22397(n36238,n39320,n35994,n34934);
  nor U22398(n34045,n29349,n29226,n28877);
  nand U22399(n30513,n29349,n30514);
  nand U22400(n30437,n29349,n30434);
  nand U22401(n30363,n29349,n30360);
  nand U22402(n30274,n29349,n30275);
  nand U22403(n30190,n29349,n30191);
  nor U22404(n41151,n36390,n36267,n35896);
  nand U22405(n37553,n36390,n37554);
  nand U22406(n37477,n36390,n37474);
  nand U22407(n37403,n36390,n37400);
  nand U22408(n37314,n36390,n37315);
  nand U22409(n37230,n36390,n37231);
  nor U22410(n27325,n22567,n22435,n22051);
  nand U22411(n23719,n22567,n23720);
  nand U22412(n23643,n22567,n23640);
  nand U22413(n23561,n22567,n23558);
  nand U22414(n23472,n22567,n23473);
  nand U22415(n23388,n22567,n23389);
  nor U22416(n28973,n27932,n29047);
  nor U22417(n22177,n21047,n22257);
  nor U22418(n36008,n34901,n36089);
  nor U22419(n28594,n28761,n28581);
  nor U22420(n21714,n21935,n21700);
  nor U22421(n35567,n35781,n35554);
  nor U22422(n28456,n28573,n28452);
  nor U22423(n21571,n21688,n21567);
  nor U22424(n35425,n35542,n35421);
  nor U22425(n28576,n32285,n28416);
  nor U22426(n35545,n39324,n35385);
  nor U22427(n21691,n25491,n21531);
  and U22428(n29194,n32147,n32282);
  and U22429(n22403,n25353,n25488);
  and U22430(n36235,n39186,n39321);
  and U22431(n28881,n28762,n28960);
  and U22432(n22055,n21936,n22164);
  and U22433(n35900,n35782,n35995);
  nor U22434(n34473,n34466,n27851);
  nor U22435(n27755,n27748,n20965);
  nor U22436(n41579,n41572,n34820);
  nor U22437(n28972,n28416,n29047);
  nor U22438(n22176,n21531,n22257);
  nor U22439(n36007,n35385,n36089);
  nor U22440(n28451,n28572,n28452);
  nor U22441(n21566,n21687,n21567);
  nor U22442(n35420,n35541,n35421);
  nor U22443(n29264,n28689,n28573);
  nor U22444(n36305,n35692,n35542);
  nor U22445(n22473,n21846,n21688);
  nand U22446(n29287,n33969,n33904,n33970);
  nand U22447(n36328,n41075,n41010,n41076);
  nand U22448(n22496,n27249,n27184,n27250);
  nand U22449(n32013,n29231,n27900);
  nand U22450(n31897,n29231,n27891);
  nand U22451(n31767,n29231,n27881);
  nand U22452(n31654,n29231,n27871);
  nand U22453(n31516,n29231,n28360);
  nand U22454(n39052,n36272,n34869);
  nand U22455(n38937,n36272,n34860);
  nand U22456(n38807,n36272,n34850);
  nand U22457(n38693,n36272,n34840);
  nand U22458(n38555,n36272,n35329);
  nand U22459(n25219,n22440,n21015);
  nand U22460(n25104,n22440,n21006);
  nand U22461(n24974,n22440,n20996);
  nand U22462(n24861,n22440,n20986);
  nand U22463(n24722,n22440,n21475);
  not U22464(n34570,n34569);
  nand U22465(n34569,n34629,n34630,n34631);
  not U22466(n28776,n28771);
  not U22467(n21950,n21945);
  not U22468(n35795,n35791);
  and U22469(n28452,n28574,n28575);
  nand U22470(n28575,n27870,n27965,n28576);
  and U22471(n21567,n21689,n21690);
  nand U22472(n21690,n20985,n21080,n21691);
  and U22473(n35421,n35543,n35544);
  nand U22474(n35544,n34839,n34934,n35545);
  not U22475(n21700,n21847);
  not U22476(n35554,n35693);
  nor U22477(n28331,n28205,n28332,n28333,n28334);
  nor U22478(n28321,n28205,n28322,n28323,n28324);
  nor U22479(n28311,n28205,n28312,n28313,n28314);
  nor U22480(n21446,n21320,n21447,n21448,n21449);
  nor U22481(n21436,n21320,n21437,n21438,n21439);
  nor U22482(n21426,n21320,n21427,n21428,n21429);
  nor U22483(n35300,n35174,n35301,n35302,n35303);
  nor U22484(n35290,n35174,n35291,n35292,n35293);
  nor U22485(n35280,n35174,n35281,n35282,n35283);
  not U22486(n28581,n28690);
  nand U22487(n28690,n28762,n28763);
  not U22488(n27943,n28689);
  nand U22489(n28689,n34366,n34367,n34368,n34369);
  not U22490(n21058,n21846);
  nand U22491(n21846,n27646,n27647,n27648,n27649);
  not U22492(n34805,n35621);
  not U22493(n34912,n35692);
  nand U22494(n35692,n41472,n41473,n41474,n41475);
  not U22495(n27851,n27852);
  not U22496(n20965,n20966);
  not U22497(n34820,n34821);
  nor U22498(n28974,n29047,n29173);
  nor U22499(n22178,n22257,n22382);
  nor U22500(n36009,n36089,n36214);
  not U22501(G1731,n34635);
  nor U22502(n34635,n34801,G59360);
  nor U22503(n29261,n32031,n32161,n32162);
  nor U22504(n32161,n27943,n32310);
  nor U22505(n22470,n25237,n25367,n25368);
  nor U22506(n25367,n21058,n25516);
  nor U22507(n36302,n39070,n39200,n39201);
  nor U22508(n39200,n34912,n39349);
  nand U22509(n21776,G59360,n34806);
  nand U22510(n34806,n34807,n34808,n34809,n34810);
  not U22511(n28963,n27993);
  nor U22512(n27993,n32286,n28416);
  nor U22513(n32417,n33639,n32332);
  not U22514(n32332,n32428);
  nor U22515(n25623,n26919,n25538);
  not U22516(n25538,n25634);
  nor U22517(n39456,n40745,n39371);
  not U22518(n39371,n39467);
  not U22519(n22167,n21108);
  nor U22520(n21108,n25492,n21531);
  not U22521(n36215,n36267);
  nor U22522(n36267,n40749,G60246);
  not U22523(n29174,n29226);
  nor U22524(n29226,n33643,G59348);
  not U22525(n35998,n34962);
  nor U22526(n34962,n39325,n35385);
  not U22527(n22383,n22435);
  nor U22528(n22435,n26923,G59797);
  nand U22529(G9273,n20963,n20964);
  nand U22530(n20964,G59356,n20965);
  nand U22531(n20963,G59790,n20966);
  nand U22532(G9272,n20967,n20968);
  nand U22533(n20968,G59357,n20965);
  nand U22534(n20967,G59791,n20966);
  nand U22535(G9271,n20969,n20970);
  nand U22536(n20970,G59358,n20965);
  nand U22537(n20969,G59792,n20966);
  nand U22538(G9270,n20971,n20972);
  nand U22539(n20972,G59359,n20965);
  nand U22540(n20971,G59793,n20966);
  nand U22541(G9269,n20973,n20974);
  nand U22542(n20974,n20975,n20976,n20977);
  nand U22543(n20973,G59393,n20978);
  nand U22544(G9268,n20979,n20980);
  nand U22545(n20980,G59394,n20978);
  nand U22546(n20979,n20981,n20977);
  nand U22547(n20981,n20976,n20975);
  not U22548(n20975,n20982);
  nand U22549(G9267,n20983,n20984);
  nand U22550(n20984,n20985,n20986,n20987,n20988);
  nand U22551(n20983,n20989,G59557);
  nand U22552(G9266,n20990,n20991);
  nand U22553(n20991,n20989,G59558);
  nand U22554(n20990,n20992,n20988);
  nand U22555(n20992,n20993,n20994);
  nand U22556(n20994,n20995,n20996);
  nand U22557(n20993,n20985,n20997);
  nand U22558(G9265,n20998,n20999);
  nand U22559(n20999,n20989,G59559);
  nand U22560(n20998,n21000,n20988);
  nand U22561(n21000,n21001,n21002,n21003);
  nand U22562(n21003,n20985,n21004);
  nand U22563(n21002,G59427,n21005,G59567);
  nand U22564(n21001,n21006,n20995);
  nand U22565(G9263,n21007,n21008);
  nand U22566(n21008,n20989,G59560);
  nand U22567(n21007,n21009,n20988);
  nand U22568(n21009,n21010,n21011,n21012);
  nand U22569(n21012,n20985,n21013);
  nand U22570(n21011,G59427,n21014,G59567);
  nand U22571(n21010,n21015,n20995);
  nand U22572(G9262,n21016,n21017);
  nand U22573(n21017,n20989,G59561);
  not U22574(n20989,n20988);
  nand U22575(n21016,n21018,n20988);
  nand U22576(n20988,n21019,n21020,n21021);
  nand U22577(n21021,n21022,n21023);
  nand U22578(n21018,n21024,n21025,n21026);
  nand U22579(n21026,n20985,n21027);
  nand U22580(n21025,G59427,n21028);
  nand U22581(n21028,G59567,n21029);
  nand U22582(n21024,n20995,n21030);
  nor U22583(n20995,n21031,G59426);
  nand U22584(G9261,n21032,n21033);
  or U22585(n21033,n20965,G59803);
  nand U22586(n21032,G59794,n20965);
  nand U22587(G9260,n21034,n21035);
  or U22588(n21035,n21036,n21037);
  nand U22589(n21034,n21038,n21036);
  nand U22590(n21036,n21039,n21040,n21041,n21042);
  nand U22591(n21041,n21043,n21044);
  nand U22592(n21040,G59427,n21045,n21046);
  nand U22593(n21038,n21047,n21048);
  nand U22594(n21048,G59428,n21049);
  nand U22595(n21049,n21050,n21045);
  nand U22596(n21050,n21051,n21052);
  nand U22597(n21052,G59426,n21053);
  nand U22598(n21053,n21054,n21055);
  nand U22599(n21055,n21056,n21057);
  nand U22600(n21056,n21058,n21059);
  nand U22601(n21054,G59797,n21060);
  nand U22602(n21051,n21061,n21058);
  nand U22603(G9259,n21062,n21063);
  nand U22604(n21063,G59800,n20965);
  nand U22605(n21062,G59804,n20966);
  nand U22606(G9258,n21064,n21065);
  nand U22607(n21065,n21066,G59803);
  nand U22608(n21064,n21067,n21068);
  nand U22609(n21067,n21069,n21070,G59426);
  nand U22610(G9257,n21071,n21072);
  nand U22611(n21072,n21066,G59804);
  not U22612(n21066,n21068);
  nand U22613(n21071,n21068,n21073);
  nand U22614(n21068,n21039,n21074);
  nand U22615(n21074,n21075,n21043);
  nand U22616(G8744,n21076,n21077,n21078,n21079);
  nand U22617(n21079,G59428,n21080,n21081);
  nand U22618(n21078,n21082,G59566);
  nand U22619(n21077,n21083,n21084);
  nand U22620(n21076,n21085,n21086);
  nand U22621(G8742,n20978,n21087);
  nand U22622(n21087,G59802,G59392);
  nand U22623(G8741,n21088,n21089);
  nand U22624(n21089,G59428,n21043,n21075);
  nand U22625(n21088,G59801,n21090);
  nand U22626(n21090,n21091,n21022);
  nand U22627(G8740,n21092,n21093,n21094);
  or U22628(n21093,n20965,G59801);
  nand U22629(n21092,G59799,n20965);
  nand U22630(G8739,n21095,n21096,n21094);
  nand U22631(n21094,n20982,n21097);
  nand U22632(n21096,G35,n20977);
  nand U22633(n21095,G59797,n20978);
  nand U22634(G8738,n21098,n21099);
  nand U22635(n21099,n21100,n21101);
  nand U22636(n21100,n21102,n21103);
  nand U22637(n21103,n21104,n21105);
  nand U22638(n21104,n21106,n21107);
  nand U22639(n21107,n21108,n20985);
  nand U22640(n21102,n21031,n21109);
  nand U22641(n21109,n21110,n21111);
  nand U22642(n21111,n20985,n21112);
  nand U22643(n21112,n21113,n21114);
  nand U22644(n21098,G59796,n21115);
  nand U22645(G8737,n21116,n21117);
  nand U22646(n21117,G59795,n21115);
  nand U22647(n21115,n21022,n21101);
  nand U22648(G8736,n21118,n21119,n21120);
  nand U22649(n21119,G59793,n21121);
  or U22650(n21118,n21121,n21122);
  nand U22651(G8735,n21120,n21123,n21124);
  nand U22652(n21124,G59792,n21121);
  not U22653(n21120,n21125);
  nand U22654(G8734,n21126,n21127,n21128);
  nand U22655(n21128,G59791,n21121);
  nand U22656(n21127,n21129,n21130,n21131);
  nand U22657(n21129,G59758,G59393);
  nand U22658(n21126,n21125,G59758);
  nor U22659(n21125,n21121,n21130);
  nand U22660(G8733,n21132,n21123,n21133);
  nand U22661(n21133,G59790,n21121);
  nand U22662(n21123,n21134,n21122,n21131);
  not U22663(n21134,G59393);
  nand U22664(n21132,n21131,n21130);
  nor U22665(n21131,n21121,G59394);
  nand U22666(n21121,n21135,n21136,n21137,n21138);
  nor U22667(n21138,n21139,n21140,n21141,n21142);
  nand U22668(n21142,n21143,n21144,n21145,n21146);
  nand U22669(n21141,n21147,n21148,n21149,n21150);
  nand U22670(n21140,n21151,n21152,n21153,n21154);
  nand U22671(n21139,n21155,n21156,n21157,n21158);
  nor U22672(n21137,n21159,n21160,G59396,G59395);
  and U22673(n21160,G59393,G59394);
  nand U22674(n21159,n21161,n21162,n21163,n21164);
  nor U22675(n21136,G59408,G59407,G59406,G59405);
  nor U22676(n21135,G59404,G59403,G59402,G59401);
  nand U22677(G8732,n21165,n21166,n21167,n21168);
  nor U22678(n21168,n21169,n21170,n21171);
  nor U22679(n21171,n21172,n21173);
  and U22680(n21170,n21174,n21175);
  nor U22681(n21169,n21176,n21177);
  nand U22682(n21167,n21178,n21179);
  nand U22683(n21166,n21180,n21181);
  nand U22684(n21165,n21182,G59757);
  nand U22685(G8731,n21183,n21184,n21185,n21186);
  nor U22686(n21186,n21187,n21188,n21189);
  nor U22687(n21189,n21190,n21173);
  nor U22688(n21188,n21191,n21192);
  nor U22689(n21187,n21193,n21177);
  nand U22690(n21185,n21194,n21179);
  nand U22691(n21184,n21180,n21195);
  nand U22692(n21183,n21182,G59756);
  nand U22693(G8730,n21196,n21197,n21198,n21199);
  nor U22694(n21199,n21200,n21201,n21202);
  nor U22695(n21202,n21203,n21173);
  nor U22696(n21201,n21191,n21204);
  nor U22697(n21200,n21205,n21177);
  nand U22698(n21198,n21206,n21179);
  nand U22699(n21197,n21207,n21180);
  nand U22700(n21196,n21182,G59755);
  nand U22701(G8729,n21208,n21209,n21210,n21211);
  nor U22702(n21211,n21212,n21213,n21214);
  nor U22703(n21214,n21215,n21173);
  nor U22704(n21213,n21191,n21216);
  nor U22705(n21212,n21217,n21177);
  nand U22706(n21210,n21218,n21179);
  nand U22707(n21209,n21180,n21219);
  nand U22708(n21208,n21182,G59754);
  nand U22709(G8728,n21220,n21221,n21222,n21223);
  nor U22710(n21223,n21224,n21225,n21226);
  nor U22711(n21226,n21227,n21173);
  nor U22712(n21225,n21191,n21228);
  nor U22713(n21224,n21229,n21177);
  nand U22714(n21222,n21230,n21179);
  nand U22715(n21221,n21180,n21231);
  nand U22716(n21220,n21182,G59753);
  nand U22717(G8727,n21232,n21233,n21234,n21235);
  nor U22718(n21235,n21236,n21237,n21238);
  nor U22719(n21238,n21239,n21173);
  nor U22720(n21237,n21191,n21240);
  nor U22721(n21236,n21241,n21177);
  nand U22722(n21234,n21242,n21179);
  nand U22723(n21233,n21180,n21243);
  nand U22724(n21232,n21182,G59752);
  nand U22725(G8726,n21244,n21245,n21246,n21247);
  nor U22726(n21247,n21248,n21249,n21250);
  nor U22727(n21250,n21251,n21173);
  and U22728(n21249,n21174,n21252);
  nor U22729(n21248,n21253,n21177);
  nand U22730(n21246,n21254,n21179);
  nand U22731(n21245,n21180,n21255);
  nand U22732(n21244,n21182,G59751);
  nand U22733(G8725,n21256,n21257,n21258,n21259);
  nor U22734(n21259,n21260,n21261,n21262);
  nor U22735(n21262,n21263,n21173);
  nor U22736(n21261,n21191,n21264);
  nor U22737(n21260,n21265,n21177);
  nand U22738(n21258,n21266,n21179);
  nand U22739(n21257,n21180,n21267);
  nand U22740(n21256,n21182,G59750);
  nand U22741(G8724,n21268,n21269,n21270,n21271);
  nor U22742(n21271,n21272,n21273,n21274);
  nor U22743(n21274,n21275,n21173);
  nor U22744(n21273,n21191,n21276);
  nor U22745(n21272,n21277,n21177);
  nand U22746(n21270,n21278,n21179);
  nand U22747(n21269,n21180,n21279);
  nand U22748(n21268,n21182,G59749);
  nand U22749(G8723,n21280,n21281,n21282,n21283);
  nor U22750(n21283,n21284,n21285,n21286);
  nor U22751(n21286,n21287,n21173);
  and U22752(n21285,n21174,n21288);
  nor U22753(n21284,n21289,n21177);
  nand U22754(n21282,n21290,n21179);
  nand U22755(n21281,n21180,n21291);
  nand U22756(n21280,n21182,G59748);
  nand U22757(G8722,n21292,n21293,n21294,n21295);
  nor U22758(n21295,n21296,n21297,n21298);
  nor U22759(n21298,n21299,n21173);
  nor U22760(n21297,n21191,n21300);
  nor U22761(n21296,n21301,n21177);
  nand U22762(n21294,n21302,n21179);
  nand U22763(n21293,n21180,n21303);
  nand U22764(n21292,n21182,G59747);
  nand U22765(G8721,n21304,n21305,n21306,n21307);
  nor U22766(n21307,n21308,n21309,n21310);
  nor U22767(n21310,n21311,n21173);
  nor U22768(n21309,n21191,n21312);
  nor U22769(n21308,n21313,n21177);
  nand U22770(n21306,n21314,n21179);
  nand U22771(n21305,n21180,n21315);
  nand U22772(n21304,n21182,G59746);
  nand U22773(G8720,n21316,n21317,n21318,n21319);
  nor U22774(n21319,n21320,n21321,n21322,n21323);
  nor U22775(n21323,n21324,n21325);
  and U22776(n21322,G59745,n21182);
  and U22777(n21321,n21326,n21180);
  nand U22778(n21318,n21327,G59777);
  nand U22779(n21317,n21328,n21174);
  nand U22780(n21316,n21329,G59618);
  nand U22781(G8719,n21330,n21331,n21332,n21333);
  nor U22782(n21333,n21320,n21334,n21335,n21336);
  nor U22783(n21336,n21324,n21337);
  and U22784(n21335,G59744,n21182);
  and U22785(n21334,n21338,n21180);
  nand U22786(n21332,n21327,G59776);
  nand U22787(n21331,n21339,n21174);
  nand U22788(n21330,n21329,G59617);
  nand U22789(G8718,n21340,n21341,n21342,n21343);
  nor U22790(n21343,n21320,n21344,n21345,n21346);
  nor U22791(n21346,n21324,n21347);
  and U22792(n21345,G59743,n21182);
  and U22793(n21344,n21348,n21180);
  nand U22794(n21342,n21327,G59775);
  nand U22795(n21341,n21349,n21174);
  nand U22796(n21340,n21329,G59616);
  nand U22797(G8717,n21350,n21351,n21352,n21353);
  nor U22798(n21353,n21320,n21354,n21355,n21356);
  nor U22799(n21356,n21324,n21357);
  and U22800(n21355,G59742,n21182);
  and U22801(n21354,n21358,n21180);
  nand U22802(n21352,n21327,G59774);
  nand U22803(n21351,n21359,n21174);
  nand U22804(n21350,n21329,G59615);
  nand U22805(G8716,n21360,n21361,n21362,n21363);
  nor U22806(n21363,n21320,n21364,n21365,n21366);
  nor U22807(n21366,n21324,n21367);
  and U22808(n21365,G59741,n21182);
  and U22809(n21364,n21368,n21180);
  nand U22810(n21362,n21327,G59773);
  nand U22811(n21361,n21369,n21174);
  nand U22812(n21360,n21329,G59614);
  nand U22813(G8715,n21370,n21371,n21372,n21373);
  nor U22814(n21373,n21320,n21374,n21375,n21376);
  nor U22815(n21376,n21324,n21377);
  and U22816(n21375,G59740,n21182);
  and U22817(n21374,n21378,n21180);
  nand U22818(n21372,n21327,G59772);
  nand U22819(n21371,n21379,n21174);
  nand U22820(n21370,n21329,G59613);
  nand U22821(G8714,n21380,n21381,n21382,n21383);
  nor U22822(n21383,n21320,n21384,n21385,n21386);
  nor U22823(n21386,n21324,n21387);
  and U22824(n21385,G59739,n21182);
  and U22825(n21384,n21180,n21388);
  nand U22826(n21382,n21327,G59771);
  nand U22827(n21381,n21389,n21174);
  nand U22828(n21380,n21329,G59612);
  nand U22829(G8713,n21390,n21391,n21392,n21393);
  nor U22830(n21393,n21320,n21394,n21395,n21396);
  nor U22831(n21396,n21324,n21397);
  and U22832(n21395,G59738,n21182);
  and U22833(n21394,n21398,n21180);
  nand U22834(n21392,n21327,G59770);
  nand U22835(n21391,n21399,n21174);
  nand U22836(n21390,n21329,G59611);
  nand U22837(G8712,n21400,n21401,n21402,n21403);
  nor U22838(n21403,n21320,n21404,n21405,n21406);
  nor U22839(n21406,n21324,n21407);
  and U22840(n21405,G59737,n21182);
  and U22841(n21404,n21408,n21180);
  nand U22842(n21402,n21327,G59769);
  nand U22843(n21401,n21409,n21174);
  nand U22844(n21400,n21329,G59610);
  nand U22845(G8711,n21410,n21411,n21412,n21413);
  nor U22846(n21413,n21320,n21414,n21415,n21416);
  nor U22847(n21416,n21324,n21417);
  nor U22848(n21415,n21418,n21419);
  nor U22849(n21414,n21420,n21421);
  nand U22850(n21412,n21327,G59768);
  nand U22851(n21411,n21422,n21174);
  nand U22852(n21410,n21329,G59609);
  nand U22853(G8710,n21423,n21424,n21425,n21426);
  nor U22854(n21429,n21324,n21430);
  and U22855(n21428,G59735,n21182);
  and U22856(n21427,n21431,n21180);
  nand U22857(n21425,n21327,G59767);
  nand U22858(n21424,n21432,n21174);
  nand U22859(n21423,n21329,G59608);
  nand U22860(G8709,n21433,n21434,n21435,n21436);
  nor U22861(n21439,n21324,n21440);
  and U22862(n21438,G59734,n21182);
  and U22863(n21437,n21180,n21441);
  nand U22864(n21435,n21327,G59766);
  nand U22865(n21434,n21442,n21174);
  nand U22866(n21433,n21329,G59607);
  nand U22867(G8708,n21443,n21444,n21445,n21446);
  nor U22868(n21449,n21324,n21450);
  and U22869(n21448,G59733,n21182);
  and U22870(n21447,n21180,n21451);
  not U22871(n21180,n21420);
  nand U22872(n21445,n21327,G59765);
  nand U22873(n21444,n21452,n21174);
  nand U22874(n21443,n21329,G59606);
  nand U22875(G8707,n21453,n21454,n21455,n21456);
  nor U22876(n21456,n21320,n21457,n21458,n21459);
  nor U22877(n21459,n21324,n21460);
  nor U22878(n21458,n21461,n21419);
  nor U22879(n21457,n21420,n21462);
  nand U22880(n21455,n21327,G59764);
  nand U22881(n21454,n21463,n21174);
  nand U22882(n21453,n21329,G59605);
  nand U22883(G8706,n21464,n21465,n21466,n21467);
  nor U22884(n21467,n21320,n21468,n21469,n21470);
  nor U22885(n21470,n21324,n21471);
  nor U22886(n21469,n21472,n21419);
  and U22887(n21468,n21473,n21474);
  nand U22888(n21466,n21327,G59763);
  nand U22889(n21465,n21475,n21476);
  nand U22890(n21464,n21329,G59604);
  nand U22891(G8705,n21477,n21478,n21479,n21480);
  nor U22892(n21480,n21320,n21481,n21482,n21483);
  nor U22893(n21483,n21324,n21484);
  not U22894(n21324,n21179);
  nor U22895(n21482,n21485,n21419);
  and U22896(n21481,n21473,n21486);
  nor U22897(n21320,G59427,G59428,n21327);
  nand U22898(n21479,n21327,G59762);
  nand U22899(n21478,n20986,n21476);
  nand U22900(n21477,n21329,G59603);
  nand U22901(G8704,n21487,n21488,n21489,n21490);
  nor U22902(n21490,n21491,n21492,n21493);
  nor U22903(n21493,n21494,n21173);
  nor U22904(n21492,n21495,n21496);
  nor U22905(n21491,n21497,n21177);
  nand U22906(n21489,n21498,n21179);
  nand U22907(n21488,n21499,n21473);
  nand U22908(n21487,n21182,G59729);
  nand U22909(G8703,n21500,n21501,n21502,n21503);
  nor U22910(n21503,n21504,n21505,n21506);
  nor U22911(n21506,n21507,n21173);
  nor U22912(n21505,n21495,n21508);
  nor U22913(n21504,n21509,n21177);
  nand U22914(n21502,n21510,n21179);
  nand U22915(n21501,n21511,n21473);
  nand U22916(n21500,n21182,G59728);
  nand U22917(G8702,n21512,n21513,n21514,n21515);
  nor U22918(n21515,n21516,n21517,n21518);
  nor U22919(n21518,n21519,n21173);
  nor U22920(n21517,n21495,n21520);
  nor U22921(n21516,n21130,n21177);
  nand U22922(n21514,n21521,n21179);
  nand U22923(n21513,n21522,n21473);
  nand U22924(n21512,n21182,G59727);
  nand U22925(G8701,n21523,n21524,n21525,n21526);
  nor U22926(n21526,n21527,n21528,n21529);
  nor U22927(n21529,n21530,n21173);
  not U22928(n21173,n21329);
  nor U22929(n21329,n21327,G59426,n21531);
  nor U22930(n21528,n21495,n21532);
  not U22931(n21495,n21476);
  nand U22932(n21476,n21191,n21533);
  nand U22933(n21533,n21534,n21057,n21535);
  not U22934(n21191,n21174);
  nand U22935(n21174,n21536,n21537);
  nand U22936(n21537,n21178,n21177,G59427);
  nand U22937(n21536,n21538,n21539,n21535);
  nor U22938(n21527,n21122,n21177);
  nand U22939(n21525,n21084,n21179);
  nand U22940(n21179,n21540,n21541);
  nand U22941(n21541,n21535,n21539,n21542,n21543);
  not U22942(n21542,n21544);
  nand U22943(n21540,G59427,n21177,n21545);
  nand U22944(n21524,n21546,n21473);
  nand U22945(n21473,n21547,n21420);
  nand U22946(n21420,n21535,n21538,n21060,n21548);
  nand U22947(n21547,n21177,n21534,n21061);
  nand U22948(n21523,n21182,G59726);
  not U22949(n21182,n21419);
  nand U22950(n21419,n21535,n21549);
  nand U22951(n21549,n21550,n21551);
  nand U22952(n21551,n21544,n21543,n21539);
  not U22953(n21543,n21538);
  nand U22954(n21550,n21548,n21552);
  nand U22955(n21552,n21538,n21060);
  nor U22956(n21535,n21044,n21327);
  not U22957(n21327,n21177);
  nand U22958(n21177,n21039,n21553,n21554,n21555);
  nor U22959(n21039,n21556,n21557);
  nor U22960(n21557,n21110,n21031);
  nor U22961(n21110,n21558,n21559);
  nor U22962(n21559,n21560,n21044,n21561);
  nor U22963(n21558,n21562,n21563);
  nand U22964(G8700,n21564,n21565);
  nand U22965(n21565,n21566,n21178);
  nand U22966(n21564,n21567,G59757);
  nand U22967(G8699,n21568,n21569,n21570);
  nand U22968(n21570,n21567,G59756);
  nand U22969(n21569,n21566,n21194);
  nand U22970(n21568,n21571,n21572);
  nand U22971(G8698,n21573,n21574,n21575);
  nand U22972(n21575,n21567,G59755);
  nand U22973(n21574,n21566,n21206);
  nand U22974(n21573,n21571,n21576);
  nand U22975(G8697,n21577,n21578,n21579);
  nand U22976(n21579,n21567,G59754);
  nand U22977(n21578,n21566,n21218);
  nand U22978(n21577,n21571,n21580);
  nand U22979(G8696,n21581,n21582,n21583);
  nand U22980(n21583,n21567,G59753);
  nand U22981(n21582,n21566,n21230);
  nand U22982(n21581,n21571,n21584);
  nand U22983(G8695,n21585,n21586,n21587);
  nand U22984(n21587,n21567,G59752);
  nand U22985(n21586,n21566,n21242);
  nand U22986(n21585,n21571,n21588);
  nand U22987(G8694,n21589,n21590,n21591);
  nand U22988(n21591,n21567,G59751);
  nand U22989(n21590,n21566,n21254);
  nand U22990(n21589,n21571,n21252);
  nand U22991(G8693,n21592,n21593,n21594);
  nand U22992(n21594,n21567,G59750);
  nand U22993(n21593,n21566,n21266);
  nand U22994(n21592,n21571,n21595);
  nand U22995(G8692,n21596,n21597,n21598);
  nand U22996(n21598,n21567,G59749);
  nand U22997(n21597,n21566,n21278);
  nand U22998(n21596,n21571,n21599);
  nand U22999(G8691,n21600,n21601,n21602);
  nand U23000(n21602,n21567,G59748);
  nand U23001(n21601,n21566,n21290);
  nand U23002(n21600,n21571,n21288);
  nand U23003(G8690,n21603,n21604,n21605);
  nand U23004(n21605,n21567,G59747);
  nand U23005(n21604,n21566,n21302);
  nand U23006(n21603,n21571,n21606);
  nand U23007(G8689,n21607,n21608,n21609);
  nand U23008(n21609,n21567,G59746);
  nand U23009(n21608,n21566,n21314);
  nand U23010(n21607,n21571,n21610);
  nand U23011(G8688,n21611,n21612,n21613);
  nand U23012(n21613,n21567,G59745);
  nand U23013(n21612,n21566,n21614);
  nand U23014(n21611,n21571,n21328);
  nand U23015(G8687,n21615,n21616,n21617);
  nand U23016(n21617,n21567,G59744);
  nand U23017(n21616,n21566,n21618);
  nand U23018(n21615,n21571,n21339);
  nand U23019(G8686,n21619,n21620,n21621);
  nand U23020(n21621,n21567,G59743);
  nand U23021(n21620,n21566,n21622);
  nand U23022(n21619,n21571,n21349);
  nand U23023(G8685,n21623,n21624,n21625);
  nand U23024(n21625,n21567,G59742);
  nand U23025(n21624,n21566,n21626);
  nand U23026(n21623,n21571,n21359);
  nand U23027(G8684,n21627,n21628,n21629);
  nand U23028(n21629,n21567,G59741);
  nand U23029(n21628,n21566,n21630);
  nand U23030(n21627,n21571,n21369);
  nand U23031(G8683,n21631,n21632,n21633);
  nand U23032(n21633,n21567,G59740);
  nand U23033(n21632,n21566,n21634);
  nand U23034(n21631,n21571,n21379);
  nand U23035(G8682,n21635,n21636,n21637);
  nand U23036(n21637,n21567,G59739);
  nand U23037(n21636,n21566,n21638);
  nand U23038(n21635,n21571,n21389);
  nand U23039(G8681,n21639,n21640,n21641);
  nand U23040(n21641,n21567,G59738);
  nand U23041(n21640,n21566,n21642);
  nand U23042(n21639,n21571,n21399);
  nand U23043(G8680,n21643,n21644,n21645);
  nand U23044(n21645,n21567,G59737);
  nand U23045(n21644,n21566,n21646);
  nand U23046(n21643,n21571,n21409);
  nand U23047(G8679,n21647,n21648,n21649);
  nand U23048(n21649,n21567,G59736);
  nand U23049(n21648,n21566,n21650);
  nand U23050(n21647,n21571,n21422);
  nand U23051(G8678,n21651,n21652,n21653);
  nand U23052(n21653,n21567,G59735);
  nand U23053(n21652,n21566,n21654);
  nand U23054(n21651,n21571,n21432);
  nand U23055(G8677,n21655,n21656,n21657);
  nand U23056(n21657,n21567,G59734);
  nand U23057(n21656,n21566,n21658);
  nand U23058(n21655,n21571,n21442);
  nand U23059(G8676,n21659,n21660,n21661);
  nand U23060(n21661,n21567,G59733);
  nand U23061(n21660,n21566,n21662);
  nand U23062(n21659,n21571,n21452);
  nand U23063(G8675,n21663,n21664,n21665);
  nand U23064(n21665,n21567,G59732);
  nand U23065(n21664,n21566,n21666);
  nand U23066(n21663,n21571,n21463);
  nand U23067(G8674,n21667,n21668,n21669);
  nand U23068(n21669,n21567,G59731);
  nand U23069(n21668,n21566,n21670);
  nand U23070(n21667,n21571,n21475);
  nand U23071(G8673,n21671,n21672,n21673);
  nand U23072(n21673,n21567,G59730);
  nand U23073(n21672,n21566,n21674);
  nand U23074(n21671,n21571,n20986);
  nand U23075(G8672,n21675,n21676,n21677);
  nand U23076(n21677,n21567,G59729);
  nand U23077(n21676,n21566,n21498);
  nand U23078(n21675,n21571,n20996);
  nand U23079(G8671,n21678,n21679,n21680);
  nand U23080(n21680,n21567,G59728);
  nand U23081(n21679,n21566,n21510);
  nand U23082(n21678,n21571,n21006);
  nand U23083(G8670,n21681,n21682,n21683);
  nand U23084(n21683,n21567,G59727);
  nand U23085(n21682,n21566,n21521);
  nand U23086(n21681,n21571,n21015);
  nand U23087(G8669,n21684,n21685,n21686);
  nand U23088(n21686,n21567,G59726);
  nand U23089(n21685,n21566,n21084);
  nand U23090(n21684,n21571,n21030);
  nand U23091(n21689,n21692,n21022);
  nand U23092(G8668,n21693,n21694,n21695,n21696);
  nand U23093(n21696,G58870,n21697);
  nand U23094(n21695,G58902,n21698);
  nand U23095(n21694,n21699,n21178);
  nand U23096(n21693,n21700,G59725);
  nand U23097(G8667,n21701,n21702,n21703,n21704);
  nor U23098(n21704,n21705,n21706,n21707);
  nor U23099(n21707,n21708,n21709);
  nor U23100(n21706,n21710,n21711);
  nor U23101(n21705,n21712,n21713);
  nand U23102(n21703,n21700,G59724);
  nand U23103(n21702,n21699,n21194);
  nand U23104(n21701,n21714,n21195);
  nand U23105(G8666,n21715,n21716,n21717,n21718);
  nor U23106(n21718,n21719,n21720,n21721);
  nor U23107(n21721,n21708,n21722);
  nor U23108(n21720,n21710,n21723);
  nor U23109(n21719,n21713,n21724);
  nand U23110(n21717,n21700,G59723);
  nand U23111(n21716,n21699,n21206);
  nand U23112(n21715,n21714,n21207);
  nand U23113(G8665,n21725,n21726,n21727,n21728);
  nor U23114(n21728,n21729,n21730,n21731);
  nor U23115(n21731,n21708,n21732);
  nor U23116(n21730,n21710,n21733);
  nor U23117(n21729,n21713,n21734);
  nand U23118(n21727,n21700,G59722);
  nand U23119(n21726,n21699,n21218);
  nand U23120(n21725,n21714,n21219);
  nand U23121(G8664,n21735,n21736,n21737,n21738);
  nor U23122(n21738,n21739,n21740,n21741);
  nor U23123(n21741,n21708,n21742);
  nor U23124(n21740,n21710,n21743);
  nor U23125(n21739,n21713,n21744);
  nand U23126(n21737,n21700,G59721);
  nand U23127(n21736,n21699,n21230);
  nand U23128(n21735,n21714,n21231);
  nand U23129(G8663,n21745,n21746,n21747,n21748);
  nor U23130(n21748,n21749,n21750,n21751);
  nor U23131(n21751,n21708,n21752);
  nor U23132(n21750,n21710,n21753);
  nor U23133(n21749,n21713,n21754);
  nand U23134(n21747,n21700,G59720);
  nand U23135(n21746,n21699,n21242);
  nand U23136(n21745,n21714,n21243);
  nand U23137(G8662,n21755,n21756,n21757,n21758);
  nor U23138(n21758,n21759,n21760,n21761);
  nor U23139(n21761,n21708,n21762);
  nor U23140(n21760,n21710,n21763);
  nor U23141(n21759,n21713,n21764);
  nand U23142(n21757,n21700,G59719);
  nand U23143(n21756,n21699,n21254);
  nand U23144(n21755,n21714,n21255);
  nand U23145(G8661,n21765,n21766,n21767,n21768);
  nor U23146(n21768,n21769,n21770,n21771);
  nor U23147(n21771,n21708,n21772);
  not U23148(n21708,n21698);
  nor U23149(n21698,n21773,n21774);
  nor U23150(n21770,n21710,n21775);
  not U23151(n21710,n21697);
  nor U23152(n21697,n21776,n21773);
  nor U23153(n21769,n21713,n21777);
  nand U23154(n21767,n21700,G59718);
  nand U23155(n21766,n21699,n21266);
  nand U23156(n21765,n21714,n21267);
  nand U23157(G8660,n21778,n21779,n21780);
  nor U23158(n21780,n21781,n21782,n21783);
  nor U23159(n21783,n21713,n21784);
  nor U23160(n21782,n21773,n21785);
  nor U23161(n21781,n21786,n21787);
  nand U23162(n21779,n21714,n21279);
  nand U23163(n21778,n21700,G59717);
  nand U23164(G8659,n21788,n21789,n21790);
  nor U23165(n21790,n21791,n21792,n21793);
  nor U23166(n21793,n21713,n21794);
  nor U23167(n21792,n21773,n21795);
  nor U23168(n21791,n21796,n21787);
  nand U23169(n21789,n21714,n21291);
  nand U23170(n21788,n21700,G59716);
  nand U23171(G8658,n21797,n21798,n21799);
  nor U23172(n21799,n21800,n21801,n21802);
  nor U23173(n21802,n21713,n21803);
  nor U23174(n21801,n21773,n21804);
  nor U23175(n21800,n21805,n21787);
  nand U23176(n21798,n21714,n21303);
  nand U23177(n21797,n21700,G59715);
  nand U23178(G8657,n21806,n21807,n21808);
  nor U23179(n21808,n21809,n21810,n21811);
  nor U23180(n21811,n21713,n21812);
  nor U23181(n21810,n21773,n21813);
  nor U23182(n21809,n21814,n21787);
  nand U23183(n21807,n21714,n21315);
  nand U23184(n21806,n21700,G59714);
  nand U23185(G8656,n21815,n21816,n21817);
  nor U23186(n21817,n21818,n21819,n21820);
  nor U23187(n21820,n21713,n21821);
  nor U23188(n21819,n21773,n21822);
  nor U23189(n21818,n21325,n21787);
  nand U23190(n21816,n21714,n21326);
  nand U23191(n21815,n21700,G59713);
  nand U23192(G8655,n21823,n21824,n21825);
  nor U23193(n21825,n21826,n21827,n21828);
  nor U23194(n21828,n21713,n21829);
  nor U23195(n21827,n21773,n21830);
  nor U23196(n21826,n21337,n21787);
  nand U23197(n21824,n21714,n21338);
  nand U23198(n21823,n21700,G59712);
  nand U23199(G8654,n21831,n21832,n21833);
  nor U23200(n21833,n21834,n21835,n21836);
  nor U23201(n21836,n21713,n21837);
  nor U23202(n21835,n21773,n21838);
  nor U23203(n21834,n21347,n21787);
  nand U23204(n21832,n21714,n21348);
  nand U23205(n21831,n21700,G59711);
  nand U23206(G8653,n21839,n21840,n21841);
  nor U23207(n21841,n21842,n21843,n21844);
  nor U23208(n21844,n21713,n21845);
  nand U23209(n21713,n21846,n21847);
  nor U23210(n21843,n21773,n21848);
  nand U23211(n21773,n21849,n21847);
  nor U23212(n21842,n21357,n21787);
  not U23213(n21787,n21699);
  nand U23214(n21840,n21714,n21358);
  nand U23215(n21839,n21700,G59710);
  nand U23216(G8652,n21850,n21851,n21852,n21853);
  nand U23217(n21853,n21854,n21855);
  nand U23218(n21852,n21699,n21630);
  nand U23219(n21851,n21714,n21368);
  nand U23220(n21850,n21700,G59709);
  nand U23221(G8651,n21856,n21857,n21858,n21859);
  nand U23222(n21859,n21854,n21860);
  nand U23223(n21858,n21699,n21634);
  nand U23224(n21857,n21714,n21378);
  nand U23225(n21856,n21700,G59708);
  nand U23226(G8650,n21861,n21862,n21863,n21864);
  nand U23227(n21864,n21854,n21865);
  nand U23228(n21863,n21699,n21638);
  nand U23229(n21862,n21714,n21388);
  nand U23230(n21861,n21700,G59707);
  nand U23231(G8649,n21866,n21867,n21868,n21869);
  nand U23232(n21869,n21854,n21870);
  nand U23233(n21868,n21699,n21642);
  nand U23234(n21867,n21714,n21398);
  nand U23235(n21866,n21700,G59706);
  nand U23236(G8648,n21871,n21872,n21873,n21874);
  nand U23237(n21874,n21854,n21875);
  nand U23238(n21873,n21699,n21646);
  nand U23239(n21872,n21714,n21408);
  nand U23240(n21871,n21700,G59705);
  nand U23241(G8647,n21876,n21877,n21878,n21879);
  nand U23242(n21879,n21854,n21880);
  nand U23243(n21878,n21699,n21650);
  nand U23244(n21877,n21714,n21881);
  nand U23245(n21876,n21700,G59704);
  nand U23246(G8646,n21882,n21883,n21884,n21885);
  nand U23247(n21885,n21854,n21886);
  nand U23248(n21884,n21699,n21654);
  nand U23249(n21883,n21714,n21431);
  nand U23250(n21882,n21700,G59703);
  nand U23251(G8645,n21887,n21888,n21889,n21890);
  nand U23252(n21890,n21854,n21891);
  nand U23253(n21889,n21699,n21658);
  nand U23254(n21888,n21714,n21441);
  nand U23255(n21887,n21700,G59702);
  nand U23256(G8644,n21892,n21893,n21894,n21895);
  nand U23257(n21895,n21854,n21896);
  nand U23258(n21894,n21699,n21662);
  nand U23259(n21893,n21714,n21451);
  nand U23260(n21892,n21700,G59701);
  nand U23261(G8643,n21897,n21898,n21899,n21900);
  nand U23262(n21900,n21854,n21901);
  nand U23263(n21899,n21699,n21666);
  nand U23264(n21898,n21714,n21902);
  nand U23265(n21897,n21700,G59700);
  nand U23266(G8642,n21903,n21904,n21905,n21906);
  nand U23267(n21906,n21854,n21907);
  nand U23268(n21905,n21699,n21670);
  nand U23269(n21904,n21714,n21474);
  nand U23270(n21903,n21700,G59699);
  nand U23271(G8641,n21908,n21909,n21910,n21911);
  nand U23272(n21911,n21854,n21912);
  nand U23273(n21910,n21699,n21674);
  nand U23274(n21909,n21714,n21486);
  nand U23275(n21908,n21700,G59698);
  nand U23276(G8640,n21913,n21914,n21915,n21916);
  nand U23277(n21916,n21854,n21917);
  nand U23278(n21915,n21699,n21498);
  nand U23279(n21914,n21714,n21499);
  nand U23280(n21913,n21700,G59697);
  nand U23281(G8639,n21918,n21919,n21920,n21921);
  nand U23282(n21921,n21854,n21922);
  nand U23283(n21920,n21699,n21510);
  nand U23284(n21919,n21714,n21511);
  nand U23285(n21918,n21700,G59696);
  nand U23286(G8638,n21923,n21924,n21925,n21926);
  nand U23287(n21926,n21854,n21927);
  nand U23288(n21925,n21699,n21521);
  nand U23289(n21924,n21714,n21522);
  nand U23290(n21923,n21700,G59695);
  nand U23291(G8637,n21928,n21929,n21930,n21931);
  nand U23292(n21931,n21854,n21932);
  nor U23293(n21854,n21700,n21933);
  nand U23294(n21930,n21699,n21084);
  nor U23295(n21699,n21934,n21700);
  nand U23296(n21929,n21714,n21546);
  nand U23297(n21928,n21700,G59694);
  nand U23298(n21847,n21936,n21937);
  nand U23299(n21937,n20985,n21938);
  nand U23300(n21938,n21939,n21940);
  nand U23301(n21940,n21941,n21080);
  nand U23302(n21941,n21113,n21942);
  or U23303(n21942,n21943,n21944);
  nor U23304(G8636,n21945,n21946);
  nand U23305(G8635,n21947,n21948,n21949);
  nand U23306(n21949,G59692,n21950);
  nand U23307(n21948,n21951,G59724);
  nand U23308(n21947,G59647,n21952);
  nand U23309(G8634,n21953,n21954,n21955);
  nand U23310(n21955,G59691,n21950);
  nand U23311(n21954,n21951,G59723);
  nand U23312(n21953,G59648,n21952);
  nand U23313(G8633,n21956,n21957,n21958);
  nand U23314(n21958,G59690,n21950);
  nand U23315(n21957,n21951,G59722);
  nand U23316(n21956,G59649,n21952);
  nand U23317(G8632,n21959,n21960,n21961);
  nand U23318(n21961,G59689,n21950);
  nand U23319(n21960,n21951,G59721);
  nand U23320(n21959,G59650,n21952);
  nand U23321(G8631,n21962,n21963,n21964);
  nand U23322(n21964,G59688,n21950);
  nand U23323(n21963,n21951,G59720);
  nand U23324(n21962,G59651,n21952);
  nand U23325(G8630,n21965,n21966,n21967);
  nand U23326(n21967,G59687,n21950);
  nand U23327(n21966,n21951,G59719);
  nand U23328(n21965,G59652,n21952);
  nand U23329(G8629,n21968,n21969,n21970);
  nand U23330(n21970,G59686,n21950);
  nand U23331(n21969,n21951,G59718);
  nand U23332(n21968,G59653,n21952);
  nand U23333(G8628,n21971,n21972,n21973);
  nand U23334(n21973,G59685,n21950);
  nand U23335(n21972,n21951,G59717);
  nand U23336(n21971,G59654,n21952);
  nand U23337(G8627,n21974,n21975,n21976);
  nand U23338(n21976,G59684,n21950);
  nand U23339(n21975,n21951,G59716);
  nand U23340(n21974,G59655,n21952);
  nand U23341(G8626,n21977,n21978,n21979);
  nand U23342(n21979,G59683,n21950);
  nand U23343(n21978,n21951,G59715);
  nand U23344(n21977,G59656,n21952);
  nand U23345(G8625,n21980,n21981,n21982);
  nand U23346(n21982,G59682,n21950);
  nand U23347(n21981,n21951,G59714);
  nand U23348(n21980,G59657,n21952);
  nand U23349(G8624,n21983,n21984,n21985);
  nand U23350(n21985,G59681,n21950);
  nand U23351(n21984,n21951,G59713);
  nand U23352(n21983,G59658,n21952);
  nand U23353(G8623,n21986,n21987,n21988);
  nand U23354(n21988,G59680,n21950);
  nand U23355(n21987,n21951,G59712);
  nand U23356(n21986,G59659,n21952);
  nand U23357(G8622,n21989,n21990,n21991);
  nand U23358(n21991,G59679,n21950);
  nand U23359(n21990,n21951,G59711);
  nand U23360(n21989,G59660,n21952);
  nand U23361(G8621,n21992,n21993,n21994);
  nand U23362(n21994,G59678,n21950);
  nand U23363(n21993,n21951,G59710);
  and U23364(n21951,n21995,n21846);
  nand U23365(n21992,G59661,n21952);
  nand U23366(G8620,n21996,n21997,n21998);
  nand U23367(n21998,G59677,n21950);
  nand U23368(n21997,G59631,n21952);
  nand U23369(n21996,n21995,G59709);
  nand U23370(G8619,n21999,n22000,n22001);
  nand U23371(n22001,G59676,n21950);
  nand U23372(n22000,G59632,n21952);
  nand U23373(n21999,n21995,G59708);
  nand U23374(G8618,n22002,n22003,n22004);
  nand U23375(n22004,G59675,n21950);
  nand U23376(n22003,G59633,n21952);
  nand U23377(n22002,n21995,G59707);
  nand U23378(G8617,n22005,n22006,n22007);
  nand U23379(n22007,G59674,n21950);
  nand U23380(n22006,G59634,n21952);
  nand U23381(n22005,n21995,G59706);
  nand U23382(G8616,n22008,n22009,n22010);
  nand U23383(n22010,G59673,n21950);
  nand U23384(n22009,G59635,n21952);
  nand U23385(n22008,n21995,G59705);
  nand U23386(G8615,n22011,n22012,n22013);
  nand U23387(n22013,G59672,n21950);
  nand U23388(n22012,G59636,n21952);
  nand U23389(n22011,n21995,G59704);
  nand U23390(G8614,n22014,n22015,n22016);
  nand U23391(n22016,G59671,n21950);
  nand U23392(n22015,G59637,n21952);
  nand U23393(n22014,n21995,G59703);
  nand U23394(G8613,n22017,n22018,n22019);
  nand U23395(n22019,G59670,n21950);
  nand U23396(n22018,G59638,n21952);
  nand U23397(n22017,n21995,G59702);
  nand U23398(G8612,n22020,n22021,n22022);
  nand U23399(n22022,G59669,n21950);
  nand U23400(n22021,G59639,n21952);
  nand U23401(n22020,n21995,G59701);
  nand U23402(G8611,n22023,n22024,n22025);
  nand U23403(n22025,G59668,n21950);
  nand U23404(n22024,G59640,n21952);
  nand U23405(n22023,n21995,G59700);
  nand U23406(G8610,n22026,n22027,n22028);
  nand U23407(n22028,G59667,n21950);
  nand U23408(n22027,G59641,n21952);
  nand U23409(n22026,n21995,G59699);
  nand U23410(G8609,n22029,n22030,n22031);
  nand U23411(n22031,G59666,n21950);
  nand U23412(n22030,G59642,n21952);
  nand U23413(n22029,n21995,G59698);
  nand U23414(G8608,n22032,n22033,n22034);
  nand U23415(n22034,G59665,n21950);
  nand U23416(n22033,G59643,n21952);
  nand U23417(n22032,n21995,G59697);
  nand U23418(G8607,n22035,n22036,n22037);
  nand U23419(n22037,G59664,n21950);
  nand U23420(n22036,G59644,n21952);
  nand U23421(n22035,n21995,G59696);
  nand U23422(G8606,n22038,n22039,n22040);
  nand U23423(n22040,G59663,n21950);
  nand U23424(n22039,G59645,n21952);
  nand U23425(n22038,n21995,G59695);
  nand U23426(G8605,n22041,n22042,n22043);
  nand U23427(n22043,G59662,n21950);
  nand U23428(n22042,G59646,n21952);
  nand U23429(n22041,n21995,G59694);
  nor U23430(n21995,n21531,n21950);
  nand U23431(n21945,n22044,n22045);
  nand U23432(n22045,n22046,n21080);
  nand U23433(n22046,n22047,n22048);
  nand U23434(n22048,n21022,n21060,n22049);
  nand U23435(n22047,n20985,n22050,n22051);
  nand U23436(n22044,n21046,G59427);
  nand U23437(G8604,n22052,n22053,n22054);
  nand U23438(n22054,n22055,G59661);
  nand U23439(n22052,n22056,G59710);
  nand U23440(G8603,n22057,n22058,n22059);
  nand U23441(n22059,n22055,G59660);
  nand U23442(n22057,n22056,G59711);
  nand U23443(G8602,n22060,n22061,n22062);
  nand U23444(n22062,n22055,G59659);
  nand U23445(n22060,n22056,G59712);
  nand U23446(G8601,n22063,n22064,n22065);
  nand U23447(n22065,n22055,G59658);
  nand U23448(n22063,n22056,G59713);
  nand U23449(G8600,n22066,n22067,n22068);
  nand U23450(n22068,n22055,G59657);
  nand U23451(n22066,n22056,G59714);
  nand U23452(G8599,n22069,n22070,n22071);
  nand U23453(n22071,n22055,G59656);
  nand U23454(n22069,n22056,G59715);
  nand U23455(G8598,n22072,n22073,n22074);
  nand U23456(n22074,n22055,G59655);
  nand U23457(n22072,n22056,G59716);
  nand U23458(G8597,n22075,n22076,n22077);
  nand U23459(n22077,n22055,G59654);
  nand U23460(n22075,n22056,G59717);
  nand U23461(G8596,n22078,n22079,n22080);
  nand U23462(n22080,n22055,G59653);
  nand U23463(n22078,n22056,G59718);
  nand U23464(G8595,n22081,n22082,n22083);
  nand U23465(n22083,n22055,G59652);
  nand U23466(n22081,n22056,G59719);
  nand U23467(G8594,n22084,n22085,n22086);
  nand U23468(n22086,n22055,G59651);
  nand U23469(n22084,n22056,G59720);
  nand U23470(G8593,n22087,n22088,n22089);
  nand U23471(n22089,n22055,G59650);
  nand U23472(n22087,n22056,G59721);
  nand U23473(G8592,n22090,n22091,n22092);
  nand U23474(n22092,n22055,G59649);
  nand U23475(n22090,n22056,G59722);
  nand U23476(G8591,n22093,n22094,n22095);
  nand U23477(n22095,n22055,G59648);
  nand U23478(n22093,n22056,G59723);
  nand U23479(G8590,n22096,n22097,n22098);
  nand U23480(n22098,n22055,G59647);
  nand U23481(n22096,n22056,G59724);
  nand U23482(G8589,n22099,n22053,n22100);
  nand U23483(n22100,n22055,G59646);
  nand U23484(n22053,n22101,n21932);
  nand U23485(n22099,n22056,G59694);
  nand U23486(G8588,n22102,n22058,n22103);
  nand U23487(n22103,n22055,G59645);
  nand U23488(n22058,n22101,n21927);
  nand U23489(n22102,n22056,G59695);
  nand U23490(G8587,n22104,n22061,n22105);
  nand U23491(n22105,n22055,G59644);
  nand U23492(n22061,n22101,n21922);
  nand U23493(n22104,n22056,G59696);
  nand U23494(G8586,n22106,n22064,n22107);
  nand U23495(n22107,n22055,G59643);
  nand U23496(n22064,n22101,n21917);
  nand U23497(n22106,n22056,G59697);
  nand U23498(G8585,n22108,n22067,n22109);
  nand U23499(n22109,n22055,G59642);
  nand U23500(n22067,n22101,n21912);
  nand U23501(n22108,n22056,G59698);
  nand U23502(G8584,n22110,n22070,n22111);
  nand U23503(n22111,n22055,G59641);
  nand U23504(n22070,n22101,n21907);
  nand U23505(n22110,n22056,G59699);
  nand U23506(G8583,n22112,n22073,n22113);
  nand U23507(n22113,n22055,G59640);
  nand U23508(n22073,n22101,n21901);
  nand U23509(n22112,n22056,G59700);
  nand U23510(G8582,n22114,n22076,n22115);
  nand U23511(n22115,n22055,G59639);
  nand U23512(n22076,n22101,n21896);
  nand U23513(n22114,n22056,G59701);
  nand U23514(G8581,n22116,n22079,n22117);
  nand U23515(n22117,n22055,G59638);
  nand U23516(n22079,n22101,n21891);
  not U23517(n21891,n21777);
  nand U23518(n21777,n22118,n22119);
  nand U23519(n22119,n21774,n22120);
  nand U23520(n22118,n21776,n22121);
  nand U23521(n22116,n22056,G59702);
  nand U23522(G8580,n22122,n22082,n22123);
  nand U23523(n22123,n22055,G59637);
  nand U23524(n22082,n22101,n21886);
  not U23525(n21886,n21764);
  nand U23526(n21764,n22124,n22125);
  nand U23527(n22125,n21774,n22126);
  nand U23528(n22124,n21776,n22127);
  nand U23529(n22122,n22056,G59703);
  nand U23530(G8579,n22128,n22085,n22129);
  nand U23531(n22129,n22055,G59636);
  nand U23532(n22085,n22101,n21880);
  not U23533(n21880,n21754);
  nand U23534(n21754,n22130,n22131);
  nand U23535(n22131,n21774,n22132);
  nand U23536(n22130,n21776,n22133);
  nand U23537(n22128,n22056,G59704);
  nand U23538(G8578,n22134,n22088,n22135);
  nand U23539(n22135,n22055,G59635);
  nand U23540(n22088,n22101,n21875);
  not U23541(n21875,n21744);
  nand U23542(n21744,n22136,n22137);
  nand U23543(n22137,n21774,n22138);
  nand U23544(n22136,n21776,n22139);
  nand U23545(n22134,n22056,G59705);
  nand U23546(G8577,n22140,n22091,n22141);
  nand U23547(n22141,n22055,G59634);
  nand U23548(n22091,n22101,n21870);
  not U23549(n21870,n21734);
  nand U23550(n21734,n22142,n22143);
  nand U23551(n22143,n21774,n22144);
  nand U23552(n22142,n21776,n22145);
  nand U23553(n22140,n22056,G59706);
  nand U23554(G8576,n22146,n22094,n22147);
  nand U23555(n22147,n22055,G59633);
  nand U23556(n22094,n22101,n21865);
  not U23557(n21865,n21724);
  nand U23558(n21724,n22148,n22149);
  nand U23559(n22149,n21774,n22150);
  nand U23560(n22148,n21776,n22151);
  nand U23561(n22146,n22056,G59707);
  nand U23562(G8575,n22152,n22097,n22153);
  nand U23563(n22153,n22055,G59632);
  nand U23564(n22097,n22101,n21860);
  not U23565(n21860,n21712);
  nand U23566(n21712,n22154,n22155);
  nand U23567(n22155,n21774,n22156);
  nand U23568(n22154,n21776,n22157);
  nand U23569(n22152,n22056,G59708);
  nand U23570(G8574,n22158,n22159,n22160);
  nand U23571(n22160,n22055,G59631);
  nand U23572(n22159,n22101,n21855);
  nand U23573(n21855,n22161,n22162);
  nand U23574(n22162,G58886,n21776);
  nand U23575(n22161,G58854,n21774);
  nor U23576(n22101,n22163,n22055);
  nand U23577(n22158,n22056,G59709);
  nand U23578(n22164,n21022,n21080,n22165);
  nand U23579(n21936,n21556,n21045);
  nor U23580(n21556,n22166,n21105,n22167);
  nand U23581(G8573,n22168,n22169,n22170,n22171);
  nor U23582(n22171,n22172,n22173);
  nor U23583(n22173,n21172,n22174);
  nor U23584(n22172,n21545,n22175);
  nand U23585(n22170,n22176,n21181);
  nand U23586(n22169,n22177,G59789);
  nand U23587(n22168,n22178,n21175);
  nand U23588(G8572,n22179,n22180,n22181,n22182);
  nor U23589(n22182,n22183,n22184);
  nor U23590(n22184,n21190,n22174);
  nor U23591(n22183,n22185,n22175);
  nand U23592(n22181,n22176,n21195);
  nand U23593(n22180,n22177,G59788);
  nand U23594(n22179,n22178,n21572);
  nand U23595(G8571,n22186,n22187,n22188,n22189);
  nor U23596(n22189,n22190,n22191);
  nor U23597(n22191,n21203,n22174);
  nor U23598(n22190,n22192,n22175);
  nand U23599(n22188,n22176,n21207);
  nand U23600(n22187,n22177,G59787);
  nand U23601(n22186,n22178,n21576);
  nand U23602(G8570,n22193,n22194,n22195,n22196);
  nor U23603(n22196,n22197,n22198);
  nor U23604(n22198,n21215,n22174);
  nor U23605(n22197,n22199,n22175);
  nand U23606(n22195,n22176,n21219);
  nand U23607(n22194,n22177,G59786);
  nand U23608(n22193,n22178,n21580);
  nand U23609(G8569,n22200,n22201,n22202,n22203);
  nor U23610(n22203,n22204,n22205);
  nor U23611(n22205,n21227,n22174);
  and U23612(n22204,n21230,n22206);
  nand U23613(n22202,n22176,n21231);
  nand U23614(n22201,n22177,G59785);
  nand U23615(n22200,n22178,n21584);
  nand U23616(G8568,n22207,n22208,n22209,n22210);
  nor U23617(n22210,n22211,n22212);
  nor U23618(n22212,n21239,n22174);
  nor U23619(n22211,n22213,n22175);
  nand U23620(n22209,n22176,n21243);
  nand U23621(n22208,n22177,G59784);
  nand U23622(n22207,n22178,n21588);
  nand U23623(G8567,n22214,n22215,n22216,n22217);
  nor U23624(n22217,n22218,n22219);
  nor U23625(n22219,n21251,n22174);
  and U23626(n22218,n21254,n22206);
  nand U23627(n22216,n22176,n21255);
  nand U23628(n22215,n22177,G59783);
  nand U23629(n22214,n22178,n21252);
  nand U23630(G8566,n22220,n22221,n22222,n22223);
  nor U23631(n22223,n22224,n22225);
  nor U23632(n22225,n21263,n22174);
  nor U23633(n22224,n22226,n22175);
  nand U23634(n22222,n22176,n21267);
  nand U23635(n22221,n22177,G59782);
  nand U23636(n22220,n22178,n21595);
  nand U23637(G8565,n22227,n22228,n22229,n22230);
  nor U23638(n22230,n22231,n22232);
  nor U23639(n22232,n21275,n22174);
  nor U23640(n22231,n21786,n22175);
  nand U23641(n22229,n22176,n21279);
  nand U23642(n22228,n22177,G59781);
  nand U23643(n22227,n22178,n21599);
  nand U23644(G8564,n22233,n22234,n22235,n22236);
  nor U23645(n22236,n22237,n22238);
  nor U23646(n22238,n21287,n22174);
  not U23647(n21287,G59621);
  nor U23648(n22237,n21796,n22175);
  nand U23649(n22235,n22176,n21291);
  nand U23650(n22234,n22177,G59780);
  nand U23651(n22233,n22178,n21288);
  nand U23652(G8563,n22239,n22240,n22241,n22242);
  nor U23653(n22242,n22243,n22244);
  nor U23654(n22244,n21299,n22174);
  not U23655(n21299,G59620);
  nor U23656(n22243,n21805,n22175);
  nand U23657(n22241,n22176,n21303);
  nand U23658(n22240,n22177,G59779);
  nand U23659(n22239,n22178,n21606);
  nand U23660(G8562,n22245,n22246,n22247,n22248);
  nor U23661(n22248,n22249,n22250);
  nor U23662(n22250,n21311,n22174);
  not U23663(n21311,G59619);
  nor U23664(n22249,n21814,n22175);
  nand U23665(n22247,n22176,n21315);
  nand U23666(n22246,n22177,G59778);
  nand U23667(n22245,n22178,n21610);
  nand U23668(G8561,n22251,n22252,n22253,n22254);
  nor U23669(n22254,n22255,n22256);
  and U23670(n22256,G59618,n22257);
  nor U23671(n22255,n21325,n22175);
  nand U23672(n22253,n22176,n21326);
  nand U23673(n22252,n22177,G59777);
  nand U23674(n22251,n22178,n21328);
  nand U23675(G8560,n22258,n22259,n22260,n22261);
  nor U23676(n22261,n22262,n22263);
  and U23677(n22263,G59617,n22257);
  nor U23678(n22262,n21337,n22175);
  nand U23679(n22260,n22176,n21338);
  nand U23680(n22259,n22177,G59776);
  nand U23681(n22258,n22178,n21339);
  nand U23682(G8559,n22264,n22265,n22266,n22267);
  nor U23683(n22267,n22268,n22269);
  and U23684(n22269,G59616,n22257);
  nor U23685(n22268,n21347,n22175);
  nand U23686(n22266,n22176,n21348);
  nand U23687(n22265,n22177,G59775);
  nand U23688(n22264,n22178,n21349);
  nand U23689(G8558,n22270,n22271,n22272,n22273);
  nor U23690(n22273,n22274,n22275);
  and U23691(n22275,G59615,n22257);
  nor U23692(n22274,n21357,n22175);
  nand U23693(n22272,n22176,n21358);
  nand U23694(n22271,n22177,G59774);
  nand U23695(n22270,n22178,n21359);
  nand U23696(G8557,n22276,n22277,n22278,n22279);
  nor U23697(n22279,n22280,n22281);
  and U23698(n22281,G59614,n22257);
  nor U23699(n22280,n21367,n22175);
  nand U23700(n22278,n22176,n21368);
  nand U23701(n22277,n22177,G59773);
  nand U23702(n22276,n22178,n21369);
  nand U23703(G8556,n22282,n22283,n22284,n22285);
  nor U23704(n22285,n22286,n22287);
  and U23705(n22287,G59613,n22257);
  nor U23706(n22286,n21377,n22175);
  nand U23707(n22284,n22176,n21378);
  nand U23708(n22283,n22177,G59772);
  nand U23709(n22282,n22178,n21379);
  nand U23710(G8555,n22288,n22289,n22290,n22291);
  nor U23711(n22291,n22292,n22293);
  and U23712(n22293,G59612,n22257);
  nor U23713(n22292,n21387,n22175);
  nand U23714(n22290,n22176,n21388);
  nand U23715(n22289,n22177,G59771);
  nand U23716(n22288,n22178,n21389);
  nand U23717(G8554,n22294,n22295,n22296,n22297);
  nor U23718(n22297,n22298,n22299);
  and U23719(n22299,G59611,n22257);
  nor U23720(n22298,n21397,n22175);
  nand U23721(n22296,n22176,n21398);
  nand U23722(n22295,n22177,G59770);
  nand U23723(n22294,n22178,n21399);
  nand U23724(G8553,n22300,n22301,n22302,n22303);
  nor U23725(n22303,n22304,n22305);
  and U23726(n22305,G59610,n22257);
  nor U23727(n22304,n21407,n22175);
  nand U23728(n22302,n22176,n21408);
  nand U23729(n22301,n22177,G59769);
  nand U23730(n22300,n22178,n21409);
  nand U23731(G8552,n22306,n22307,n22308);
  nor U23732(n22308,n22309,n22310,n22311);
  nor U23733(n22311,n22312,n22313);
  nor U23734(n22310,n22314,n22315);
  and U23735(n22309,n21881,n22176);
  nand U23736(n22307,n22206,n21650);
  nand U23737(n22306,n22257,G59609);
  nand U23738(G8551,n22316,n22317,n22318,n22319);
  nor U23739(n22319,n22320,n22321);
  and U23740(n22321,G59608,n22257);
  nor U23741(n22320,n21430,n22175);
  nand U23742(n22318,n22176,n21431);
  nand U23743(n22317,n22177,G59767);
  nand U23744(n22316,n22178,n21432);
  nand U23745(G8550,n22322,n22323,n22324,n22325);
  nor U23746(n22325,n22326,n22327);
  and U23747(n22327,G59607,n22257);
  nor U23748(n22326,n21440,n22175);
  not U23749(n21440,n21658);
  nand U23750(n22324,n22176,n21441);
  nand U23751(n22323,n22177,G59766);
  nand U23752(n22322,n22178,n21442);
  nand U23753(G8549,n22328,n22329,n22330,n22331);
  nor U23754(n22331,n22332,n22333);
  and U23755(n22333,G59606,n22257);
  nor U23756(n22332,n21450,n22175);
  nand U23757(n22330,n22176,n21451);
  nand U23758(n22329,n22177,G59765);
  nand U23759(n22328,n22178,n21452);
  nand U23760(G8548,n22334,n22335,n22336,n22337);
  nor U23761(n22337,n22338,n22339);
  nor U23762(n22339,n22340,n22174);
  nor U23763(n22338,n21460,n22175);
  nand U23764(n22336,n22176,n21902);
  nand U23765(n22335,n22177,G59764);
  nand U23766(n22334,n22178,n21463);
  nand U23767(G8547,n22341,n22342,n22343,n22344);
  nor U23768(n22344,n22345,n22346);
  nor U23769(n22346,n22347,n22174);
  nor U23770(n22345,n21471,n22175);
  nand U23771(n22343,n22176,n21474);
  nand U23772(n22342,n22177,G59763);
  nand U23773(n22341,n22178,n21475);
  nand U23774(G8546,n22348,n22349,n22350,n22351);
  nor U23775(n22351,n22352,n22353);
  nor U23776(n22353,n22354,n22174);
  nor U23777(n22352,n21484,n22175);
  nand U23778(n22350,n22176,n21486);
  nand U23779(n22349,n22177,G59762);
  nand U23780(n22348,n22178,n20986);
  nand U23781(G8545,n22355,n22356,n22357,n22358);
  nor U23782(n22358,n22359,n22360);
  nor U23783(n22360,n21494,n22174);
  nor U23784(n22359,n22361,n22175);
  nand U23785(n22357,n22176,n21499);
  nand U23786(n22356,n22177,G59761);
  nand U23787(n22355,n22178,n20996);
  nand U23788(G8544,n22362,n22363,n22364,n22365);
  nor U23789(n22365,n22366,n22367);
  nor U23790(n22367,n21507,n22174);
  nor U23791(n22366,n22368,n22175);
  nand U23792(n22364,n22176,n21511);
  nand U23793(n22363,n22177,G59760);
  nand U23794(n22362,n22178,n21006);
  nand U23795(G8543,n22369,n22370,n22371,n22372);
  nor U23796(n22372,n22373,n22374);
  nor U23797(n22374,n21519,n22174);
  nor U23798(n22373,n22375,n22175);
  not U23799(n22175,n22206);
  nand U23800(n22371,n22176,n21522);
  nand U23801(n22370,n22177,G59759);
  nand U23802(n22369,n22178,n21015);
  nand U23803(G8542,n22376,n22377,n22378,n22379);
  nand U23804(n22379,n22176,n21546);
  nor U23805(n22378,n22380,n22381);
  nor U23806(n22381,n21532,n22313);
  not U23807(n22313,n22178);
  nor U23808(n22380,n21122,n22315);
  not U23809(n22315,n22177);
  nand U23810(n22377,n22206,n21084);
  nor U23811(n22206,n22383,n22257);
  nand U23812(n22376,n22257,G59599);
  not U23813(n22257,n22174);
  nand U23814(n22174,n21116,n21042);
  nand U23815(n21042,n21043,n21531,n22384);
  or U23816(n21116,n21106,n21105);
  nand U23817(n21106,n22385,G59426,n22386);
  nand U23818(G8541,n22387,n22388,n22389,n22390);
  nor U23819(n22390,n22391,n22392,n22393);
  nor U23820(n22393,G59598,n22394,n22395);
  nor U23821(n22392,n22396,n22397);
  nor U23822(n22396,n22398,n22399);
  and U23823(n22398,n22395,n22400);
  nor U23824(n22391,n21176,n22401);
  nand U23825(n22389,n22402,n21178);
  nand U23826(n22388,n22403,n21181);
  nand U23827(n21181,n22404,n22405);
  nand U23828(n22405,n22406,n22407);
  nand U23829(n22407,n22408,n22409);
  nand U23830(n22408,n22410,n22411,n22412);
  nand U23831(n22404,n22413,n22409,n22414);
  nand U23832(n22409,n22415,n22416,n22417);
  nand U23833(n22415,n22418,n22414);
  nand U23834(n22413,n22412,n22418);
  not U23835(n22412,n22416);
  nand U23836(n22416,n22419,n22420,n22421,n22422);
  nand U23837(n22422,n21175,n22423);
  nand U23838(n22421,n22406,n21178);
  not U23839(n21178,n21545);
  xor U23840(n21545,n22424,n22425);
  nand U23841(n22424,n22426,n22427);
  nand U23842(n22427,n22428,n21108);
  nand U23843(n22426,n22429,n22167);
  nand U23844(n22429,n22430,n22431,n22428);
  and U23845(n22428,n22432,n22433);
  nand U23846(n22433,G59757,n22434);
  nand U23847(n22432,G59630,n22435);
  nand U23848(n22431,G59598,n22436);
  nand U23849(n22430,G59725,n22437);
  nand U23850(n22420,G59598,n22438);
  nand U23851(n22419,n22439,G59789);
  nand U23852(n22387,n22440,n21175);
  xor U23853(n21175,n22441,n22442);
  nor U23854(n22442,n22443,n22444,n22445);
  nor U23855(n22445,n22382,n21172);
  not U23856(n21172,G59630);
  nor U23857(n22444,n22446,n22397);
  nor U23858(n22443,n22167,n21176);
  not U23859(n21176,G59789);
  nand U23860(G8540,n22447,n22448,n22449,n22450);
  nor U23861(n22450,n22451,n22452,n22453);
  nor U23862(n22453,n21193,n22401);
  nor U23863(n22452,n22454,n22394);
  nor U23864(n22451,n22455,n22456);
  nand U23865(n22449,n22402,n21194);
  nand U23866(n22448,n22403,n21195);
  nand U23867(n21195,n22457,n22458);
  nand U23868(n22458,n22406,n22459);
  nand U23869(n22459,n22418,n22417);
  nand U23870(n22417,n22410,n22411);
  not U23871(n22410,n22460);
  nand U23872(n22418,n22460,n22461);
  nand U23873(n22457,n22462,n22414);
  xnor U23874(n22462,n22460,n22411);
  not U23875(n22411,n22461);
  nand U23876(n22461,n22463,n22464,n22465,n22466);
  nor U23877(n22466,n22467,n22468);
  nor U23878(n22468,n21193,n22469);
  nor U23879(n22467,n22470,n22455);
  nand U23880(n22465,n22406,n21194);
  nand U23881(n22464,n22471,n22472,n22473);
  nand U23882(n22472,n21572,n22474);
  nand U23883(n22471,n22475,n21192);
  nand U23884(n22475,n22476,n22474);
  nor U23885(n22474,n21204,n21216);
  nand U23886(n22463,n21572,n22477);
  nand U23887(n22460,n22478,n22479);
  nand U23888(n22479,n22406,n22480);
  nand U23889(n22480,n22481,n22482);
  or U23890(n22478,n22482,n22481);
  nand U23891(n22447,n22440,n21572);
  not U23892(n21572,n21192);
  nand U23893(n21192,n22483,n22441);
  nand U23894(n22441,n22484,n22485,n22486);
  xnor U23895(n22486,n22487,n22383);
  nand U23896(n22483,n22488,n22489);
  nand U23897(n22489,n22485,n22484);
  xnor U23898(n22488,n22435,n22487);
  nand U23899(n22487,n22490,n22491,n22492,n22493);
  nor U23900(n22493,n22494,n22495);
  nor U23901(n22495,n22382,n21190);
  not U23902(n21190,G59629);
  nor U23903(n22494,n22167,n21193);
  not U23904(n21193,G59788);
  nand U23905(n22492,G59597,n22496);
  nand U23906(n22491,n21194,n22497);
  not U23907(n21194,n22185);
  nand U23908(n22185,n22425,n22498);
  nand U23909(n22498,n22499,n22500);
  or U23910(n22425,n22500,n22499);
  xor U23911(n22499,n22501,n22167);
  nand U23912(n22501,n22502,n22503,n22504,n22505);
  nor U23913(n22505,n22506,n22507);
  and U23914(n22507,n22437,G59724);
  nor U23915(n22506,n22508,n22455);
  not U23916(n22455,G59597);
  nand U23917(n22504,G59629,n22435);
  or U23918(n22503,n22454,n21114);
  nand U23919(n22454,n22509,n22395);
  nand U23920(n22395,n22510,n22511);
  or U23921(n22509,n22511,n22510);
  nand U23922(n22511,n22512,n22513);
  nand U23923(n22513,G59597,n21058);
  nand U23924(n22512,n22514,n21846);
  nand U23925(n22514,n22515,n22516,n22517,n22518);
  nor U23926(n22518,n22519,n22520,n22521,n22522);
  nor U23927(n22522,n22523,n22524);
  nor U23928(n22521,n22525,n22526);
  nor U23929(n22520,n22527,n22528);
  nor U23930(n22519,n22529,n22530);
  nor U23931(n22517,n22531,n22532,n22533,n22534);
  nor U23932(n22534,n22535,n22536);
  nor U23933(n22533,n22537,n22538);
  nor U23934(n22532,n22539,n22540);
  nor U23935(n22531,n22541,n22542);
  nor U23936(n22516,n22543,n22544,n22545,n22546);
  nor U23937(n22546,n22547,n22548);
  nor U23938(n22545,n22549,n22550);
  nor U23939(n22544,n22551,n22552);
  nor U23940(n22543,n22553,n22554);
  nor U23941(n22515,n22555,n22556,n22557,n22558);
  nor U23942(n22558,n22559,n22560);
  nor U23943(n22557,n22561,n22562);
  nor U23944(n22556,n22563,n22564);
  nor U23945(n22555,n22565,n22566);
  nand U23946(n22502,G59756,n22434);
  nand U23947(n22490,n22567,n22568);
  nand U23948(G8539,n22569,n22570,n22571,n22572);
  nor U23949(n22572,n22573,n22574,n22575);
  nor U23950(n22575,n21205,n22401);
  nor U23951(n22574,n22576,n22394);
  nor U23952(n22573,n22577,n22456);
  nand U23953(n22571,n22402,n21206);
  nand U23954(n22570,n22403,n21207);
  xnor U23955(n21207,n22481,n22578);
  xnor U23956(n22578,n22406,n22482);
  nand U23957(n22482,n22579,n22580);
  nand U23958(n22580,n22581,n22414);
  nand U23959(n22581,n22582,n22583);
  or U23960(n22579,n22582,n22583);
  and U23961(n22481,n22584,n22585,n22586,n22587);
  nor U23962(n22587,n22588,n22589);
  nor U23963(n22589,n21205,n22469);
  nor U23964(n22588,n22470,n22577);
  nand U23965(n22586,n22406,n21206);
  nand U23966(n22585,n22590,n22591,n22473);
  nand U23967(n22591,n21216,n21204);
  nand U23968(n22590,n21580,n22592);
  nand U23969(n22592,n22476,n21204);
  nand U23970(n22584,n21576,n22477);
  nand U23971(n22569,n22440,n21576);
  not U23972(n21576,n21204);
  xnor U23973(n21204,n22484,n22485);
  nor U23974(n22485,n22593,n22594);
  xnor U23975(n22484,n22595,n22383);
  nand U23976(n22595,n22596,n22597,n22598,n22599);
  nor U23977(n22599,n22600,n22601);
  nor U23978(n22601,n22382,n21203);
  not U23979(n21203,G59628);
  nor U23980(n22600,n22167,n21205);
  not U23981(n21205,G59787);
  nand U23982(n22598,G59596,n22496);
  nand U23983(n22597,n21206,n22497);
  not U23984(n21206,n22192);
  nand U23985(n22192,n22500,n22602);
  nand U23986(n22602,n22603,n22604);
  or U23987(n22500,n22604,n22603);
  xor U23988(n22603,n22605,n22167);
  nand U23989(n22605,n22606,n22607,n22608,n22609);
  nor U23990(n22609,n22610,n22611);
  and U23991(n22611,n22434,G59755);
  and U23992(n22610,n22437,G59723);
  nand U23993(n22608,G59628,n22435);
  or U23994(n22607,n22576,n21114);
  nand U23995(n22576,n22612,n22613);
  nand U23996(n22613,n22614,n22615);
  not U23997(n22612,n22510);
  nor U23998(n22510,n22615,n22614);
  nand U23999(n22614,n22616,n22617);
  nand U24000(n22617,n21058,n22577);
  not U24001(n22577,G59596);
  nand U24002(n22616,n22618,n22619,n22620,n21846);
  nor U24003(n22620,n22621,n22622);
  nand U24004(n22622,n22623,n22624,n22625,n22626);
  nand U24005(n22626,n22627,G59550);
  nand U24006(n22625,n22628,G59542);
  nand U24007(n22624,n22629,G59534);
  nand U24008(n22623,n22630,G59526);
  nand U24009(n22621,n22631,n22632,n22633,n22634);
  nand U24010(n22634,n22635,G59518);
  nand U24011(n22633,n22636,G59510);
  nand U24012(n22632,n22637,G59502);
  nand U24013(n22631,n22638,G59494);
  nor U24014(n22619,n22639,n22640,n22641,n22642);
  nor U24015(n22642,n22643,n22524);
  nor U24016(n22641,n22644,n22526);
  nor U24017(n22640,n22645,n22528);
  nor U24018(n22639,n22646,n22530);
  nor U24019(n22618,n22647,n22648,n22649,n22650);
  nor U24020(n22650,n22651,n22536);
  nor U24021(n22649,n22652,n22538);
  nor U24022(n22648,n22653,n22540);
  nor U24023(n22647,n22654,n22542);
  nand U24024(n22606,G59596,n22436);
  nand U24025(n22596,n22567,n22655);
  nand U24026(G8538,n22656,n22657,n22658,n22659);
  nor U24027(n22659,n22660,n22661,n22662);
  nor U24028(n22662,n21217,n22401);
  nor U24029(n22661,n22663,n22394);
  nor U24030(n22660,n22664,n22456);
  nand U24031(n22658,n22402,n21218);
  nand U24032(n22657,n22403,n21219);
  xor U24033(n21219,n22665,n22583);
  nand U24034(n22583,n22666,n22667,n22668,n22669);
  nor U24035(n22669,n22670,n22671);
  nor U24036(n22671,n22470,n22664);
  nor U24037(n22670,n22199,n22414);
  nand U24038(n22668,n22439,G59786);
  nand U24039(n22667,n21580,n22477);
  nand U24040(n22666,n22476,n22473,n21216);
  xnor U24041(n22665,n22414,n22582);
  nand U24042(n22582,n22672,n22673);
  nand U24043(n22673,n22406,n22674);
  or U24044(n22674,n22675,n22676);
  nand U24045(n22672,n22676,n22675);
  nand U24046(n22656,n22440,n21580);
  not U24047(n21580,n21216);
  xnor U24048(n21216,n22593,n22594);
  xor U24049(n22594,n22677,n22383);
  nand U24050(n22677,n22678,n22679,n22680,n22681);
  nor U24051(n22681,n22682,n22683);
  nor U24052(n22683,n22382,n21215);
  not U24053(n21215,G59627);
  nor U24054(n22682,n22167,n21217);
  not U24055(n21217,G59786);
  nand U24056(n22680,G59595,n22496);
  nand U24057(n22679,n21218,n22497);
  not U24058(n21218,n22199);
  nand U24059(n22199,n22604,n22684);
  nand U24060(n22684,n22685,n22686);
  nand U24061(n22686,n22687,n22688);
  nand U24062(n22604,n22688,n22687,n22689);
  not U24063(n22689,n22685);
  xor U24064(n22685,n22690,n22167);
  nand U24065(n22690,n22691,n22692,n22693,n22694);
  nor U24066(n22694,n22695,n22696);
  and U24067(n22696,n22437,G59722);
  nor U24068(n22695,n22508,n22664);
  nand U24069(n22693,G59627,n22435);
  or U24070(n22692,n22663,n21114);
  nand U24071(n22663,n22615,n22697);
  nand U24072(n22697,n22698,n22699);
  or U24073(n22615,n22699,n22698);
  nand U24074(n22698,n22700,n22701);
  nand U24075(n22701,n21058,n22664);
  not U24076(n22664,G59595);
  nand U24077(n22700,n22702,n22703,n22704,n21846);
  nor U24078(n22704,n22705,n22706);
  nand U24079(n22706,n22707,n22708,n22709,n22710);
  nand U24080(n22710,n22627,G59551);
  nand U24081(n22709,n22628,G59543);
  nand U24082(n22708,n22629,G59535);
  nand U24083(n22707,n22630,G59527);
  nand U24084(n22705,n22711,n22712,n22713,n22714);
  nand U24085(n22714,n22635,G59519);
  nand U24086(n22713,n22636,G59511);
  nand U24087(n22712,n22637,G59503);
  nand U24088(n22711,n22638,G59495);
  nor U24089(n22703,n22715,n22716,n22717,n22718);
  nor U24090(n22718,n22719,n22524);
  nor U24091(n22717,n22720,n22526);
  nor U24092(n22716,n22721,n22528);
  nor U24093(n22715,n22722,n22530);
  nor U24094(n22702,n22723,n22724,n22725,n22726);
  nor U24095(n22726,n22727,n22536);
  nor U24096(n22725,n22728,n22538);
  nor U24097(n22724,n22729,n22540);
  nor U24098(n22723,n22730,n22542);
  nand U24099(n22691,G59754,n22434);
  nand U24100(n22678,n22567,n22731);
  nand U24101(G8537,n22732,n22733,n22734,n22735);
  nor U24102(n22735,n22736,n22737,n22738);
  nor U24103(n22738,n21229,n22401);
  nor U24104(n22737,n22739,n22394);
  nor U24105(n22736,n22740,n22456);
  nand U24106(n22734,n22402,n21230);
  nand U24107(n22733,n22403,n21231);
  xor U24108(n21231,n22741,n22676);
  nand U24109(n22676,n22742,n22743,n22744,n22745);
  nor U24110(n22745,n22746,n22747);
  nor U24111(n22747,n21229,n22469);
  nor U24112(n22746,n22470,n22740);
  nand U24113(n22744,n22406,n21230);
  nand U24114(n22743,n21588,n22748,n22473,n22749);
  nand U24115(n22742,n21584,n22477);
  nand U24116(n22477,n22750,n22751);
  nand U24117(n22751,n22473,n22749);
  not U24118(n22749,n22476);
  nor U24119(n22476,n21240,n22752,n21228);
  xnor U24120(n22741,n22414,n22675);
  nand U24121(n22675,n22753,n22754);
  nand U24122(n22754,n22406,n22755);
  or U24123(n22755,n22756,n22757);
  nand U24124(n22753,n22757,n22756);
  nand U24125(n22732,n22440,n21584);
  not U24126(n21584,n21228);
  nand U24127(n21228,n22758,n22593);
  or U24128(n22593,n22759,n22760);
  nand U24129(n22758,n22760,n22759);
  or U24130(n22759,n22761,n22762,n22763);
  xor U24131(n22760,n22764,n22383);
  nand U24132(n22764,n22765,n22766,n22767,n22768);
  nor U24133(n22768,n22769,n22770);
  nor U24134(n22770,n22382,n21227);
  not U24135(n21227,G59626);
  nor U24136(n22769,n22167,n21229);
  not U24137(n21229,G59785);
  nand U24138(n22767,G59594,n22496);
  nand U24139(n22766,n21230,n22497);
  xor U24140(n21230,n22687,n22688);
  xnor U24141(n22688,n22771,n22167);
  nand U24142(n22771,n22772,n22773,n22774,n22775);
  nor U24143(n22775,n22776,n22777);
  and U24144(n22777,n22437,G59721);
  nor U24145(n22776,n22508,n22740);
  nand U24146(n22774,G59626,n22435);
  or U24147(n22773,n22739,n21114);
  nand U24148(n22739,n22699,n22778);
  nand U24149(n22778,n22779,n22780);
  or U24150(n22699,n22780,n22779);
  nand U24151(n22779,n22781,n22782);
  nand U24152(n22782,n21058,n22740);
  not U24153(n22740,G59594);
  nand U24154(n22781,n22783,n22784,n22785,n21846);
  nor U24155(n22785,n22786,n22787);
  nand U24156(n22787,n22788,n22789,n22790,n22791);
  nand U24157(n22791,n22627,G59552);
  nand U24158(n22790,n22628,G59544);
  nand U24159(n22789,n22629,G59536);
  nand U24160(n22788,n22630,G59528);
  nand U24161(n22786,n22792,n22793,n22794,n22795);
  nand U24162(n22795,n22635,G59520);
  nand U24163(n22794,n22636,G59512);
  nand U24164(n22793,n22637,G59504);
  nand U24165(n22792,n22638,G59496);
  nor U24166(n22784,n22796,n22797,n22798,n22799);
  nor U24167(n22799,n22800,n22524);
  nor U24168(n22798,n22801,n22526);
  nor U24169(n22797,n22802,n22528);
  nor U24170(n22796,n22803,n22530);
  nor U24171(n22783,n22804,n22805,n22806,n22807);
  nor U24172(n22807,n22808,n22536);
  nor U24173(n22806,n22809,n22538);
  nor U24174(n22805,n22810,n22540);
  nor U24175(n22804,n22811,n22542);
  nand U24176(n22772,G59753,n22434);
  and U24177(n22687,n22812,n22813);
  nand U24178(n22765,n22567,n22814);
  nand U24179(G8536,n22815,n22816,n22817,n22818);
  nor U24180(n22818,n22819,n22820,n22821);
  nor U24181(n22821,n21241,n22401);
  nor U24182(n22820,n22822,n22394);
  nor U24183(n22819,n22823,n22456);
  nand U24184(n22817,n22402,n21242);
  nand U24185(n22816,n22403,n21243);
  xor U24186(n21243,n22824,n22757);
  nand U24187(n22757,n22825,n22826,n22827,n22828);
  nor U24188(n22828,n22829,n22830);
  nor U24189(n22830,n22470,n22823);
  nor U24190(n22829,n22213,n22414);
  nand U24191(n22827,n22439,G59784);
  nand U24192(n22826,n21588,n22831);
  nand U24193(n22825,n22748,n22473,n21240);
  not U24194(n22748,n22752);
  xnor U24195(n22824,n22414,n22756);
  nand U24196(n22756,n22832,n22833);
  nand U24197(n22833,n22406,n22834);
  or U24198(n22834,n22835,n22836);
  nand U24199(n22832,n22836,n22835);
  nand U24200(n22815,n22440,n21588);
  not U24201(n21588,n21240);
  xor U24202(n21240,n22762,n22837);
  nor U24203(n22837,n22761,n22763);
  xnor U24204(n22762,n22838,n22435);
  nand U24205(n22838,n22839,n22840,n22841,n22842);
  nor U24206(n22842,n22843,n22844);
  nor U24207(n22844,n22382,n21239);
  not U24208(n21239,G59625);
  nor U24209(n22843,n22167,n21241);
  not U24210(n21241,G59784);
  nand U24211(n22841,G59593,n22496);
  nand U24212(n22840,n21242,n22497);
  not U24213(n21242,n22213);
  xnor U24214(n22213,n22813,n22812);
  xnor U24215(n22813,n22845,n22167);
  nand U24216(n22845,n22846,n22847,n22848,n22849);
  nor U24217(n22849,n22850,n22851);
  and U24218(n22851,n22437,G59720);
  nor U24219(n22850,n22508,n22823);
  nand U24220(n22848,G59625,n22435);
  or U24221(n22847,n22822,n21114);
  nand U24222(n22822,n22780,n22852);
  nand U24223(n22852,n22853,n22854);
  or U24224(n22780,n22854,n22853);
  nand U24225(n22853,n22855,n22856);
  nand U24226(n22856,n21058,n22823);
  not U24227(n22823,G59593);
  nand U24228(n22855,n22857,n22858,n22859,n21846);
  nor U24229(n22859,n22860,n22861);
  nand U24230(n22861,n22862,n22863,n22864,n22865);
  nand U24231(n22865,n22627,G59553);
  nand U24232(n22864,n22628,G59545);
  nand U24233(n22863,n22629,G59537);
  nand U24234(n22862,n22630,G59529);
  nand U24235(n22860,n22866,n22867,n22868,n22869);
  nand U24236(n22869,n22635,G59521);
  nand U24237(n22868,n22636,G59513);
  nand U24238(n22867,n22637,G59505);
  nand U24239(n22866,n22638,G59497);
  nor U24240(n22858,n22870,n22871,n22872,n22873);
  nor U24241(n22873,n22874,n22524);
  nor U24242(n22872,n22875,n22526);
  nor U24243(n22871,n22876,n22528);
  nor U24244(n22870,n22877,n22530);
  nor U24245(n22857,n22878,n22879,n22880,n22881);
  nor U24246(n22881,n22882,n22536);
  nor U24247(n22880,n22883,n22538);
  nor U24248(n22879,n22884,n22540);
  nor U24249(n22878,n22885,n22542);
  nand U24250(n22846,G59752,n22434);
  nand U24251(n22839,n22567,n22886);
  nand U24252(G8535,n22887,n22888,n22889,n22890);
  nor U24253(n22890,n22891,n22892,n22893);
  nor U24254(n22893,n21253,n22401);
  nor U24255(n22892,n22894,n22394);
  nor U24256(n22891,n22895,n22456);
  nand U24257(n22889,n22402,n21254);
  nand U24258(n22888,n22403,n21255);
  xor U24259(n21255,n22896,n22836);
  nand U24260(n22836,n22897,n22898,n22899,n22900);
  nor U24261(n22900,n22901,n22902);
  nor U24262(n22902,n21253,n22469);
  nor U24263(n22901,n22470,n22895);
  nand U24264(n22899,n22406,n21254);
  nand U24265(n22898,n21595,n22752,n22903);
  nand U24266(n22897,n21252,n22831);
  nand U24267(n22831,n22750,n22904);
  nand U24268(n22904,n22473,n22752);
  nand U24269(n22752,n22905,n21595,n21252,n21599);
  xnor U24270(n22896,n22414,n22835);
  nand U24271(n22835,n22906,n22907);
  nand U24272(n22907,n22406,n22908);
  or U24273(n22908,n22909,n22910);
  nand U24274(n22906,n22910,n22909);
  nand U24275(n22887,n22440,n21252);
  xor U24276(n21252,n22763,n22761);
  xor U24277(n22761,n22911,n22383);
  nand U24278(n22911,n22912,n22913,n22914,n22915);
  nor U24279(n22915,n22916,n22917);
  nor U24280(n22917,n22382,n21251);
  not U24281(n21251,G59624);
  nor U24282(n22916,n22167,n21253);
  not U24283(n21253,G59783);
  nand U24284(n22914,G59592,n22496);
  nand U24285(n22913,n21254,n22497);
  nor U24286(n21254,n22918,n22812);
  nor U24287(n22812,n22919,n22920);
  and U24288(n22918,n22920,n22919);
  nand U24289(n22919,n22921,n22922,n22923);
  xor U24290(n22920,n22924,n22167);
  nand U24291(n22924,n22925,n22926,n22927,n22928);
  nor U24292(n22928,n22929,n22930);
  and U24293(n22930,n22437,G59719);
  nor U24294(n22929,n22508,n22895);
  nand U24295(n22927,G59624,n22435);
  or U24296(n22926,n22894,n21114);
  nand U24297(n22894,n22854,n22931);
  nand U24298(n22931,n22932,n22933);
  or U24299(n22854,n22933,n22932);
  nand U24300(n22932,n22934,n22935);
  nand U24301(n22935,n21058,n22895);
  not U24302(n22895,G59592);
  nand U24303(n22934,n22936,n22937,n22938,n21846);
  nor U24304(n22938,n22939,n22940);
  nand U24305(n22940,n22941,n22942,n22943,n22944);
  nand U24306(n22944,n22627,G59554);
  not U24307(n22627,n22566);
  nand U24308(n22943,n22628,G59546);
  not U24309(n22628,n22564);
  nand U24310(n22942,n22629,G59538);
  not U24311(n22629,n22562);
  nand U24312(n22941,n22630,G59530);
  not U24313(n22630,n22560);
  nand U24314(n22939,n22945,n22946,n22947,n22948);
  nand U24315(n22948,n22635,G59522);
  not U24316(n22635,n22554);
  nand U24317(n22947,n22636,G59514);
  not U24318(n22636,n22552);
  nand U24319(n22946,n22637,G59506);
  not U24320(n22637,n22550);
  nand U24321(n22945,n22638,G59498);
  not U24322(n22638,n22548);
  nor U24323(n22937,n22949,n22950,n22951,n22952);
  nor U24324(n22952,n22953,n22524);
  nor U24325(n22951,n22954,n22526);
  nor U24326(n22950,n22955,n22528);
  nor U24327(n22949,n22956,n22530);
  nor U24328(n22936,n22957,n22958,n22959,n22960);
  nor U24329(n22960,n22961,n22536);
  nor U24330(n22959,n22962,n22538);
  nor U24331(n22958,n22963,n22540);
  nor U24332(n22957,n22964,n22542);
  nand U24333(n22933,n22965,n22966);
  nand U24334(n22925,G59751,n22434);
  nand U24335(n22912,n22567,n22967);
  nand U24336(G8534,n22968,n22969,n22970,n22971);
  nor U24337(n22971,n22972,n22973,n22974);
  nor U24338(n22974,n21265,n22401);
  nor U24339(n22973,n22226,n22975);
  nor U24340(n22972,n22976,n22456);
  nand U24341(n22970,n22440,n21595);
  nand U24342(n22969,n22400,n22977);
  nand U24343(n22968,n22403,n21267);
  xor U24344(n21267,n22978,n22910);
  nand U24345(n22910,n22979,n22980,n22981,n22982);
  nor U24346(n22982,n22983,n22984);
  nor U24347(n22984,n22470,n22976);
  nor U24348(n22983,n22226,n22414);
  not U24349(n22226,n21266);
  nand U24350(n22981,n22439,G59782);
  nand U24351(n22980,n22903,n21264);
  nor U24352(n22903,n21276,n21935,n22985);
  nand U24353(n22979,n21595,n22986);
  nand U24354(n22986,n22987,n22988);
  nand U24355(n22988,n22473,n21276);
  not U24356(n22987,n22989);
  not U24357(n21595,n21264);
  nand U24358(n21264,n22763,n22990);
  nand U24359(n22990,n22991,n22992);
  or U24360(n22763,n22992,n22991);
  and U24361(n22991,n22993,n22994);
  nand U24362(n22993,n22995,n22996);
  xor U24363(n22992,n22997,n22383);
  nand U24364(n22997,n22998,n22999,n23000,n23001);
  nor U24365(n23001,n23002,n23003);
  nor U24366(n23003,n22382,n21263);
  not U24367(n21263,G59623);
  nor U24368(n23002,n22167,n21265);
  not U24369(n21265,G59782);
  nand U24370(n23000,G59591,n22496);
  nand U24371(n22999,n21266,n22497);
  xnor U24372(n21266,n23004,n22923);
  xor U24373(n22923,n23005,n21108);
  nand U24374(n23005,n23006,n23007,n23008,n23009);
  nor U24375(n23009,n23010,n23011);
  and U24376(n23011,n22437,G59718);
  nor U24377(n23010,n22508,n22976);
  not U24378(n22976,G59591);
  nand U24379(n23008,G59623,n22435);
  nand U24380(n23007,n21691,n22977);
  xor U24381(n22977,n22965,n22966);
  nand U24382(n22966,n23012,n23013);
  nand U24383(n23013,G59591,n21058);
  nand U24384(n23012,n23014,n21846);
  nand U24385(n23014,n23015,n23016,n23017,n23018);
  nor U24386(n23018,n23019,n23020,n23021,n23022);
  nor U24387(n23022,n23023,n22524);
  nor U24388(n23021,n23024,n22526);
  nor U24389(n23020,n23025,n22528);
  nor U24390(n23019,n23026,n22530);
  nor U24391(n23017,n23027,n23028,n23029,n23030);
  nor U24392(n23030,n23031,n22536);
  nor U24393(n23029,n23032,n22538);
  nor U24394(n23028,n23033,n22540);
  nor U24395(n23027,n23034,n22542);
  nor U24396(n23016,n23035,n23036,n23037,n23038);
  nor U24397(n23038,n23039,n22548);
  nor U24398(n23037,n23040,n22550);
  nor U24399(n23036,n23041,n22552);
  nor U24400(n23035,n23042,n22554);
  nor U24401(n23015,n23043,n23044,n23045,n23046);
  nor U24402(n23046,n23047,n22560);
  nor U24403(n23045,n23048,n22562);
  nor U24404(n23044,n23049,n22564);
  nor U24405(n23043,n23050,n22566);
  and U24406(n22965,n23051,n23052);
  nand U24407(n23006,G59750,n22434);
  nand U24408(n23004,n22922,n22921);
  nand U24409(n22998,n22567,n23053);
  xnor U24410(n22978,n22414,n22909);
  nand U24411(n22909,n23054,n23055);
  nand U24412(n23055,n22406,n23056);
  or U24413(n23056,n23057,n23058);
  nand U24414(n23054,n23058,n23057);
  nand U24415(G8533,n23059,n23060,n23061,n23062);
  nor U24416(n23062,n23063,n23064,n23065);
  nor U24417(n23065,n21277,n22401);
  nor U24418(n23064,n21786,n22975);
  nor U24419(n23063,n23066,n22456);
  nand U24420(n23061,n22440,n21599);
  nand U24421(n23060,n22400,n23067);
  nand U24422(n23059,n22403,n21279);
  xor U24423(n21279,n23068,n23058);
  nand U24424(n23058,n23069,n23070,n23071,n23072);
  nor U24425(n23072,n23073,n23074);
  nor U24426(n23074,n22470,n23066);
  nor U24427(n23073,n21786,n22414);
  not U24428(n21786,n21278);
  nand U24429(n23071,n22439,G59781);
  nand U24430(n23070,n21599,n22989);
  not U24431(n21599,n21276);
  nand U24432(n23069,n22905,n22473,n21276);
  xnor U24433(n21276,n22995,n23075);
  and U24434(n23075,n22994,n22996);
  nand U24435(n22996,n23076,n23077,n23078);
  nand U24436(n23078,n22567,n23079);
  nand U24437(n22994,n23080,n23079,n22567);
  nand U24438(n23080,n23076,n23077);
  or U24439(n23077,n23081,n22383);
  nand U24440(n23076,n22383,n23081);
  nand U24441(n23081,n23082,n23083,n23084,n23085);
  nor U24442(n23085,n23086,n23087);
  nor U24443(n23087,n22382,n21275);
  not U24444(n21275,G59622);
  nor U24445(n23086,n22167,n21277);
  not U24446(n21277,G59781);
  nand U24447(n23084,G59590,n22496);
  nand U24448(n23083,n21278,n22497);
  xor U24449(n21278,n22921,n22922);
  xnor U24450(n22921,n23088,n22167);
  nand U24451(n23088,n23089,n23090,n23091,n23092);
  nor U24452(n23092,n23093,n23094);
  and U24453(n23094,n22437,G59717);
  nor U24454(n23093,n22508,n23066);
  not U24455(n23066,G59590);
  nand U24456(n23091,G59622,n22435);
  nand U24457(n23090,n21691,n23067);
  xor U24458(n23067,n23052,n23051);
  nand U24459(n23051,n23095,n23096);
  nand U24460(n23096,G59590,n21058);
  nand U24461(n23095,n23097,n21846);
  nand U24462(n23097,n23098,n23099,n23100,n23101);
  nor U24463(n23101,n23102,n23103,n23104,n23105);
  nor U24464(n23105,n23106,n22524);
  nand U24465(n22524,n23107,n23108);
  nor U24466(n23104,n23109,n22526);
  nand U24467(n22526,n23110,n23108);
  nor U24468(n23103,n23111,n22528);
  nand U24469(n22528,n23112,n23108);
  nor U24470(n23102,n23113,n22530);
  nand U24471(n22530,n23114,n23108);
  and U24472(n23108,n23115,n23116);
  nor U24473(n23100,n23117,n23118,n23119,n23120);
  nor U24474(n23120,n23121,n22536);
  nand U24475(n22536,n23122,n23107);
  nor U24476(n23119,n23123,n22538);
  nand U24477(n22538,n23122,n23110);
  nor U24478(n23118,n23124,n22540);
  nand U24479(n22540,n23122,n23112);
  nor U24480(n23117,n23125,n22542);
  nand U24481(n22542,n23122,n23114);
  and U24482(n23122,n23126,n23116);
  nor U24483(n23099,n23127,n23128,n23129,n23130);
  nor U24484(n23130,n23131,n22548);
  nand U24485(n22548,n23132,n23107);
  nor U24486(n23129,n23133,n22550);
  nand U24487(n22550,n23132,n23110);
  nor U24488(n23128,n23134,n22552);
  nand U24489(n22552,n23132,n23112);
  nor U24490(n23127,n23135,n22554);
  nand U24491(n22554,n23132,n23114);
  nor U24492(n23132,n23116,n23126);
  not U24493(n23126,n23115);
  nor U24494(n23098,n23136,n23137,n23138,n23139);
  nor U24495(n23139,n23140,n22560);
  nand U24496(n22560,n23141,n23107);
  nor U24497(n23107,n23142,n23143);
  nor U24498(n23138,n23144,n22562);
  nand U24499(n22562,n23141,n23110);
  nor U24500(n23110,G59561,n23143);
  nor U24501(n23137,n23145,n22564);
  nand U24502(n22564,n23141,n23112);
  nor U24503(n23112,n23146,n23142);
  nor U24504(n23136,n23147,n22566);
  nand U24505(n22566,n23141,n23114);
  nor U24506(n23114,n23146,G59561);
  nor U24507(n23141,n23116,n23115);
  nand U24508(n23052,n23148,n23149);
  nand U24509(n23149,n23150,G59589);
  nand U24510(n23148,n21846,n22568);
  nand U24511(n22568,n23151,n23152,n23153,n23154);
  nor U24512(n23154,n23155,n23156,n23157,n23158);
  nor U24513(n23158,n22525,n23159);
  nor U24514(n23157,n22527,n23160);
  nor U24515(n23156,n22539,n23161);
  nor U24516(n23155,n22551,n23162);
  nor U24517(n23153,n23163,n23164,n23165,n23166);
  nor U24518(n23166,n22537,n23167);
  nor U24519(n23165,n22541,n23168);
  nor U24520(n23164,n22565,n23169);
  nor U24521(n23163,n22523,n23170);
  nor U24522(n23152,n23171,n23172,n23173,n23174);
  nor U24523(n23174,n22549,n23175);
  nor U24524(n23173,n22553,n23176);
  nor U24525(n23172,n22559,n23177);
  nor U24526(n23171,n22535,n23178);
  nor U24527(n23151,n23179,n23180,n23181,n23182);
  nor U24528(n23182,n22563,n23183);
  nor U24529(n23181,n22561,n23184);
  nor U24530(n23180,n22547,n23185);
  nor U24531(n23179,n22529,n23186);
  nand U24532(n23089,G59749,n22434);
  nand U24533(n23082,n22567,n23187);
  nand U24534(n22995,n23188,n23189);
  nand U24535(n23189,n23190,n23191);
  not U24536(n22905,n22985);
  xnor U24537(n23068,n22414,n23057);
  nand U24538(n23057,n23192,n23193);
  nand U24539(n23193,n22406,n23194);
  or U24540(n23194,n23195,n23196);
  nand U24541(n23192,n23196,n23195);
  nand U24542(G8532,n23197,n23198,n23199,n23200);
  nor U24543(n23200,n23201,n23202,n23203);
  nor U24544(n23203,n21289,n22401);
  and U24545(n23202,n23204,n22400);
  nor U24546(n23201,n23205,n22456);
  nand U24547(n23199,n22402,n21290);
  nand U24548(n23198,n22403,n21291);
  xor U24549(n21291,n23206,n23196);
  nand U24550(n23196,n23207,n23208,n23209,n23210);
  nor U24551(n23210,n23211,n23212);
  nor U24552(n23212,n21289,n22469);
  not U24553(n21289,G59780);
  nor U24554(n23211,n22470,n23205);
  nand U24555(n23209,n22406,n21290);
  nand U24556(n23208,n21606,n22985,n23213);
  nand U24557(n23207,n21288,n22989);
  nand U24558(n22989,n22750,n23214);
  nand U24559(n23214,n22473,n22985);
  nand U24560(n22985,n21288,n23215,n21606,n21610);
  xnor U24561(n23206,n22414,n23195);
  nand U24562(n23195,n23216,n23217);
  nand U24563(n23217,n22406,n23218);
  or U24564(n23218,n23219,n23220);
  nand U24565(n23216,n23220,n23219);
  nand U24566(n23197,n22440,n21288);
  xor U24567(n21288,n23191,n23221);
  and U24568(n23221,n23188,n23190);
  nand U24569(n23190,n23222,n23223,n23224);
  nand U24570(n23224,n22567,n23225);
  nand U24571(n23188,n23226,n23225,n22567);
  nand U24572(n23226,n23222,n23223);
  nand U24573(n23223,n22435,n21796,n23227);
  not U24574(n21796,n21290);
  nand U24575(n23222,n23228,n22383);
  nand U24576(n23228,n23227,n23229);
  nand U24577(n23229,n21290,n22497);
  nor U24578(n21290,n23230,n22922);
  nor U24579(n22922,n23231,n23232,n23233);
  and U24580(n23230,n23231,n23234);
  or U24581(n23234,n23233,n23232);
  xor U24582(n23231,n21108,n23235);
  nor U24583(n23235,n23236,n23237,n23238);
  and U24584(n23238,n22437,G59716);
  nor U24585(n23237,n22508,n23205);
  nand U24586(n23236,n23239,n23240,n23241);
  nand U24587(n23241,G59621,n22435);
  nand U24588(n23240,n21691,n23204);
  nand U24589(n23204,n23242,n23243,n23244);
  nand U24590(n23244,n23150,n23205);
  not U24591(n23205,G59589);
  not U24592(n23150,n23245);
  nand U24593(n23243,G59589,n23245,n21058);
  nand U24594(n23245,G59588,n23246);
  nand U24595(n23242,n22655,n21846);
  nand U24596(n22655,n23247,n23248,n23249,n23250);
  nor U24597(n23250,n23251,n23252,n23253,n23254);
  nor U24598(n23254,n23255,n23177);
  nor U24599(n23253,n23256,n23184);
  nor U24600(n23252,n23257,n23183);
  nor U24601(n23251,n23258,n23169);
  nor U24602(n23249,n23259,n23260,n23261,n23262);
  nor U24603(n23262,n23263,n23185);
  nor U24604(n23261,n23264,n23175);
  nor U24605(n23260,n23265,n23162);
  nor U24606(n23259,n23266,n23176);
  nor U24607(n23248,n23267,n23268,n23269,n23270);
  nor U24608(n23270,n22651,n23178);
  nor U24609(n23269,n22652,n23167);
  nor U24610(n23268,n22653,n23161);
  nor U24611(n23267,n22654,n23168);
  nor U24612(n23247,n23271,n23272,n23273,n23274);
  nor U24613(n23274,n22643,n23170);
  nor U24614(n23273,n22644,n23159);
  nor U24615(n23272,n22645,n23160);
  nor U24616(n23271,n22646,n23186);
  nand U24617(n23239,G59748,n22434);
  and U24618(n23227,n23275,n23276,n23277);
  nand U24619(n23277,G59621,n23278);
  nand U24620(n23276,G59589,n22496);
  nand U24621(n23275,G59780,n21108);
  nand U24622(n23191,n23279,n23280);
  nand U24623(n23280,n23281,n23282);
  nand U24624(G8531,n23283,n23284,n23285,n23286);
  nor U24625(n23286,n23287,n23288,n23289);
  nor U24626(n23289,n21301,n22401);
  not U24627(n21301,G59779);
  and U24628(n23288,n23290,n22400);
  nor U24629(n23287,n23291,n22456);
  nand U24630(n23285,n22402,n21302);
  nand U24631(n23284,n22403,n21303);
  xor U24632(n21303,n23292,n23220);
  nand U24633(n23220,n23293,n23294,n23295,n23296);
  nor U24634(n23296,n23297,n23298);
  nor U24635(n23298,n22470,n23291);
  nor U24636(n23297,n21805,n22414);
  nand U24637(n23295,n22439,G59779);
  nand U24638(n23294,n21300,n23213);
  nor U24639(n23213,n21312,n21935,n23299);
  nand U24640(n23293,n21606,n23300);
  nand U24641(n23300,n23301,n23302);
  nand U24642(n23302,n22473,n21312);
  not U24643(n23301,n23303);
  xnor U24644(n23292,n22414,n23219);
  nand U24645(n23219,n23304,n23305);
  nand U24646(n23305,n22406,n23306);
  or U24647(n23306,n23307,n23308);
  nand U24648(n23304,n23308,n23307);
  nand U24649(n23283,n22440,n21606);
  not U24650(n21606,n21300);
  xnor U24651(n21300,n23282,n23309);
  and U24652(n23309,n23279,n23281);
  nand U24653(n23281,n23310,n23311,n23312);
  nand U24654(n23312,n22567,n23313);
  nand U24655(n23279,n23314,n23313,n22567);
  nand U24656(n23314,n23310,n23311);
  nand U24657(n23311,n22435,n21805,n23315);
  nand U24658(n23310,n23316,n22383);
  nand U24659(n23316,n23315,n23317);
  nand U24660(n23317,n21302,n22497);
  not U24661(n21302,n21805);
  xnor U24662(n21805,n23233,n23232);
  xor U24663(n23232,n21108,n23318);
  nor U24664(n23318,n23319,n23320,n23321);
  and U24665(n23321,n22437,G59715);
  nor U24666(n23320,n22508,n23291);
  nand U24667(n23319,n23322,n23323,n23324);
  nand U24668(n23324,G59620,n22435);
  nand U24669(n23323,n21691,n23290);
  nand U24670(n23290,n23325,n23326);
  nand U24671(n23326,n22731,n21846);
  nand U24672(n22731,n23327,n23328,n23329,n23330);
  nor U24673(n23330,n23331,n23332,n23333,n23334);
  nor U24674(n23334,n23335,n23177);
  nor U24675(n23333,n23336,n23184);
  nor U24676(n23332,n23337,n23183);
  nor U24677(n23331,n23338,n23169);
  nor U24678(n23329,n23339,n23340,n23341,n23342);
  nor U24679(n23342,n23343,n23185);
  nor U24680(n23341,n23344,n23175);
  nor U24681(n23340,n23345,n23162);
  nor U24682(n23339,n23346,n23176);
  nor U24683(n23328,n23347,n23348,n23349,n23350);
  nor U24684(n23350,n22727,n23178);
  nor U24685(n23349,n22728,n23167);
  nor U24686(n23348,n22729,n23161);
  nor U24687(n23347,n22730,n23168);
  nor U24688(n23327,n23351,n23352,n23353,n23354);
  nor U24689(n23354,n22719,n23170);
  nor U24690(n23353,n22720,n23159);
  nor U24691(n23352,n22721,n23160);
  nor U24692(n23351,n22722,n23186);
  nand U24693(n23325,n23355,n21058);
  xnor U24694(n23355,n23291,n23246);
  nor U24695(n23246,n23356,n23357);
  not U24696(n23291,G59588);
  nand U24697(n23322,G59747,n22434);
  and U24698(n23315,n23358,n23359,n23360);
  nand U24699(n23360,G59620,n23278);
  nand U24700(n23359,G59588,n22496);
  nand U24701(n23358,G59779,n21108);
  nand U24702(n23282,n23361,n23362);
  nand U24703(n23362,n23363,n23364);
  nand U24704(G8530,n23365,n23366,n23367,n23368);
  nor U24705(n23368,n23369,n23370,n23371);
  nor U24706(n23371,n21313,n22401);
  not U24707(n21313,G59778);
  and U24708(n23370,n23372,n22400);
  nor U24709(n23369,n23357,n22456);
  nand U24710(n23367,n22402,n21314);
  nand U24711(n23366,n22403,n21315);
  xor U24712(n21315,n23373,n23308);
  nand U24713(n23308,n23374,n23375,n23376,n23377);
  nor U24714(n23377,n23378,n23379);
  nor U24715(n23379,n22470,n23357);
  nor U24716(n23378,n21814,n22414);
  nand U24717(n23376,n22439,G59778);
  nand U24718(n23375,n21610,n23303);
  nand U24719(n23374,n23215,n22473,n21312);
  not U24720(n23215,n23299);
  xnor U24721(n23373,n22414,n23307);
  nand U24722(n23307,n23380,n23381);
  nand U24723(n23381,n22406,n23382);
  or U24724(n23382,n23383,n23384);
  nand U24725(n23380,n23384,n23383);
  nand U24726(n23365,n22440,n21610);
  not U24727(n21610,n21312);
  xnor U24728(n21312,n23364,n23385);
  and U24729(n23385,n23361,n23363);
  nand U24730(n23363,n23386,n23387,n23388);
  nand U24731(n23361,n23390,n23389,n22567);
  nand U24732(n23390,n23386,n23387);
  nand U24733(n23387,n22435,n21814,n23391);
  nand U24734(n23386,n23392,n22383);
  nand U24735(n23392,n23391,n23393);
  nand U24736(n23393,n21314,n22497);
  not U24737(n21314,n21814);
  nand U24738(n21814,n23233,n23394);
  nand U24739(n23394,n23395,n23396);
  or U24740(n23233,n23396,n23395);
  xor U24741(n23395,n21108,n23397);
  nor U24742(n23397,n23398,n23399,n23400);
  and U24743(n23400,n22437,G59714);
  nor U24744(n23399,n22508,n23357);
  not U24745(n23357,G59587);
  nand U24746(n23398,n23401,n23402,n23403);
  nand U24747(n23403,G59619,n22435);
  nand U24748(n23402,n21691,n23372);
  nand U24749(n23372,n23404,n23405,n23406);
  or U24750(n23406,n23356,G59587);
  nand U24751(n23405,G59587,n23356,n21058);
  nand U24752(n23356,n23407,G59586);
  nand U24753(n23404,n22814,n21846);
  nand U24754(n22814,n23408,n23409,n23410,n23411);
  nor U24755(n23411,n23412,n23413,n23414,n23415);
  nor U24756(n23415,n23416,n23177);
  nor U24757(n23414,n23417,n23184);
  nor U24758(n23413,n23418,n23183);
  nor U24759(n23412,n23419,n23169);
  nor U24760(n23410,n23420,n23421,n23422,n23423);
  nor U24761(n23423,n23424,n23185);
  nor U24762(n23422,n23425,n23175);
  nor U24763(n23421,n23426,n23162);
  nor U24764(n23420,n23427,n23176);
  nor U24765(n23409,n23428,n23429,n23430,n23431);
  nor U24766(n23431,n22808,n23178);
  nor U24767(n23430,n22809,n23167);
  nor U24768(n23429,n22810,n23161);
  nor U24769(n23428,n22811,n23168);
  nor U24770(n23408,n23432,n23433,n23434,n23435);
  nor U24771(n23435,n22800,n23170);
  nor U24772(n23434,n22801,n23159);
  nor U24773(n23433,n22802,n23160);
  nor U24774(n23432,n22803,n23186);
  nand U24775(n23401,G59746,n22434);
  and U24776(n23391,n23436,n23437,n23438);
  nand U24777(n23438,G59619,n23278);
  nand U24778(n23437,G59587,n22496);
  nand U24779(n23436,G59778,n21108);
  nand U24780(n23364,n23439,n23440);
  nand U24781(n23440,n23441,n23442);
  nand U24782(G8529,n23443,n23444,n23445,n23446);
  nor U24783(n23446,n23447,n23448,n23449);
  nor U24784(n23449,n23450,n22401);
  and U24785(n23448,n23451,n22400);
  nor U24786(n23447,n23452,n22456);
  nand U24787(n23445,n22402,n21614);
  nand U24788(n23444,n22403,n21326);
  xor U24789(n21326,n23453,n23384);
  nand U24790(n23384,n23454,n23455,n23456,n23457);
  nor U24791(n23457,n23458,n23459);
  nor U24792(n23459,n23450,n22469);
  not U24793(n23450,G59777);
  nor U24794(n23458,n22470,n23452);
  nand U24795(n23456,n22406,n21614);
  nand U24796(n23455,n21349,n23460,n21339,n23299);
  nand U24797(n23454,n21328,n23303);
  nand U24798(n23303,n22750,n23461);
  nand U24799(n23461,n22473,n23299);
  nand U24800(n23299,n21359,n23462,n21339,n23463);
  and U24801(n23463,n21328,n21349);
  xnor U24802(n23453,n22414,n23383);
  nand U24803(n23383,n23464,n23465);
  nand U24804(n23465,n22406,n23466);
  or U24805(n23466,n23467,n23468);
  nand U24806(n23464,n23468,n23467);
  nand U24807(n23443,n22440,n21328);
  xor U24808(n21328,n23442,n23469);
  and U24809(n23469,n23439,n23441);
  nand U24810(n23441,n23470,n23471,n23472);
  nand U24811(n23439,n23474,n23473,n22567);
  nand U24812(n23474,n23470,n23471);
  nand U24813(n23471,n22435,n21325,n23475);
  nand U24814(n23470,n23476,n22383);
  nand U24815(n23476,n23475,n23477);
  nand U24816(n23477,n21614,n22497);
  not U24817(n21614,n21325);
  nand U24818(n21325,n23478,n23396);
  or U24819(n23396,n23479,n23480,n23481);
  nand U24820(n23478,n23479,n23482);
  or U24821(n23482,n23481,n23480);
  xor U24822(n23479,n21108,n23483);
  nor U24823(n23483,n23484,n23485,n23486);
  and U24824(n23486,n22437,G59713);
  nor U24825(n23485,n22508,n23452);
  nand U24826(n23484,n23487,n23488,n23489);
  nand U24827(n23489,G59618,n22435);
  nand U24828(n23488,n21691,n23451);
  nand U24829(n23451,n23490,n23491);
  nand U24830(n23491,n22886,n21846);
  nand U24831(n22886,n23492,n23493,n23494,n23495);
  nor U24832(n23495,n23496,n23497,n23498,n23499);
  nor U24833(n23499,n23500,n23177);
  nor U24834(n23498,n23501,n23184);
  nor U24835(n23497,n23502,n23183);
  nor U24836(n23496,n23503,n23169);
  nor U24837(n23494,n23504,n23505,n23506,n23507);
  nor U24838(n23507,n23508,n23185);
  nor U24839(n23506,n23509,n23175);
  nor U24840(n23505,n23510,n23162);
  nor U24841(n23504,n23511,n23176);
  nor U24842(n23493,n23512,n23513,n23514,n23515);
  nor U24843(n23515,n22882,n23178);
  nor U24844(n23514,n22883,n23167);
  nor U24845(n23513,n22884,n23161);
  nor U24846(n23512,n22885,n23168);
  nor U24847(n23492,n23516,n23517,n23518,n23519);
  nor U24848(n23519,n22874,n23170);
  nor U24849(n23518,n22875,n23159);
  nor U24850(n23517,n22876,n23160);
  nor U24851(n23516,n22877,n23186);
  nand U24852(n23490,n23520,n21058);
  xnor U24853(n23520,n23452,n23407);
  nor U24854(n23407,n23521,n23522);
  not U24855(n23452,G59586);
  nand U24856(n23487,G59745,n22434);
  and U24857(n23475,n23523,n23524,n23525);
  nand U24858(n23525,G59618,n23278);
  nand U24859(n23524,G59586,n22496);
  nand U24860(n23523,G59777,n21108);
  nand U24861(n23442,n23526,n23527);
  nand U24862(n23527,n23528,n23529);
  nand U24863(G8528,n23530,n23531,n23532,n23533);
  nor U24864(n23533,n23534,n23535,n23536);
  nor U24865(n23536,n23537,n22401);
  not U24866(n23537,G59776);
  and U24867(n23535,n23538,n22400);
  nor U24868(n23534,n23521,n22456);
  nand U24869(n23532,n22402,n21618);
  nand U24870(n23531,n22403,n21338);
  xor U24871(n21338,n23539,n23468);
  nand U24872(n23468,n23540,n23541,n23542,n23543);
  nor U24873(n23543,n23544,n23545);
  nor U24874(n23545,n22470,n23521);
  nor U24875(n23544,n21337,n22414);
  nand U24876(n23542,n22439,G59776);
  nand U24877(n23541,n21339,n23546);
  nand U24878(n23546,n23547,n23548);
  nand U24879(n23548,n22473,n23549);
  nand U24880(n23540,n23460,n21349,n23550);
  xnor U24881(n23539,n22414,n23467);
  nand U24882(n23467,n23551,n23552);
  nand U24883(n23552,n22406,n23553);
  or U24884(n23553,n23554,n23555);
  nand U24885(n23551,n23555,n23554);
  nand U24886(n23530,n22440,n21339);
  not U24887(n21339,n23550);
  xnor U24888(n23550,n23528,n23556);
  and U24889(n23556,n23529,n23526);
  nand U24890(n23526,n23557,n23558,n22567);
  nand U24891(n23557,n23559,n23560);
  nand U24892(n23529,n23559,n23560,n23561);
  nand U24893(n23560,n22435,n21337,n23562);
  nand U24894(n23559,n23563,n22383);
  nand U24895(n23563,n23562,n23564);
  nand U24896(n23564,n21618,n22497);
  not U24897(n21618,n21337);
  xnor U24898(n21337,n23481,n23480);
  xor U24899(n23480,n21108,n23565);
  nor U24900(n23565,n23566,n23567,n23568);
  and U24901(n23568,n22437,G59712);
  nor U24902(n23567,n22508,n23521);
  not U24903(n23521,G59585);
  nand U24904(n23566,n23569,n23570,n23571);
  nand U24905(n23571,G59617,n22435);
  nand U24906(n23570,n21691,n23538);
  nand U24907(n23538,n23572,n23573,n23574);
  or U24908(n23574,n23522,G59585);
  nand U24909(n23573,G59585,n23522,n21058);
  nand U24910(n23522,n23575,n23576);
  nand U24911(n23572,n22967,n21846);
  nand U24912(n22967,n23577,n23578,n23579,n23580);
  nor U24913(n23580,n23581,n23582,n23583,n23584);
  nor U24914(n23584,n23585,n23177);
  nor U24915(n23583,n23586,n23184);
  nor U24916(n23582,n23587,n23183);
  nor U24917(n23581,n23588,n23169);
  nor U24918(n23579,n23589,n23590,n23591,n23592);
  nor U24919(n23592,n23593,n23185);
  nor U24920(n23591,n23594,n23175);
  nor U24921(n23590,n23595,n23162);
  nor U24922(n23589,n23596,n23176);
  nor U24923(n23578,n23597,n23598,n23599,n23600);
  nor U24924(n23600,n22961,n23178);
  nor U24925(n23599,n22962,n23167);
  nor U24926(n23598,n22963,n23161);
  nor U24927(n23597,n22964,n23168);
  nor U24928(n23577,n23601,n23602,n23603,n23604);
  nor U24929(n23604,n22953,n23170);
  nor U24930(n23603,n22954,n23159);
  nor U24931(n23602,n22955,n23160);
  nor U24932(n23601,n22956,n23186);
  nand U24933(n23569,G59744,n22434);
  and U24934(n23562,n23605,n23606,n23607);
  nand U24935(n23607,G59617,n23278);
  nand U24936(n23606,G59585,n22496);
  nand U24937(n23605,G59776,n21108);
  nand U24938(n23528,n23608,n23609);
  nand U24939(n23609,n23610,n23611);
  nand U24940(G8527,n23612,n23613,n23614,n23615);
  nor U24941(n23615,n23616,n23617,n23618);
  nor U24942(n23618,n23619,n22401);
  not U24943(n23619,G59775);
  and U24944(n23617,n23620,n22400);
  nor U24945(n23616,n23621,n22456);
  nand U24946(n23614,n22402,n21622);
  nand U24947(n23613,n22403,n21348);
  xor U24948(n21348,n23622,n23555);
  nand U24949(n23555,n23623,n23624,n23625,n23626);
  nor U24950(n23626,n23627,n23628);
  nor U24951(n23628,n22470,n23621);
  nor U24952(n23627,n21347,n22414);
  nand U24953(n23625,n22439,G59775);
  nand U24954(n23624,n23460,n23549);
  nor U24955(n23460,n23629,n23630,n21935);
  or U24956(n23623,n23549,n23547);
  nor U24957(n23547,n23631,n23632);
  nor U24958(n23632,n21359,n21935);
  xnor U24959(n23622,n22414,n23554);
  nand U24960(n23554,n23633,n23634);
  nand U24961(n23634,n22406,n23635);
  or U24962(n23635,n23636,n23637);
  nand U24963(n23633,n23637,n23636);
  nand U24964(n23612,n22440,n21349);
  not U24965(n21349,n23549);
  xnor U24966(n23549,n23610,n23638);
  and U24967(n23638,n23611,n23608);
  nand U24968(n23608,n23639,n23640,n22567);
  nand U24969(n23639,n23641,n23642);
  nand U24970(n23611,n23641,n23642,n23643);
  nand U24971(n23642,n22435,n21347,n23644);
  nand U24972(n23641,n23645,n22383);
  nand U24973(n23645,n23644,n23646);
  nand U24974(n23646,n21622,n22497);
  not U24975(n21622,n21347);
  nand U24976(n21347,n23481,n23647);
  nand U24977(n23647,n23648,n23649);
  or U24978(n23481,n23649,n23648);
  xor U24979(n23648,n21108,n23650);
  nor U24980(n23650,n23651,n23652,n23653);
  and U24981(n23653,n22437,G59711);
  nor U24982(n23652,n22508,n23621);
  nand U24983(n23651,n23654,n23655,n23656);
  nand U24984(n23656,G59616,n22435);
  nand U24985(n23655,n21691,n23620);
  nand U24986(n23620,n23657,n23658);
  nand U24987(n23658,n23053,n21846);
  nand U24988(n23053,n23659,n23660,n23661,n23662);
  nor U24989(n23662,n23663,n23664,n23665,n23666);
  nor U24990(n23666,n23047,n23177);
  nor U24991(n23665,n23048,n23184);
  nor U24992(n23664,n23049,n23183);
  nor U24993(n23663,n23050,n23169);
  nor U24994(n23661,n23667,n23668,n23669,n23670);
  nor U24995(n23670,n23039,n23185);
  nor U24996(n23669,n23040,n23175);
  nor U24997(n23668,n23041,n23162);
  nor U24998(n23667,n23042,n23176);
  nor U24999(n23660,n23671,n23672,n23673,n23674);
  nor U25000(n23674,n23031,n23178);
  nor U25001(n23673,n23032,n23167);
  nor U25002(n23672,n23033,n23161);
  nor U25003(n23671,n23034,n23168);
  nor U25004(n23659,n23675,n23676,n23677,n23678);
  nor U25005(n23678,n23023,n23170);
  nor U25006(n23677,n23024,n23159);
  nor U25007(n23676,n23025,n23160);
  nor U25008(n23675,n23026,n23186);
  xnor U25009(n23657,n23576,n23575);
  nor U25010(n23575,n23679,n23680);
  nor U25011(n23576,n23621,n21846);
  not U25012(n23621,G59584);
  nand U25013(n23654,G59743,n22434);
  and U25014(n23644,n23681,n23682,n23683);
  nand U25015(n23683,G59616,n23278);
  nand U25016(n23682,G59584,n22496);
  nand U25017(n23681,G59775,n21108);
  nand U25018(n23610,n23684,n23685);
  nand U25019(n23685,n23686,n23687);
  not U25020(n23686,n23688);
  nand U25021(G8526,n23689,n23690,n23691,n23692);
  nor U25022(n23692,n23693,n23694,n23695);
  nor U25023(n23695,n23696,n22401);
  not U25024(n23696,G59774);
  and U25025(n23694,n23697,n22400);
  nor U25026(n23693,n23680,n22456);
  nand U25027(n23691,n22402,n21626);
  nand U25028(n23690,n22403,n21358);
  xor U25029(n21358,n23698,n23637);
  nand U25030(n23637,n23699,n23700);
  nand U25031(n23700,n22406,n23701);
  or U25032(n23701,n23702,n23703);
  nand U25033(n23699,n23703,n23702);
  xnor U25034(n23698,n23636,n22414);
  nand U25035(n23636,n23704,n23705,n23706,n23707);
  nor U25036(n23707,n23708,n23709);
  nor U25037(n23709,n22470,n23680);
  nor U25038(n23708,n21357,n22414);
  nand U25039(n23706,n22439,G59774);
  nand U25040(n23705,n21359,n23631);
  nand U25041(n23631,n22750,n23710);
  nand U25042(n23710,n23630,n22473);
  not U25043(n23630,n23462);
  nand U25044(n23704,n22473,n23462,n23629);
  not U25045(n23629,n21359);
  nand U25046(n23462,n23711,n23712);
  nand U25047(n23712,n23713,n23714);
  or U25048(n23713,n23715,n21369);
  nand U25049(n23711,n21369,n23715);
  nand U25050(n23689,n22440,n21359);
  xor U25051(n21359,n23716,n23688);
  nand U25052(n23716,n23684,n23687);
  nand U25053(n23687,n23717,n23718,n23719);
  nand U25054(n23684,n23721,n23720,n22567);
  nand U25055(n23721,n23717,n23718);
  nand U25056(n23718,n22435,n21357,n23722);
  nand U25057(n23717,n23723,n22383);
  nand U25058(n23723,n23722,n23724);
  nand U25059(n23724,n21626,n22497);
  not U25060(n21626,n21357);
  nand U25061(n21357,n23649,n23725);
  nand U25062(n23725,n23726,n23727);
  or U25063(n23649,n23727,n23726);
  and U25064(n23726,n23728,n23729);
  nand U25065(n23729,n23730,n23731);
  xor U25066(n23727,n21108,n23732);
  nor U25067(n23732,n23733,n23734,n23735);
  and U25068(n23735,n22437,G59710);
  nor U25069(n23734,n22508,n23680);
  nand U25070(n23733,n23736,n23737,n23738);
  nand U25071(n23738,G59615,n22435);
  nand U25072(n23737,n21691,n23697);
  nand U25073(n23697,n23739,n23740,n23741);
  nand U25074(n23741,n23742,n23680);
  not U25075(n23680,G59583);
  nand U25076(n23740,G59583,n23679,n21058);
  not U25077(n23679,n23742);
  nor U25078(n23742,n23743,n23744,n23745);
  nand U25079(n23739,n23187,n21846);
  nand U25080(n23187,n23746,n23747,n23748,n23749);
  nor U25081(n23749,n23750,n23751,n23752,n23753);
  nor U25082(n23753,n23140,n23177);
  nor U25083(n23752,n23144,n23184);
  nor U25084(n23751,n23145,n23183);
  nor U25085(n23750,n23147,n23169);
  nor U25086(n23748,n23754,n23755,n23756,n23757);
  nor U25087(n23757,n23131,n23185);
  nor U25088(n23756,n23133,n23175);
  nor U25089(n23755,n23134,n23162);
  nor U25090(n23754,n23135,n23176);
  nor U25091(n23747,n23758,n23759,n23760,n23761);
  nor U25092(n23761,n23121,n23178);
  nor U25093(n23760,n23123,n23167);
  nor U25094(n23759,n23124,n23161);
  nor U25095(n23758,n23125,n23168);
  nor U25096(n23746,n23762,n23763,n23764,n23765);
  nor U25097(n23765,n23106,n23170);
  nor U25098(n23764,n23109,n23159);
  nor U25099(n23763,n23111,n23160);
  nor U25100(n23762,n23113,n23186);
  nand U25101(n23736,G59742,n22434);
  and U25102(n23722,n23766,n23767,n23768);
  nand U25103(n23768,G59615,n23278);
  nand U25104(n23767,G59583,n22496);
  nand U25105(n23766,G59774,n21108);
  nand U25106(G8525,n23769,n23770,n23771,n23772);
  nor U25107(n23772,n23773,n23774,n23775);
  nor U25108(n23775,G59582,n22394,n23776,n23745);
  nor U25109(n23774,n23777,n23744);
  nor U25110(n23777,n23778,n22399);
  nor U25111(n23778,n23779,n22394);
  nor U25112(n23779,n23776,n23745);
  nor U25113(n23773,n23780,n22401);
  nand U25114(n23771,n22402,n21630);
  nand U25115(n23770,n22403,n21368);
  xor U25116(n21368,n23781,n23703);
  nand U25117(n23703,n23782,n23783,n23784,n23785);
  nor U25118(n23785,n23786,n23787);
  nor U25119(n23787,n23780,n22469);
  not U25120(n23780,G59773);
  nor U25121(n23786,n22470,n23744);
  not U25122(n23744,G59582);
  nand U25123(n23784,n22406,n21630);
  nand U25124(n23783,n22473,n23788);
  xor U25125(n23788,n23715,n23789);
  xor U25126(n23789,n21369,n23714);
  nand U25127(n23715,n23790,n23791);
  nand U25128(n23791,n23792,n23793);
  nand U25129(n23792,n23794,n23795);
  or U25130(n23790,n23794,n23795);
  nand U25131(n23782,n21369,n22423);
  xnor U25132(n23781,n22414,n23702);
  nand U25133(n23702,n23796,n23797);
  nand U25134(n23797,n22406,n23798);
  or U25135(n23798,n23799,n23800);
  nand U25136(n23796,n23800,n23799);
  nand U25137(n23769,n22440,n21369);
  and U25138(n21369,n23688,n23801);
  nand U25139(n23801,n23802,n23803);
  xnor U25140(n23802,n22435,n23804);
  nand U25141(n23688,n23805,n23806);
  xnor U25142(n23805,n23804,n22383);
  nand U25143(n23804,n23807,n23808,n23809,n23810);
  nand U25144(n23810,n21630,n22497);
  not U25145(n21630,n21367);
  xor U25146(n21367,n23811,n23730);
  nand U25147(n23730,n23812,n23813);
  nand U25148(n23813,n23814,n23815);
  nand U25149(n23811,n23731,n23728);
  nand U25150(n23728,n23816,n23714,n21691);
  nand U25151(n23731,n23817,n23818,n23819);
  nand U25152(n23819,n21691,n23714);
  nand U25153(n23714,n23820,n23821,n23822,n23823);
  nor U25154(n23823,n23824,n23825,n23826,n23827);
  nor U25155(n23827,n22563,n23828);
  nor U25156(n23826,n22561,n23829);
  nor U25157(n23825,n22559,n23830);
  nor U25158(n23824,n22551,n23831);
  nor U25159(n23822,n23832,n23833,n23834,n23835);
  nor U25160(n23835,n22549,n23836);
  nor U25161(n23834,n22547,n23837);
  nor U25162(n23833,n22539,n23838);
  nor U25163(n23832,n22537,n23839);
  nor U25164(n23821,n23840,n23841,n23842,n23843);
  nor U25165(n23843,n22535,n23844);
  nor U25166(n23842,n22527,n23845);
  nor U25167(n23841,n22525,n23846);
  nor U25168(n23840,n22523,n23847);
  nor U25169(n23820,n23848,n23849,n23850,n23851);
  nor U25170(n23851,n22565,n23852);
  nor U25171(n23850,n22553,n23853);
  nor U25172(n23849,n22541,n23854);
  nor U25173(n23848,n22529,n23855);
  nand U25174(n23818,n23856,n21108);
  nand U25175(n23817,n23816,n22167);
  nand U25176(n23816,n23857,n23858,n23856);
  and U25177(n23856,n23859,n23860);
  nand U25178(n23860,G59741,n22434);
  nand U25179(n23859,G59614,n22435);
  nand U25180(n23858,G59582,n22436);
  nand U25181(n23857,G59709,n22437);
  nand U25182(n23809,G59582,n22496);
  nand U25183(n23808,G59773,n21108);
  nand U25184(n23807,G59614,n23278);
  nand U25185(G8524,n23861,n23862,n23863,n23864);
  nor U25186(n23864,n23865,n23866,n23867);
  nor U25187(n23867,n21377,n22975);
  nor U25188(n23866,n23794,n23868);
  nor U25189(n23865,n23869,n22401);
  nand U25190(n23863,n22403,n21378);
  xor U25191(n21378,n23870,n23800);
  nand U25192(n23800,n23871,n23872,n23873,n23874);
  nor U25193(n23874,n23875,n23876);
  nor U25194(n23876,n23869,n22469);
  not U25195(n23869,G59772);
  nor U25196(n23875,n22470,n23776);
  not U25197(n23776,G59581);
  nand U25198(n23873,n22406,n21634);
  nand U25199(n23872,n23877,n22473);
  xor U25200(n23877,n23795,n23878);
  xnor U25201(n23878,n23793,n21379);
  nand U25202(n23795,n23879,n23880);
  nand U25203(n23880,n23881,n23882);
  or U25204(n23882,n23883,n23884);
  nand U25205(n23879,n23884,n23883);
  nand U25206(n23871,n21379,n22423);
  not U25207(n21379,n23794);
  nand U25208(n23794,n23803,n23885);
  nand U25209(n23885,n23886,n23887);
  not U25210(n23803,n23806);
  nor U25211(n23806,n23887,n23886);
  xor U25212(n23886,n23888,n22383);
  nand U25213(n23888,n23889,n23890,n23891,n23892);
  nand U25214(n23892,n21634,n22497);
  not U25215(n21634,n21377);
  xor U25216(n21377,n23893,n23815);
  nand U25217(n23815,n23894,n23895);
  nand U25218(n23895,n23896,n23897);
  nand U25219(n23893,n23812,n23814);
  nand U25220(n23814,n23898,n23899);
  nand U25221(n23899,n21691,n23793);
  xnor U25222(n23898,n21108,n23900);
  nand U25223(n23812,n23900,n23793,n21691);
  nand U25224(n23793,n23901,n23902,n23903,n23904);
  nor U25225(n23904,n23905,n23906,n23907,n23908);
  nor U25226(n23908,n23257,n23828);
  nor U25227(n23907,n23256,n23829);
  nor U25228(n23906,n23255,n23830);
  nor U25229(n23905,n23265,n23831);
  nor U25230(n23903,n23909,n23910,n23911,n23912);
  nor U25231(n23912,n23264,n23836);
  nor U25232(n23911,n23263,n23837);
  nor U25233(n23910,n22653,n23838);
  nor U25234(n23909,n22652,n23839);
  nor U25235(n23902,n23913,n23914,n23915,n23916);
  nor U25236(n23916,n22651,n23844);
  nor U25237(n23915,n22645,n23845);
  nor U25238(n23914,n22644,n23846);
  nor U25239(n23913,n22643,n23847);
  nor U25240(n23901,n23917,n23918,n23919,n23920);
  nor U25241(n23920,n23258,n23852);
  nor U25242(n23919,n23266,n23853);
  nor U25243(n23918,n22654,n23854);
  nor U25244(n23917,n22646,n23855);
  nand U25245(n23900,n23921,n23922,n23923,n23924);
  nand U25246(n23924,G59740,n22434);
  nand U25247(n23923,G59613,n22435);
  nand U25248(n23922,G59581,n22436);
  nand U25249(n23921,G59708,n22437);
  nand U25250(n23891,G59581,n22496);
  nand U25251(n23890,G59772,n21108);
  nand U25252(n23889,G59613,n23278);
  xnor U25253(n23870,n22414,n23799);
  nand U25254(n23799,n23925,n23926);
  nand U25255(n23926,n22406,n23927);
  nand U25256(n23927,n23928,n23929);
  or U25257(n23925,n23929,n23928);
  nand U25258(n23862,n23930,n23743,n22400);
  nand U25259(n23743,G59581,n21058);
  nand U25260(n23861,G59581,n23931);
  nand U25261(n23931,n22456,n23932);
  nand U25262(n23932,n22400,n23745);
  not U25263(n23745,n23930);
  nor U25264(n23930,n23933,n23934,n23935);
  nand U25265(G8523,n23936,n23937,n23938,n23939);
  nor U25266(n23939,n23940,n23941,n23942);
  nor U25267(n23942,G59580,n22394,n23943,n23935);
  nor U25268(n23941,n23944,n23934);
  nor U25269(n23944,n23945,n22399);
  nor U25270(n23945,n23946,n22394);
  nor U25271(n23946,n23943,n23935);
  nor U25272(n23940,n23947,n22401);
  nand U25273(n23938,n22402,n21638);
  nand U25274(n23937,n22403,n21388);
  xnor U25275(n21388,n23928,n23948);
  xnor U25276(n23948,n22406,n23929);
  nand U25277(n23929,n23949,n23950);
  nand U25278(n23950,n23951,n22414);
  nand U25279(n23951,n23952,n23953);
  or U25280(n23949,n23952,n23953);
  and U25281(n23928,n23954,n23955,n23956,n23957);
  nor U25282(n23957,n23958,n23959);
  nor U25283(n23959,n23947,n22469);
  not U25284(n23947,G59771);
  nor U25285(n23958,n22470,n23934);
  not U25286(n23934,G59580);
  nand U25287(n23956,n22406,n21638);
  nand U25288(n23955,n23960,n22473);
  xor U25289(n23960,n23884,n23961);
  xnor U25290(n23961,n23881,n23883);
  not U25291(n23881,n23962);
  nand U25292(n23884,n23963,n23964);
  nand U25293(n23964,n23965,n23966);
  or U25294(n23966,n23967,n23968);
  not U25295(n23965,n23969);
  nand U25296(n23963,n23968,n23967);
  nand U25297(n23954,n21389,n22423);
  nand U25298(n23936,n22440,n21389);
  not U25299(n21389,n23883);
  nand U25300(n23883,n23887,n23970);
  nand U25301(n23970,n23971,n23972);
  or U25302(n23887,n23972,n23971);
  xor U25303(n23971,n23973,n22383);
  nand U25304(n23973,n23974,n23975,n23976,n23977);
  nand U25305(n23977,n21638,n22497);
  not U25306(n21638,n21387);
  xor U25307(n21387,n23978,n23896);
  or U25308(n23896,n23979,n23980);
  nor U25309(n23980,n23981,n23982);
  nand U25310(n23978,n23897,n23894);
  nand U25311(n23894,n23983,n23962,n21691);
  nand U25312(n23897,n23984,n23985,n23986);
  nand U25313(n23986,n21691,n23962);
  nand U25314(n23962,n23987,n23988,n23989,n23990);
  nor U25315(n23990,n23991,n23992,n23993,n23994);
  nor U25316(n23994,n23337,n23828);
  nor U25317(n23993,n23336,n23829);
  nor U25318(n23992,n23335,n23830);
  nor U25319(n23991,n23345,n23831);
  nor U25320(n23989,n23995,n23996,n23997,n23998);
  nor U25321(n23998,n23344,n23836);
  nor U25322(n23997,n23343,n23837);
  nor U25323(n23996,n22729,n23838);
  nor U25324(n23995,n22728,n23839);
  nor U25325(n23988,n23999,n24000,n24001,n24002);
  nor U25326(n24002,n22727,n23844);
  nor U25327(n24001,n22721,n23845);
  nor U25328(n24000,n22720,n23846);
  nor U25329(n23999,n22719,n23847);
  nor U25330(n23987,n24003,n24004,n24005,n24006);
  nor U25331(n24006,n23338,n23852);
  nor U25332(n24005,n23346,n23853);
  nor U25333(n24004,n22730,n23854);
  nor U25334(n24003,n22722,n23855);
  nand U25335(n23985,n24007,n21108);
  nand U25336(n23984,n23983,n22167);
  nand U25337(n23983,n24008,n24009,n24007);
  and U25338(n24007,n24010,n24011);
  nand U25339(n24011,G59739,n22434);
  nand U25340(n24010,G59612,n22435);
  nand U25341(n24009,G59580,n22436);
  nand U25342(n24008,G59707,n22437);
  nand U25343(n23976,G59580,n22496);
  nand U25344(n23975,G59771,n21108);
  nand U25345(n23974,G59612,n23278);
  nand U25346(n23972,n24012,n24013);
  nand U25347(G8522,n24014,n24015,n24016,n24017);
  nor U25348(n24017,n24018,n24019,n24020);
  nor U25349(n24020,n21397,n22975);
  not U25350(n21397,n21642);
  nor U25351(n24019,n23968,n23868);
  nor U25352(n24018,n24021,n22401);
  nand U25353(n24016,n22403,n21398);
  xnor U25354(n21398,n23953,n24022);
  xnor U25355(n24022,n22406,n23952);
  nand U25356(n23952,n24023,n24024,n24025,n24026);
  nor U25357(n24026,n24027,n24028);
  nor U25358(n24028,n24021,n22469);
  not U25359(n24021,G59770);
  nor U25360(n24027,n22470,n23943);
  not U25361(n23943,G59579);
  nand U25362(n24025,n22406,n21642);
  nand U25363(n24024,n22473,n24029);
  xnor U25364(n24029,n23968,n24030);
  xnor U25365(n24030,n23967,n23969);
  nand U25366(n23967,n24031,n24032);
  nand U25367(n24032,n24033,n24034);
  or U25368(n24034,n24035,n24036);
  not U25369(n24033,n24037);
  nand U25370(n24031,n24036,n24035);
  nand U25371(n24023,n21399,n22423);
  not U25372(n21399,n23968);
  xnor U25373(n23968,n24013,n24012);
  xnor U25374(n24013,n24038,n22383);
  nand U25375(n24038,n24039,n24040,n24041,n24042);
  nand U25376(n24042,n21642,n22497);
  xnor U25377(n21642,n23981,n24043);
  nor U25378(n24043,n23979,n23982);
  and U25379(n23982,n24044,n24045,n24046);
  nand U25380(n24046,n24047,n21108);
  nor U25381(n23979,n24045,n24044);
  nand U25382(n24044,n21691,n23969);
  nand U25383(n23969,n24048,n24049,n24050,n24051);
  nor U25384(n24051,n24052,n24053,n24054,n24055);
  nor U25385(n24055,n22801,n23846);
  nor U25386(n24054,n22802,n23845);
  nor U25387(n24053,n22810,n23838);
  nor U25388(n24052,n23426,n23831);
  nor U25389(n24050,n24056,n24057,n24058,n24059);
  nor U25390(n24059,n22809,n23839);
  nor U25391(n24058,n22811,n23854);
  nor U25392(n24057,n23419,n23852);
  nor U25393(n24056,n22800,n23847);
  nor U25394(n24049,n24060,n24061,n24062,n24063);
  nor U25395(n24063,n23425,n23836);
  nor U25396(n24062,n23427,n23853);
  nor U25397(n24061,n23416,n23830);
  nor U25398(n24060,n22808,n23844);
  nor U25399(n24048,n24064,n24065,n24066,n24067);
  nor U25400(n24067,n23417,n23829);
  nor U25401(n24066,n23424,n23837);
  nor U25402(n24065,n22803,n23855);
  nor U25403(n24064,n23418,n23828);
  nand U25404(n24045,n24068,n22167);
  nand U25405(n24068,n24069,n24070,n24047);
  and U25406(n24047,n24071,n24072);
  nand U25407(n24072,G59738,n22434);
  nand U25408(n24071,G59611,n22435);
  nand U25409(n24070,G59579,n22436);
  nand U25410(n24069,G59706,n22437);
  nand U25411(n23981,n24073,n24074);
  nand U25412(n24074,n24075,n24076,n24077);
  nand U25413(n24041,G59579,n22496);
  nand U25414(n24040,G59770,n21108);
  nand U25415(n24039,G59611,n23278);
  nand U25416(n23953,n24078,n24079,n24080);
  or U25417(n24080,n22414,n24081);
  nor U25418(n24081,n24082,n24083,n24084);
  nand U25419(n24078,n24084,n24085,n24083);
  nand U25420(n24015,n24086,n23933,n22400);
  nand U25421(n23933,G59579,n21058);
  nand U25422(n24014,G59579,n24087);
  nand U25423(n24087,n22456,n24088);
  nand U25424(n24088,n22400,n23935);
  not U25425(n23935,n24086);
  nor U25426(n24086,n24089,n24090,n24091,n24092);
  nand U25427(G8521,n24093,n24094,n24095,n24096);
  nor U25428(n24096,n24097,n24098,n24099);
  nor U25429(n24099,G59578,n24092,n24100);
  nor U25430(n24098,n24101,n24090);
  nor U25431(n24101,n24102,n24103);
  nor U25432(n24102,G59577,n22394);
  nor U25433(n24097,n24104,n22401);
  nand U25434(n24095,n22402,n21646);
  nand U25435(n24094,n22403,n21408);
  xnor U25436(n21408,n24105,n24106);
  nor U25437(n24106,n24082,n24107);
  not U25438(n24082,n24108);
  xnor U25439(n24105,n24084,n22414);
  nand U25440(n24084,n24109,n24110,n24111,n24112);
  nor U25441(n24112,n24113,n24114);
  nor U25442(n24114,n24104,n22469);
  not U25443(n24104,G59769);
  nor U25444(n24113,n22470,n24090);
  not U25445(n24090,G59578);
  nand U25446(n24111,n22406,n21646);
  nand U25447(n24110,n24115,n22473);
  xnor U25448(n24115,n24116,n24036);
  not U25449(n24036,n21409);
  xnor U25450(n24116,n24035,n24037);
  nand U25451(n24035,n24117,n24118);
  nand U25452(n24118,n24119,n24120);
  nand U25453(n24120,n21422,n24121);
  nand U25454(n24117,n24122,n22312);
  nand U25455(n24109,n21409,n22423);
  nand U25456(n24093,n22440,n21409);
  nor U25457(n21409,n24012,n24123);
  and U25458(n24123,n24124,n24125);
  nor U25459(n24012,n24125,n24124);
  xor U25460(n24124,n24126,n22383);
  nand U25461(n24126,n24127,n24128,n24129,n24130);
  nand U25462(n24130,n21646,n22497);
  not U25463(n21646,n21407);
  xnor U25464(n21407,n24131,n24132);
  and U25465(n24132,n24077,n24073);
  nand U25466(n24073,n24133,n24134,n24135);
  nand U25467(n24135,n21691,n24037);
  nand U25468(n24134,n24136,n22167);
  nand U25469(n24133,n24137,n21108);
  nand U25470(n24077,n24136,n24037,n21691);
  nand U25471(n24037,n24138,n24139,n24140,n24141);
  nor U25472(n24141,n24142,n24143,n24144,n24145);
  nor U25473(n24145,n22875,n23846);
  nor U25474(n24144,n22876,n23845);
  nor U25475(n24143,n22884,n23838);
  nor U25476(n24142,n23510,n23831);
  nor U25477(n24140,n24146,n24147,n24148,n24149);
  nor U25478(n24149,n22883,n23839);
  nor U25479(n24148,n22885,n23854);
  nor U25480(n24147,n23503,n23852);
  nor U25481(n24146,n22874,n23847);
  nor U25482(n24139,n24150,n24151,n24152,n24153);
  nor U25483(n24153,n23509,n23836);
  nor U25484(n24152,n23511,n23853);
  nor U25485(n24151,n23500,n23830);
  nor U25486(n24150,n22882,n23844);
  nor U25487(n24138,n24154,n24155,n24156,n24157);
  nor U25488(n24157,n23501,n23829);
  nor U25489(n24156,n23508,n23837);
  nor U25490(n24155,n22877,n23855);
  nor U25491(n24154,n23502,n23828);
  nand U25492(n24136,n24158,n24159,n24137);
  and U25493(n24137,n24160,n24161);
  nand U25494(n24161,G59737,n22434);
  nand U25495(n24160,G59610,n22435);
  nand U25496(n24159,G59578,n22436);
  nand U25497(n24158,G59705,n22437);
  nand U25498(n24131,n24076,n24075);
  nand U25499(n24129,G59578,n22496);
  nand U25500(n24128,G59769,n21108);
  nand U25501(n24127,G59610,n23278);
  nand U25502(G8520,n24162,n24163,n24164,n24165);
  nor U25503(n24165,n24166,n24167,n24168);
  nor U25504(n24168,G59577,n24100);
  nand U25505(n24100,n24169,G59576,n22400);
  and U25506(n24167,n24103,G59577);
  nand U25507(n24103,n24170,n24171);
  nand U25508(n24171,n22400,n24091);
  nor U25509(n24166,n22314,n22401);
  nand U25510(n24164,n22402,n21650);
  nand U25511(n24163,n22403,n21881);
  not U25512(n21881,n21421);
  nand U25513(n21421,n24172,n24173);
  nand U25514(n24173,n24174,n24079,n24175);
  nand U25515(n24175,n24176,n24108);
  nand U25516(n24172,n24108,n24107);
  nand U25517(n24107,n24079,n24177);
  nand U25518(n24177,n24083,n24176);
  or U25519(n24176,n24085,n22406);
  not U25520(n24083,n24174);
  nand U25521(n24174,n24178,n24179);
  nand U25522(n24179,n24180,n22414);
  nand U25523(n24108,n22406,n24085);
  nand U25524(n24085,n24181,n24182,n24183,n24184);
  nor U25525(n24184,n24185,n24186);
  nor U25526(n24186,n22314,n22469);
  not U25527(n22314,G59768);
  nor U25528(n24185,n22470,n24092);
  nand U25529(n24183,n22406,n21650);
  nand U25530(n24182,n22473,n24187);
  xnor U25531(n24187,n21422,n24188);
  xnor U25532(n24188,n24119,n24122);
  and U25533(n24119,n24189,n24190);
  nand U25534(n24190,n24191,n24192,n21442);
  nand U25535(n24181,n21422,n22423);
  nand U25536(n24162,n22440,n21422);
  not U25537(n21422,n22312);
  nand U25538(n22312,n24193,n24125);
  nand U25539(n24125,n24194,n24195,n24196);
  xnor U25540(n24196,n24197,n22383);
  nand U25541(n24193,n24198,n24199);
  nand U25542(n24199,n24195,n24194);
  xnor U25543(n24198,n22435,n24197);
  nand U25544(n24197,n24200,n24201,n24202,n24203);
  nand U25545(n24203,n21650,n22497);
  not U25546(n21650,n21417);
  nand U25547(n21417,n24204,n24205);
  or U25548(n24205,n24075,n24206);
  nand U25549(n24075,n24207,n24208);
  nand U25550(n24208,n24209,n24210);
  nand U25551(n24204,n24211,n24210,n24209);
  nand U25552(n24209,n24212,n24213);
  nand U25553(n24211,n24207,n24076);
  not U25554(n24076,n24206);
  nor U25555(n24206,n21114,n24122,n24214);
  not U25556(n24122,n24121);
  nand U25557(n24207,n24214,n24215);
  nand U25558(n24215,n21691,n24121);
  nand U25559(n24121,n24216,n24217,n24218,n24219);
  nor U25560(n24219,n24220,n24221,n24222,n24223);
  nor U25561(n24223,n23587,n23828);
  nor U25562(n24222,n23586,n23829);
  nor U25563(n24221,n23585,n23830);
  nor U25564(n24220,n23595,n23831);
  nor U25565(n24218,n24224,n24225,n24226,n24227);
  nor U25566(n24227,n23594,n23836);
  nor U25567(n24226,n23593,n23837);
  nor U25568(n24225,n22963,n23838);
  nor U25569(n24224,n22962,n23839);
  nor U25570(n24217,n24228,n24229,n24230,n24231);
  nor U25571(n24231,n22961,n23844);
  nor U25572(n24230,n22955,n23845);
  nor U25573(n24229,n22954,n23846);
  nor U25574(n24228,n22953,n23847);
  nor U25575(n24216,n24232,n24233,n24234,n24235);
  nor U25576(n24235,n23588,n23852);
  nor U25577(n24234,n23596,n23853);
  nor U25578(n24233,n22964,n23854);
  nor U25579(n24232,n22956,n23855);
  xor U25580(n24214,n21108,n24236);
  nor U25581(n24236,n24237,n24238,n24239,n24240);
  and U25582(n24240,n22437,G59704);
  nor U25583(n24239,n22508,n24092);
  not U25584(n24092,G59577);
  and U25585(n24238,n22435,G59609);
  nor U25586(n24237,n24241,n21418);
  not U25587(n21418,G59736);
  nand U25588(n24202,G59577,n22496);
  nand U25589(n24201,G59768,n21108);
  nand U25590(n24200,G59609,n23278);
  nand U25591(G8519,n24242,n24243,n24244,n24245);
  nor U25592(n24245,n24246,n24247,n24248);
  nor U25593(n24248,G59576,n24089,n22394);
  nor U25594(n24247,n24170,n24091);
  and U25595(n24170,n22456,n24249);
  nand U25596(n24249,n22400,n24089);
  not U25597(n24089,n24169);
  nor U25598(n24169,n24250,n24251,n24252);
  nor U25599(n24246,n24253,n22401);
  nand U25600(n24244,n22402,n21654);
  nand U25601(n24243,n22403,n21431);
  nand U25602(n21431,n24254,n24255,n24256);
  or U25603(n24256,n24079,n24257);
  nand U25604(n24079,n22406,n24258);
  nand U25605(n24255,n24257,n24180,n22406);
  not U25606(n24180,n24258);
  nand U25607(n24254,n24259,n22414);
  xnor U25608(n24259,n24258,n24257);
  not U25609(n24257,n24178);
  nand U25610(n24178,n24260,n24261);
  nand U25611(n24261,n22406,n24262);
  or U25612(n24262,n24263,n24264);
  nand U25613(n24260,n24264,n24263);
  nand U25614(n24258,n24265,n24266,n24267,n24268);
  nor U25615(n24268,n24269,n24270);
  nor U25616(n24270,n24253,n22469);
  not U25617(n24253,G59767);
  nor U25618(n24269,n22470,n24091);
  not U25619(n24091,G59576);
  nand U25620(n24267,n22406,n21654);
  nand U25621(n24266,n22473,n24271);
  xor U25622(n24271,n24272,n24273);
  nand U25623(n24273,n21442,n24192);
  nand U25624(n24272,n24191,n24189);
  nand U25625(n24189,n21432,n24274);
  or U25626(n24191,n24274,n21432);
  nand U25627(n24265,n21432,n22423);
  nand U25628(n24242,n22440,n21432);
  xor U25629(n21432,n24195,n24194);
  xor U25630(n24194,n24275,n22435);
  nand U25631(n24275,n24276,n24277,n24278,n24279);
  nand U25632(n24279,n21654,n22497);
  not U25633(n21654,n21430);
  xnor U25634(n21430,n24213,n24280);
  and U25635(n24280,n24212,n24210);
  nand U25636(n24210,n24281,n24274,n21691);
  nand U25637(n24212,n24282,n24283,n24284);
  nand U25638(n24284,n21691,n24274);
  nand U25639(n24274,n24285,n24286,n24287,n24288);
  nor U25640(n24288,n24289,n24290,n24291,n24292);
  nor U25641(n24292,n23049,n23828);
  nor U25642(n24291,n23048,n23829);
  nor U25643(n24290,n23047,n23830);
  nor U25644(n24289,n23041,n23831);
  nor U25645(n24287,n24293,n24294,n24295,n24296);
  nor U25646(n24296,n23040,n23836);
  nor U25647(n24295,n23039,n23837);
  nor U25648(n24294,n23033,n23838);
  nor U25649(n24293,n23032,n23839);
  nor U25650(n24286,n24297,n24298,n24299,n24300);
  nor U25651(n24300,n23031,n23844);
  nor U25652(n24299,n23025,n23845);
  nor U25653(n24298,n23024,n23846);
  nor U25654(n24297,n23023,n23847);
  nor U25655(n24285,n24301,n24302,n24303,n24304);
  nor U25656(n24304,n23050,n23852);
  nor U25657(n24303,n23042,n23853);
  nor U25658(n24302,n23034,n23854);
  nor U25659(n24301,n23026,n23855);
  nand U25660(n24283,n24281,n22167);
  nand U25661(n24281,n24305,n24306,n24307);
  nand U25662(n24306,G59576,n22436);
  nand U25663(n24305,G59703,n22437);
  nand U25664(n24282,n24307,n21108);
  and U25665(n24307,n24308,n24309);
  nand U25666(n24309,G59735,n22434);
  nand U25667(n24308,G59608,n22435);
  nand U25668(n24213,n24310,n24311);
  nand U25669(n24311,n24312,n24313);
  not U25670(n24312,n24314);
  nand U25671(n24278,G59576,n22496);
  nand U25672(n24277,G59767,n21108);
  nand U25673(n24276,G59608,n23278);
  nand U25674(G8518,n24315,n24316,n24317,n24318);
  nor U25675(n24318,n24319,n24320,n24321);
  nor U25676(n24321,G59575,n22394,n24251,n24252);
  not U25677(n24251,G59574);
  nor U25678(n24320,n24322,n24250);
  nor U25679(n24322,n24323,n24324);
  nor U25680(n24323,G59574,n22394);
  nor U25681(n24319,n24325,n22401);
  nand U25682(n24317,n22402,n21658);
  nand U25683(n24316,n22403,n21441);
  xnor U25684(n21441,n24326,n24263);
  nand U25685(n24263,n24327,n24328,n24329,n24330);
  nor U25686(n24330,n24331,n24332);
  nor U25687(n24332,n24325,n22469);
  not U25688(n24325,G59766);
  nor U25689(n24331,n22470,n24250);
  not U25690(n24250,G59575);
  nand U25691(n24329,n22406,n21658);
  nand U25692(n24328,n24333,n22473);
  xor U25693(n24333,n21442,n24192);
  nand U25694(n24327,n21442,n22423);
  xnor U25695(n24326,n22406,n24264);
  nor U25696(n24264,n24334,n24335);
  nor U25697(n24334,n24336,n24337);
  nand U25698(n24315,n22440,n21442);
  nor U25699(n21442,n24195,n24338);
  and U25700(n24338,n24339,n24340);
  nor U25701(n24195,n24340,n24339);
  xor U25702(n24339,n24341,n22383);
  nand U25703(n24341,n24342,n24343,n24344,n24345);
  nand U25704(n24345,n21658,n22497);
  xor U25705(n21658,n24346,n24314);
  nand U25706(n24346,n24310,n24313);
  nand U25707(n24313,n24347,n24348,n24349);
  nand U25708(n24349,n21691,n24192);
  nand U25709(n24348,n24350,n21108);
  nand U25710(n24347,n24351,n22167);
  nand U25711(n24310,n24351,n24192,n21691);
  nand U25712(n24192,n24352,n24353,n24354,n24355);
  nor U25713(n24355,n24356,n24357,n24358,n24359);
  nor U25714(n24359,n23111,n23845);
  nand U25715(n23845,n24360,n24361);
  nor U25716(n24358,n23113,n23855);
  nand U25717(n23855,n24360,n24362);
  nor U25718(n24357,n23125,n23854);
  nand U25719(n23854,n24363,n24362);
  nor U25720(n24356,n23135,n23853);
  nand U25721(n23853,n24364,n24362);
  nor U25722(n24354,n24365,n24366,n24367,n24368);
  nor U25723(n24368,n23124,n23838);
  nand U25724(n23838,n24363,n24361);
  nor U25725(n24367,n23131,n23837);
  nand U25726(n23837,n24364,n24369);
  nor U25727(n24366,n23106,n23847);
  nand U25728(n23847,n24360,n24369);
  nor U25729(n24365,n23109,n23846);
  nand U25730(n23846,n24360,n24370);
  nor U25731(n24360,n24371,n24372);
  nor U25732(n24353,n24373,n24374,n24375,n24376);
  nor U25733(n24376,n23134,n23831);
  nand U25734(n23831,n24364,n24361);
  nor U25735(n24375,n23140,n23830);
  nand U25736(n23830,n24377,n24369);
  nor U25737(n24374,n23144,n23829);
  nand U25738(n23829,n24377,n24370);
  nor U25739(n24373,n23123,n23839);
  nand U25740(n23839,n24363,n24370);
  nor U25741(n24352,n24378,n24379,n24380,n24381);
  nor U25742(n24381,n23147,n23852);
  nand U25743(n23852,n24377,n24362);
  nor U25744(n24380,n23145,n23828);
  nand U25745(n23828,n24377,n24361);
  nor U25746(n24377,n24382,n24383);
  nor U25747(n24379,n23133,n23836);
  nand U25748(n23836,n24364,n24370);
  nor U25749(n24364,n24383,n24371);
  not U25750(n24371,n24382);
  nor U25751(n24378,n23121,n23844);
  nand U25752(n23844,n24363,n24369);
  nor U25753(n24363,n24382,n24372);
  not U25754(n24372,n24383);
  nand U25755(n24383,n24384,n24385,n24386);
  not U25756(n24386,n24387);
  nand U25757(n24385,G59558,n24388);
  nand U25758(n24384,n24389,G59560);
  xnor U25759(n24382,G59559,n24388);
  nand U25760(n24351,n24390,n24391,n24350);
  and U25761(n24350,n24392,n24393);
  nand U25762(n24393,G59734,n22434);
  nand U25763(n24392,G59607,n22435);
  nand U25764(n24391,G59575,n22436);
  nand U25765(n24390,G59702,n22437);
  nand U25766(n24344,G59575,n22496);
  nand U25767(n24343,G59766,n21108);
  nand U25768(n24342,G59607,n23278);
  or U25769(n24340,n24394,n24395);
  nand U25770(G8517,n24396,n24397,n24398,n24399);
  nor U25771(n24399,n24400,n24401,n24402);
  nor U25772(n24402,G59574,n24252,n22394);
  and U25773(n24401,n24324,G59574);
  nand U25774(n24324,n22456,n24403);
  nand U25775(n24403,n22400,n24252);
  or U25776(n24252,n24404,n24405);
  nor U25777(n24400,n24406,n22401);
  not U25778(n24406,G59765);
  nand U25779(n24398,n22402,n21662);
  nand U25780(n24397,n22403,n21451);
  xor U25781(n21451,n24336,n24407);
  nor U25782(n24407,n24337,n24335);
  nor U25783(n24335,n24408,n24409);
  and U25784(n24337,n24409,n24408);
  nand U25785(n24408,n24410,n24411,n24412,n24413);
  nand U25786(n24413,n24414,n21452);
  nand U25787(n24412,n21662,n22406);
  nand U25788(n24411,G59574,n22438);
  nand U25789(n24410,n22439,G59765);
  xnor U25790(n24409,n22414,n24415);
  nand U25791(n24415,n24416,n24417,n24418,n24419);
  nand U25792(n24419,n24420,n24421,n24422,n24423);
  nor U25793(n24423,n24424,n24425,n24426,n24427);
  nor U25794(n24427,n22541,n24428);
  nor U25795(n24426,n22553,n24429);
  nor U25796(n24425,n22529,n24430);
  nand U25797(n24424,n24431,n24432);
  nand U25798(n24432,n24433,G59445);
  nand U25799(n24431,n24434,G59437);
  nor U25800(n24422,n24435,n24436,n24437,n24438);
  nor U25801(n24438,n22539,n24439);
  nor U25802(n24437,n22547,n24440);
  nor U25803(n24436,n22565,n24441);
  nor U25804(n24435,n22523,n24442);
  nor U25805(n24421,n24443,n24444,n24445,n24446);
  nor U25806(n24446,n22551,n24447);
  nor U25807(n24445,n22549,n24448);
  nor U25808(n24444,n22535,n24449);
  nor U25809(n24443,n22537,n24450);
  nor U25810(n24420,n24451,n24452,n24453,n22414);
  nor U25811(n24453,n22561,n24454);
  nor U25812(n24452,n22563,n24455);
  nor U25813(n24451,n22559,n24456);
  nand U25814(n24418,n24457,n23079);
  nand U25815(n23079,n24458,n24459,n24460,n24461);
  nor U25816(n24461,n24462,n24463,n24464,n24465);
  nor U25817(n24465,n22563,n24466);
  nor U25818(n24464,n22561,n24467);
  nor U25819(n24463,n22559,n24468);
  nor U25820(n24462,n22551,n24469);
  nor U25821(n24460,n24470,n24471,n24472,n24473);
  nor U25822(n24473,n22549,n24474);
  nor U25823(n24472,n22547,n24475);
  nor U25824(n24471,n22539,n24476);
  nor U25825(n24470,n22537,n24477);
  nor U25826(n24459,n24478,n24479,n24480,n24481);
  nor U25827(n24481,n22535,n24482);
  nor U25828(n24480,n22527,n24483);
  nor U25829(n24479,n22525,n24484);
  nor U25830(n24478,n22523,n24485);
  nor U25831(n24458,n24486,n24487,n24488,n24489);
  nor U25832(n24489,n22565,n24490);
  nor U25833(n24488,n22553,n24491);
  nor U25834(n24487,n22541,n24492);
  nor U25835(n24486,n22529,n24493);
  nand U25836(n24417,n22473,n24494);
  nand U25837(n24494,n24495,n24496,n24497,n24498);
  nor U25838(n24498,n24499,n24500,n24501,n24502);
  nor U25839(n24502,n22565,n24503);
  nor U25840(n24501,n22563,n24504);
  nor U25841(n24500,n22561,n24505);
  nor U25842(n24499,n22559,n24506);
  nor U25843(n24497,n24507,n24508,n24509,n24510);
  nor U25844(n24510,n22553,n24511);
  nor U25845(n24509,n22551,n24512);
  nor U25846(n24508,n22549,n24513);
  nor U25847(n24507,n22547,n24514);
  nor U25848(n24496,n24515,n24516,n24517,n24518);
  nor U25849(n24518,n22541,n24519);
  nor U25850(n24517,n22539,n24520);
  nor U25851(n24516,n22537,n24521);
  nor U25852(n24515,n22535,n24522);
  nor U25853(n24495,n24523,n24524,n24525,n24526);
  nor U25854(n24526,n22529,n24527);
  nor U25855(n24525,n22527,n24528);
  nor U25856(n24524,n22525,n24529);
  nor U25857(n24523,n22523,n24530);
  nand U25858(n24416,n24531,n24532);
  nand U25859(n24336,n24533,n24534);
  nand U25860(n24396,n22440,n21452);
  nand U25861(n21452,n24535,n24536);
  nand U25862(n24536,n24537,n24538);
  or U25863(n24537,n24395,n24539);
  not U25864(n24395,n24540);
  nand U25865(n24535,n24394,n24540);
  nand U25866(n24540,n24541,n24542);
  nand U25867(n24542,n21691,G59549);
  nor U25868(n24394,n24538,n24539);
  nor U25869(n24539,n22565,n24541,n21114);
  nor U25870(n24541,n24543,n24544);
  and U25871(n24544,n24545,n22383);
  nor U25872(n24543,n24545,n21662,n22383);
  not U25873(n21662,n21450);
  nand U25874(n21450,n24314,n24546);
  nand U25875(n24546,n24547,n24548);
  xnor U25876(n24547,n22167,n24549);
  nand U25877(n24314,n24550,n24551);
  xnor U25878(n24550,n21108,n24549);
  and U25879(n24549,n24552,n24553,n24554,n24555);
  nand U25880(n24555,G59733,n22434);
  nand U25881(n24554,G59606,n22435);
  nand U25882(n24553,G59574,n22436);
  nand U25883(n24552,G59701,n22437);
  nand U25884(n24545,n24556,n24557,n24558);
  nand U25885(n24558,G59606,n23278);
  nand U25886(n24557,G59574,n22496);
  nand U25887(n24556,G59765,n21108);
  or U25888(n24538,n24559,n24560);
  and U25889(n24560,n24561,n24562);
  nand U25890(G8516,n24563,n24564,n24565,n24566);
  nor U25891(n24566,n24567,n24568,n24569);
  nor U25892(n24569,n21460,n22975);
  and U25893(n24568,n21463,n22440);
  nor U25894(n24567,n24570,n22401);
  not U25895(n24570,G59764);
  nand U25896(n24565,n22403,n21902);
  not U25897(n21902,n21462);
  nand U25898(n21462,n24571,n24572);
  nand U25899(n24572,n24573,n24574,n24575);
  nand U25900(n24573,n24576,n24533);
  nand U25901(n24571,n24577,n24533);
  nand U25902(n24533,n24578,n24579);
  xnor U25903(n24578,n24580,n22414);
  not U25904(n24577,n24534);
  nand U25905(n24534,n24576,n24581);
  nand U25906(n24581,n24575,n24574);
  nand U25907(n24575,n24582,n24583);
  nand U25908(n24576,n24584,n24585);
  xnor U25909(n24585,n22406,n24580);
  nand U25910(n24580,n24586,n24587,n24588,n24589);
  nand U25911(n24589,n24590,n24591,n24592,n24593);
  nor U25912(n24593,n24594,n24595,n24596,n24597);
  nor U25913(n24597,n22654,n24428);
  nor U25914(n24596,n23266,n24429);
  nor U25915(n24595,n22646,n24430);
  nand U25916(n24594,n24598,n24599);
  nand U25917(n24599,n24433,G59446);
  nand U25918(n24598,n24434,G59438);
  nor U25919(n24592,n24600,n24601,n24602,n24603);
  nor U25920(n24603,n22653,n24439);
  nor U25921(n24602,n23263,n24440);
  nor U25922(n24601,n23258,n24441);
  nor U25923(n24600,n22643,n24442);
  nor U25924(n24591,n24604,n24605,n24606,n24607);
  nor U25925(n24607,n23265,n24447);
  nor U25926(n24606,n23264,n24448);
  nor U25927(n24605,n22651,n24449);
  nor U25928(n24604,n22652,n24450);
  nor U25929(n24590,n24608,n24609,n24610,n22414);
  nor U25930(n24610,n23256,n24454);
  nor U25931(n24609,n23257,n24455);
  nor U25932(n24608,n23255,n24456);
  nand U25933(n24588,n24457,n23225);
  nand U25934(n23225,n24611,n24612,n24613,n24614);
  nor U25935(n24614,n24615,n24616,n24617,n24618);
  nor U25936(n24618,n23257,n24466);
  nor U25937(n24617,n23256,n24467);
  nor U25938(n24616,n23255,n24468);
  nor U25939(n24615,n23265,n24469);
  nor U25940(n24613,n24619,n24620,n24621,n24622);
  nor U25941(n24622,n23264,n24474);
  nor U25942(n24621,n23263,n24475);
  nor U25943(n24620,n22653,n24476);
  nor U25944(n24619,n22652,n24477);
  nor U25945(n24612,n24623,n24624,n24625,n24626);
  nor U25946(n24626,n22651,n24482);
  nor U25947(n24625,n22645,n24483);
  nor U25948(n24624,n22644,n24484);
  nor U25949(n24623,n22643,n24485);
  nor U25950(n24611,n24627,n24628,n24629,n24630);
  nor U25951(n24630,n23258,n24490);
  nor U25952(n24629,n23266,n24491);
  nor U25953(n24628,n22654,n24492);
  nor U25954(n24627,n22646,n24493);
  nand U25955(n24587,n24531,n24631);
  nand U25956(n24631,n24632,n24633,n24634,n24635);
  nor U25957(n24635,n24636,n24637,n24638,n24639);
  nor U25958(n24639,n23256,n24640);
  nor U25959(n24638,n23255,n24641);
  nor U25960(n24637,n23266,n24642);
  nor U25961(n24636,n23264,n24643);
  nor U25962(n24634,n24644,n24645,n24646,n24647);
  nor U25963(n24647,n23263,n24648);
  nor U25964(n24646,n22654,n24649);
  nor U25965(n24645,n22652,n24650);
  nor U25966(n24644,n22651,n24651);
  nor U25967(n24633,n24652,n24653,n24654,n24655);
  nor U25968(n24655,n22646,n24656);
  nor U25969(n24654,n22644,n24657);
  nor U25970(n24653,n22643,n24658);
  nor U25971(n24652,n23258,n24659);
  nor U25972(n24632,n24660,n24661,n24662,n24663);
  nor U25973(n24663,n23257,n24664);
  nor U25974(n24662,n23265,n24665);
  nor U25975(n24661,n22653,n24666);
  nor U25976(n24660,n22645,n24667);
  nand U25977(n24586,n22473,n24668);
  nand U25978(n24668,n24669,n24670,n24671,n24672);
  nor U25979(n24672,n24673,n24674,n24675,n24676);
  nor U25980(n24676,n23258,n24503);
  nor U25981(n24675,n23257,n24504);
  nor U25982(n24674,n23256,n24505);
  nor U25983(n24673,n23255,n24506);
  nor U25984(n24671,n24677,n24678,n24679,n24680);
  nor U25985(n24680,n23266,n24511);
  nor U25986(n24679,n23265,n24512);
  nor U25987(n24678,n23264,n24513);
  nor U25988(n24677,n23263,n24514);
  nor U25989(n24670,n24681,n24682,n24683,n24684);
  nor U25990(n24684,n22654,n24519);
  nor U25991(n24683,n22653,n24520);
  nor U25992(n24682,n22652,n24521);
  nor U25993(n24681,n22651,n24522);
  nor U25994(n24669,n24685,n24686,n24687,n24688);
  nor U25995(n24688,n22646,n24527);
  nor U25996(n24687,n22645,n24528);
  nor U25997(n24686,n22644,n24529);
  nor U25998(n24685,n22643,n24530);
  not U25999(n24584,n24579);
  nand U26000(n24579,n24689,n24690,n24691,n24692);
  nand U26001(n24692,n21463,n24414);
  xor U26002(n21463,n24562,n24693);
  nor U26003(n24693,n24559,n24694);
  not U26004(n24694,n24561);
  nand U26005(n24561,n24695,n24696);
  nand U26006(n24696,n21691,G59550);
  nor U26007(n24559,n21114,n23258,n24695);
  xor U26008(n24695,n24697,n22383);
  nand U26009(n24697,n24698,n24699,n24700,n24701);
  nand U26010(n24701,n21666,n22497);
  nand U26011(n24700,G59573,n22496);
  nand U26012(n24699,G59764,n21108);
  nand U26013(n24698,G59605,n23278);
  nand U26014(n24562,n24702,n24703);
  nand U26015(n24703,n24704,n24705);
  nand U26016(n24704,n24706,n24707);
  nand U26017(n24707,n21691,G59551);
  not U26018(n24702,n24708);
  nand U26019(n24691,n22406,n21666);
  not U26020(n21666,n21460);
  nand U26021(n21460,n24548,n24709);
  nand U26022(n24709,n24710,n24711);
  not U26023(n24548,n24551);
  nor U26024(n24551,n24711,n24710);
  xor U26025(n24710,n21108,n24712);
  nor U26026(n24712,n24713,n24714,n24715,n24716);
  and U26027(n24716,n22437,G59700);
  and U26028(n24715,n22436,G59573);
  nor U26029(n24714,n22383,n22340);
  not U26030(n22340,G59605);
  nor U26031(n24713,n24241,n21461);
  not U26032(n21461,G59732);
  nand U26033(n24690,G59573,n22438);
  nand U26034(n24689,n22439,G59764);
  nand U26035(n24564,n24717,n24405,n22400);
  nand U26036(n24405,G59573,n21058);
  nand U26037(n24563,G59573,n24718);
  nand U26038(n24718,n22456,n24719);
  nand U26039(n24719,n22400,n24404);
  not U26040(n24404,n24717);
  nor U26041(n24717,n24720,n24721);
  nand U26042(G8515,n24722,n24723,n24724,n24725);
  nor U26043(n24725,n24726,n24727,n24728);
  nor U26044(n24728,G59572,n24720,n22394);
  nand U26045(n24720,G59571,G59570,n24729);
  nor U26046(n24727,n24730,n24721);
  nor U26047(n24730,n24731,n24732);
  nor U26048(n24731,G59571,n22394);
  nor U26049(n24726,n24733,n22401);
  not U26050(n24733,G59763);
  nand U26051(n24724,n22402,n21670);
  nand U26052(n24723,n22403,n21474);
  xor U26053(n21474,n24583,n24734);
  and U26054(n24734,n24582,n24574);
  nand U26055(n24574,n24735,n24736);
  or U26056(n24582,n24736,n24735);
  xnor U26057(n24735,n24737,n22414);
  nand U26058(n24737,n24738,n24739,n24740,n24741);
  nand U26059(n24741,n24742,n24743,n24744,n24745);
  nor U26060(n24745,n24746,n24747,n24748,n24749);
  nor U26061(n24749,n22730,n24428);
  nor U26062(n24748,n23346,n24429);
  nor U26063(n24747,n22722,n24430);
  nand U26064(n24746,n24750,n24751);
  nand U26065(n24751,n24433,G59447);
  nand U26066(n24750,n24434,G59439);
  nor U26067(n24744,n24752,n24753,n24754,n24755);
  nor U26068(n24755,n22729,n24439);
  nor U26069(n24754,n23343,n24440);
  nor U26070(n24753,n23338,n24441);
  nor U26071(n24752,n22719,n24442);
  nor U26072(n24743,n24756,n24757,n24758,n24759);
  nor U26073(n24759,n23345,n24447);
  nor U26074(n24758,n23344,n24448);
  nor U26075(n24757,n22727,n24449);
  nor U26076(n24756,n22728,n24450);
  nor U26077(n24742,n24760,n24761,n24762,n22414);
  nor U26078(n24762,n23336,n24454);
  nor U26079(n24761,n23337,n24455);
  nor U26080(n24760,n23335,n24456);
  nand U26081(n24740,n24457,n23313);
  nand U26082(n23313,n24763,n24764,n24765,n24766);
  nor U26083(n24766,n24767,n24768,n24769,n24770);
  nor U26084(n24770,n23337,n24466);
  nor U26085(n24769,n23336,n24467);
  nor U26086(n24768,n23335,n24468);
  nor U26087(n24767,n23345,n24469);
  nor U26088(n24765,n24771,n24772,n24773,n24774);
  nor U26089(n24774,n23344,n24474);
  nor U26090(n24773,n23343,n24475);
  nor U26091(n24772,n22729,n24476);
  nor U26092(n24771,n22728,n24477);
  nor U26093(n24764,n24775,n24776,n24777,n24778);
  nor U26094(n24778,n22727,n24482);
  nor U26095(n24777,n22721,n24483);
  nor U26096(n24776,n22720,n24484);
  nor U26097(n24775,n22719,n24485);
  nor U26098(n24763,n24779,n24780,n24781,n24782);
  nor U26099(n24782,n23338,n24490);
  nor U26100(n24781,n23346,n24491);
  nor U26101(n24780,n22730,n24492);
  nor U26102(n24779,n22722,n24493);
  nand U26103(n24739,n24531,n24783);
  nand U26104(n24783,n24784,n24785,n24786,n24787);
  nor U26105(n24787,n24788,n24789,n24790,n24791);
  nor U26106(n24791,n23336,n24640);
  nor U26107(n24790,n23335,n24641);
  nor U26108(n24789,n23346,n24642);
  nor U26109(n24788,n23344,n24643);
  nor U26110(n24786,n24792,n24793,n24794,n24795);
  nor U26111(n24795,n23343,n24648);
  nor U26112(n24794,n22730,n24649);
  nor U26113(n24793,n22728,n24650);
  nor U26114(n24792,n22727,n24651);
  nor U26115(n24785,n24796,n24797,n24798,n24799);
  nor U26116(n24799,n22722,n24656);
  nor U26117(n24798,n22720,n24657);
  nor U26118(n24797,n22719,n24658);
  nor U26119(n24796,n23338,n24659);
  nor U26120(n24784,n24800,n24801,n24802,n24803);
  nor U26121(n24803,n23337,n24664);
  nor U26122(n24802,n23345,n24665);
  nor U26123(n24801,n22729,n24666);
  nor U26124(n24800,n22721,n24667);
  nand U26125(n24738,n22473,n24804);
  nand U26126(n24804,n24805,n24806,n24807,n24808);
  nor U26127(n24808,n24809,n24810,n24811,n24812);
  nor U26128(n24812,n23338,n24503);
  nor U26129(n24811,n23337,n24504);
  nor U26130(n24810,n23336,n24505);
  nor U26131(n24809,n23335,n24506);
  nor U26132(n24807,n24813,n24814,n24815,n24816);
  nor U26133(n24816,n23346,n24511);
  nor U26134(n24815,n23345,n24512);
  nor U26135(n24814,n23344,n24513);
  nor U26136(n24813,n23343,n24514);
  nor U26137(n24806,n24817,n24818,n24819,n24820);
  nor U26138(n24820,n22730,n24519);
  nor U26139(n24819,n22729,n24520);
  nor U26140(n24818,n22728,n24521);
  nor U26141(n24817,n22727,n24522);
  nor U26142(n24805,n24821,n24822,n24823,n24824);
  nor U26143(n24824,n22722,n24527);
  nor U26144(n24823,n22721,n24528);
  nor U26145(n24822,n22720,n24529);
  nor U26146(n24821,n22719,n24530);
  nand U26147(n24736,n24825,n24826,n24827,n24828);
  nand U26148(n24828,n21475,n24414);
  nand U26149(n24827,n21670,n22406);
  nand U26150(n24826,G59572,n22438);
  nand U26151(n24825,n22439,G59763);
  nand U26152(n24583,n24829,n24830);
  nand U26153(n24830,n24831,n24832);
  nand U26154(n24831,n24833,n24834);
  or U26155(n24829,n24834,n24833);
  xor U26156(n21475,n24705,n24835);
  nor U26157(n24835,n24836,n24708);
  nor U26158(n24708,n23338,n24706,n21114);
  nor U26159(n24836,n24837,n24838);
  not U26160(n24838,n24706);
  nor U26161(n24706,n24839,n24840);
  and U26162(n24840,n24841,n22383);
  nor U26163(n24839,n24841,n21670,n22383);
  not U26164(n21670,n21471);
  nand U26165(n21471,n24711,n24842);
  nand U26166(n24842,n24843,n24844);
  or U26167(n24711,n24844,n24843);
  xor U26168(n24843,n21108,n24845);
  nor U26169(n24845,n24846,n24847,n24848,n24849);
  and U26170(n24849,n22437,G59699);
  nor U26171(n24848,n22508,n24721);
  not U26172(n24721,G59572);
  nor U26173(n24847,n22383,n22347);
  not U26174(n22347,G59604);
  nor U26175(n24846,n24241,n21472);
  not U26176(n21472,G59731);
  nand U26177(n24844,n24850,n24851);
  nand U26178(n24841,n24852,n24853,n24854);
  nand U26179(n24854,G59604,n23278);
  nand U26180(n24853,G59572,n22496);
  nand U26181(n24852,G59763,n21108);
  nor U26182(n24837,n23338,n21114);
  nand U26183(n24705,n24855,n24856);
  nand U26184(n24856,n24857,n24858);
  nand U26185(G8514,n24859,n24860,n24861,n24862);
  nor U26186(n24862,n24863,n24864,n24865);
  nor U26187(n24865,G59571,n22394,n24866,n24867);
  and U26188(n24864,n24732,G59571);
  nand U26189(n24732,n22456,n24868);
  nand U26190(n24868,n22400,n24869);
  nand U26191(n24869,n24729,G59570);
  nor U26192(n24863,n24870,n22401);
  nand U26193(n24860,n22403,n21486);
  xor U26194(n21486,n24871,n24834);
  xor U26195(n24834,n24872,n22414);
  nand U26196(n24872,n24873,n24874,n24875,n24876);
  nor U26197(n24876,n24877,n24878);
  nor U26198(n24878,n24879,n24880);
  and U26199(n24877,n23389,n24457);
  nand U26200(n23389,n24881,n24882,n24883,n24884);
  nor U26201(n24884,n24885,n24886,n24887,n24888);
  nor U26202(n24888,n23418,n24466);
  nor U26203(n24887,n23417,n24467);
  nor U26204(n24886,n23416,n24468);
  nor U26205(n24885,n23426,n24469);
  nor U26206(n24883,n24889,n24890,n24891,n24892);
  nor U26207(n24892,n23425,n24474);
  nor U26208(n24891,n23424,n24475);
  nor U26209(n24890,n22810,n24476);
  nor U26210(n24889,n22809,n24477);
  nor U26211(n24882,n24893,n24894,n24895,n24896);
  nor U26212(n24896,n22808,n24482);
  nor U26213(n24895,n22802,n24483);
  nor U26214(n24894,n22801,n24484);
  nor U26215(n24893,n22800,n24485);
  nor U26216(n24881,n24897,n24898,n24899,n24900);
  nor U26217(n24900,n23419,n24490);
  nor U26218(n24899,n23427,n24491);
  nor U26219(n24898,n22811,n24492);
  nor U26220(n24897,n22803,n24493);
  nand U26221(n24875,n22473,n24901);
  nand U26222(n24901,n24902,n24903,n24904,n24905);
  nor U26223(n24905,n24906,n24907,n24908,n24909);
  nor U26224(n24909,n23419,n24503);
  nor U26225(n24908,n23418,n24504);
  nor U26226(n24907,n23417,n24505);
  nor U26227(n24906,n23416,n24506);
  nor U26228(n24904,n24910,n24911,n24912,n24913);
  nor U26229(n24913,n23427,n24511);
  nor U26230(n24912,n23426,n24512);
  nor U26231(n24911,n23425,n24513);
  nor U26232(n24910,n23424,n24514);
  nor U26233(n24903,n24914,n24915,n24916,n24917);
  nor U26234(n24917,n22811,n24519);
  nor U26235(n24916,n22810,n24520);
  nor U26236(n24915,n22809,n24521);
  nor U26237(n24914,n22808,n24522);
  nor U26238(n24902,n24918,n24919,n24920,n24921);
  nor U26239(n24921,n22803,n24527);
  nor U26240(n24920,n22802,n24528);
  nor U26241(n24919,n22801,n24529);
  nor U26242(n24918,n22800,n24530);
  nand U26243(n24874,n24922,n24923,n24924,n24925);
  nor U26244(n24925,n24926,n24927,n24928,n24929);
  nor U26245(n24929,n22811,n24428);
  nor U26246(n24928,n23427,n24429);
  nor U26247(n24927,n22803,n24430);
  nand U26248(n24926,n24930,n24931);
  nand U26249(n24931,n24433,G59448);
  nand U26250(n24930,n24434,G59440);
  nor U26251(n24924,n24932,n24933,n24934,n24935);
  nor U26252(n24935,n22810,n24439);
  nor U26253(n24934,n23424,n24440);
  nor U26254(n24933,n23419,n24441);
  nor U26255(n24932,n22800,n24442);
  nor U26256(n24923,n24936,n24937,n24938,n24939);
  nor U26257(n24939,n23426,n24447);
  nor U26258(n24938,n23425,n24448);
  nor U26259(n24937,n22808,n24449);
  nor U26260(n24936,n22809,n24450);
  nor U26261(n24922,n24940,n24941,n24942,n22414);
  nor U26262(n24942,n23417,n24454);
  nor U26263(n24941,n23418,n24455);
  nor U26264(n24940,n23416,n24456);
  nand U26265(n24873,n24531,n24943);
  nand U26266(n24943,n24944,n24945,n24946,n24947);
  nor U26267(n24947,n24948,n24949,n24950,n24951);
  nor U26268(n24951,n23417,n24640);
  nor U26269(n24950,n23416,n24641);
  nor U26270(n24949,n23427,n24642);
  nor U26271(n24948,n23425,n24643);
  nor U26272(n24946,n24952,n24953,n24954,n24955);
  nor U26273(n24955,n23424,n24648);
  nor U26274(n24954,n22811,n24649);
  nor U26275(n24953,n22809,n24650);
  nor U26276(n24952,n22808,n24651);
  nor U26277(n24945,n24956,n24957,n24958,n24959);
  nor U26278(n24959,n22803,n24656);
  nor U26279(n24958,n22801,n24657);
  nor U26280(n24957,n22800,n24658);
  nor U26281(n24956,n23419,n24659);
  nor U26282(n24944,n24960,n24961,n24962,n24963);
  nor U26283(n24963,n23418,n24664);
  nor U26284(n24962,n23426,n24665);
  nor U26285(n24961,n22810,n24666);
  nor U26286(n24960,n22802,n24667);
  xor U26287(n24871,n24832,n24833);
  and U26288(n24833,n24964,n24965,n24966,n24967);
  nand U26289(n24967,n20986,n24414);
  nand U26290(n24966,G59571,n22438);
  nand U26291(n24965,n22406,n21674);
  nand U26292(n24964,n22439,G59762);
  nand U26293(n24832,n24968,n24969);
  nand U26294(n24969,n24970,n24971);
  nand U26295(n24859,n22402,n21674);
  nand U26296(G8513,n24972,n24973,n24974,n24975);
  nor U26297(n24975,n24976,n24977,n24978);
  nor U26298(n24978,G59570,n24867,n22394);
  nor U26299(n24977,n24979,n24866);
  nor U26300(n24979,n24980,n22399);
  nor U26301(n24980,n24729,n22394);
  not U26302(n24729,n24867);
  nand U26303(n24867,n21058,n24981);
  nand U26304(n24981,n24982,n24983);
  nor U26305(n24976,n21497,n22401);
  nand U26306(n24973,n22403,n21499);
  xor U26307(n21499,n24971,n24984);
  and U26308(n24984,n24968,n24970);
  or U26309(n24970,n24985,n24986);
  nand U26310(n24968,n24986,n24985);
  nand U26311(n24985,n24987,n24988,n24989,n24990);
  nand U26312(n24990,n20996,n24414);
  nand U26313(n24989,G59570,n22438);
  nand U26314(n24988,n22406,n21498);
  nand U26315(n24987,n22439,G59761);
  xnor U26316(n24986,n22414,n24991);
  nand U26317(n24991,n24992,n24993,n24994,n24995);
  nor U26318(n24995,n24996,n24997);
  nor U26319(n24997,n24879,n24998);
  nor U26320(n24996,n24999,n21935);
  nor U26321(n24999,n25000,n25001,n25002,n25003);
  nand U26322(n25003,n25004,n25005,n25006,n25007);
  nand U26323(n25007,n25008,G59433);
  nand U26324(n25006,n25009,G59441);
  nand U26325(n25005,n25010,G59449);
  nand U26326(n25004,n25011,G59457);
  nand U26327(n25002,n25012,n25013,n25014,n25015);
  nand U26328(n25015,n25016,G59465);
  nand U26329(n25014,n25017,G59473);
  nand U26330(n25013,n25018,G59481);
  nand U26331(n25012,n25019,G59489);
  nand U26332(n25001,n25020,n25021,n25022,n25023);
  nand U26333(n25023,n25024,G59497);
  nand U26334(n25022,n25025,G59505);
  nand U26335(n25021,n25026,G59513);
  nand U26336(n25020,n25027,G59521);
  nand U26337(n25000,n25028,n25029,n25030,n25031);
  nand U26338(n25031,n25032,G59529);
  nand U26339(n25030,n25033,G59537);
  nand U26340(n25029,n25034,G59545);
  nand U26341(n25028,n25035,G59553);
  nand U26342(n24994,n24457,n23473);
  nand U26343(n23473,n25036,n25037,n25038,n25039);
  nor U26344(n25039,n25040,n25041,n25042,n25043);
  nor U26345(n25043,n23502,n24466);
  nor U26346(n25042,n23501,n24467);
  nor U26347(n25041,n23500,n24468);
  nor U26348(n25040,n23510,n24469);
  nor U26349(n25038,n25044,n25045,n25046,n25047);
  nor U26350(n25047,n23509,n24474);
  nor U26351(n25046,n23508,n24475);
  nor U26352(n25045,n22884,n24476);
  nor U26353(n25044,n22883,n24477);
  nor U26354(n25037,n25048,n25049,n25050,n25051);
  nor U26355(n25051,n22882,n24482);
  nor U26356(n25050,n22876,n24483);
  nor U26357(n25049,n22875,n24484);
  nor U26358(n25048,n22874,n24485);
  nor U26359(n25036,n25052,n25053,n25054,n25055);
  nor U26360(n25055,n23503,n24490);
  nor U26361(n25054,n23511,n24491);
  nor U26362(n25053,n22885,n24492);
  nor U26363(n25052,n22877,n24493);
  nand U26364(n24993,n25056,n25057,n25058,n25059);
  nor U26365(n25059,n25060,n25061,n25062,n25063);
  nor U26366(n25063,n22885,n24428);
  nor U26367(n25062,n23511,n24429);
  nor U26368(n25061,n22877,n24430);
  nand U26369(n25060,n25064,n25065);
  nand U26370(n25065,n24433,G59449);
  nand U26371(n25064,n24434,G59441);
  nor U26372(n25058,n25066,n25067,n25068,n25069);
  nor U26373(n25069,n22884,n24439);
  nor U26374(n25068,n23508,n24440);
  nor U26375(n25067,n23503,n24441);
  nor U26376(n25066,n22874,n24442);
  nor U26377(n25057,n25070,n25071,n25072,n25073);
  nor U26378(n25073,n23510,n24447);
  nor U26379(n25072,n23509,n24448);
  nor U26380(n25071,n22882,n24449);
  nor U26381(n25070,n22883,n24450);
  nor U26382(n25056,n25074,n25075,n25076,n22414);
  nor U26383(n25076,n23501,n24454);
  nor U26384(n25075,n23502,n24455);
  nor U26385(n25074,n23500,n24456);
  nand U26386(n24992,n24531,n25077);
  nand U26387(n25077,n25078,n25079,n25080,n25081);
  nor U26388(n25081,n25082,n25083,n25084,n25085);
  nor U26389(n25085,n23501,n24640);
  nor U26390(n25084,n23500,n24641);
  nor U26391(n25083,n23511,n24642);
  nor U26392(n25082,n23509,n24643);
  nor U26393(n25080,n25086,n25087,n25088,n25089);
  nor U26394(n25089,n23508,n24648);
  nor U26395(n25088,n22885,n24649);
  nor U26396(n25087,n22883,n24650);
  nor U26397(n25086,n22882,n24651);
  nor U26398(n25079,n25090,n25091,n25092,n25093);
  nor U26399(n25093,n22877,n24656);
  nor U26400(n25092,n22875,n24657);
  nor U26401(n25091,n22874,n24658);
  nor U26402(n25090,n23503,n24659);
  nor U26403(n25078,n25094,n25095,n25096,n25097);
  nor U26404(n25097,n23502,n24664);
  nor U26405(n25096,n23510,n24665);
  nor U26406(n25095,n22884,n24666);
  nor U26407(n25094,n22876,n24667);
  nand U26408(n24971,n25098,n25099);
  nand U26409(n25099,n25100,n25101);
  nand U26410(n24972,n22402,n21498);
  nand U26411(G8512,n25102,n25103,n25104,n25105);
  nor U26412(n25105,n25106,n25107,n25108);
  and U26413(n25108,n24982,n24983,n22400);
  not U26414(n22400,n22394);
  nor U26415(n25107,n25109,n24982);
  nor U26416(n25109,n25110,n22399);
  nor U26417(n25110,n22394,n24983);
  nand U26418(n24983,G59567,n21058,G59568);
  nor U26419(n25106,n21509,n22401);
  not U26420(n21509,G59760);
  nand U26421(n25103,n22403,n21511);
  xor U26422(n21511,n25100,n25111);
  and U26423(n25111,n25101,n25098);
  nand U26424(n25098,n25112,n25113);
  nand U26425(n25113,n25114,n25115);
  nand U26426(n25101,n25114,n25115,n25116);
  not U26427(n25116,n25112);
  nand U26428(n25112,n25117,n25118,n25119,n25120);
  nand U26429(n25120,n21006,n24414);
  nand U26430(n24414,n22750,n21935);
  nand U26431(n25119,G59569,n22438);
  not U26432(n22438,n22470);
  nand U26433(n25118,n22406,n21510);
  nand U26434(n25117,n22439,G59760);
  not U26435(n22439,n22469);
  nand U26436(n25115,n22406,n25121,n25122);
  nand U26437(n25121,n25123,n25124,n25125,n25126);
  nor U26438(n25126,n25127,n25128,n25129,n25130);
  nor U26439(n25130,n22955,n25131);
  nor U26440(n25129,n22956,n24430);
  nor U26441(n25128,n22964,n24428);
  nor U26442(n25127,n23596,n24429);
  nor U26443(n25125,n25132,n25133,n25134,n25135);
  nor U26444(n25135,n23593,n24440);
  nor U26445(n25134,n23588,n24441);
  nor U26446(n25133,n22953,n24442);
  nor U26447(n25132,n22954,n25136);
  nor U26448(n25124,n25137,n25138,n25139,n25140);
  nor U26449(n25140,n23594,n24448);
  nor U26450(n25139,n22961,n24449);
  nor U26451(n25138,n22962,n24450);
  nor U26452(n25137,n22963,n24439);
  nor U26453(n25123,n25141,n25142,n25143,n25144);
  nor U26454(n25144,n23586,n24454);
  nor U26455(n25143,n23587,n24455);
  nor U26456(n25142,n23585,n24456);
  nor U26457(n25141,n23595,n24447);
  nand U26458(n25114,n25145,n22414);
  nand U26459(n25145,n25122,n25146,n25147,n25148);
  nand U26460(n25147,n24531,n25149);
  nand U26461(n25149,n25150,n25151,n25152,n25153);
  nor U26462(n25153,n25154,n25155,n25156,n25157);
  nor U26463(n25157,n23586,n24640);
  nor U26464(n25156,n23585,n24641);
  nor U26465(n25155,n23596,n24642);
  nor U26466(n25154,n23594,n24643);
  nor U26467(n25152,n25158,n25159,n25160,n25161);
  nor U26468(n25161,n23593,n24648);
  nor U26469(n25160,n22964,n24649);
  nor U26470(n25159,n22962,n24650);
  nor U26471(n25158,n22961,n24651);
  nor U26472(n25151,n25162,n25163,n25164,n25165);
  nor U26473(n25165,n22956,n24656);
  nor U26474(n25164,n22954,n24657);
  nor U26475(n25163,n22953,n24658);
  nor U26476(n25162,n23588,n24659);
  nor U26477(n25150,n25166,n25167,n25168,n25169);
  nor U26478(n25169,n23587,n24664);
  nor U26479(n25168,n23595,n24665);
  nor U26480(n25167,n22963,n24666);
  nor U26481(n25166,n22955,n24667);
  nand U26482(n25146,n24457,n23558);
  nand U26483(n23558,n25170,n25171,n25172,n25173);
  nor U26484(n25173,n25174,n25175,n25176,n25177);
  nor U26485(n25177,n23587,n24466);
  nor U26486(n25176,n23586,n24467);
  nor U26487(n25175,n23585,n24468);
  nor U26488(n25174,n23595,n24469);
  nor U26489(n25172,n25178,n25179,n25180,n25181);
  nor U26490(n25181,n23594,n24474);
  nor U26491(n25180,n23593,n24475);
  nor U26492(n25179,n22963,n24476);
  nor U26493(n25178,n22962,n24477);
  nor U26494(n25171,n25182,n25183,n25184,n25185);
  nor U26495(n25185,n22961,n24482);
  nor U26496(n25184,n22955,n24483);
  nor U26497(n25183,n22954,n24484);
  nor U26498(n25182,n22953,n24485);
  nor U26499(n25170,n25186,n25187,n25188,n25189);
  nor U26500(n25189,n23588,n24490);
  nor U26501(n25188,n23596,n24491);
  nor U26502(n25187,n22964,n24492);
  nor U26503(n25186,n22956,n24493);
  and U26504(n25122,n25190,n25191);
  nand U26505(n25191,n22473,n25192);
  nand U26506(n25192,n25193,n25194,n25195,n25196);
  nor U26507(n25196,n25197,n25198,n25199,n25200);
  nor U26508(n25200,n23588,n24503);
  nor U26509(n25199,n23587,n24504);
  nor U26510(n25198,n23586,n24505);
  nor U26511(n25197,n23585,n24506);
  nor U26512(n25195,n25201,n25202,n25203,n25204);
  nor U26513(n25204,n23596,n24511);
  nor U26514(n25203,n23595,n24512);
  nor U26515(n25202,n23594,n24513);
  nor U26516(n25201,n23593,n24514);
  nor U26517(n25194,n25205,n25206,n25207,n25208);
  nor U26518(n25208,n22964,n24519);
  nor U26519(n25207,n22963,n24520);
  nor U26520(n25206,n22962,n24521);
  nor U26521(n25205,n22961,n24522);
  nor U26522(n25193,n25209,n25210,n25211,n25212);
  nor U26523(n25212,n22956,n24527);
  nor U26524(n25211,n22955,n24528);
  nor U26525(n25210,n22954,n24529);
  nor U26526(n25209,n22953,n24530);
  nand U26527(n25190,G59559,n21849);
  nand U26528(n25100,n25213,n25214);
  nand U26529(n25214,n25215,n25216);
  nand U26530(n25102,n22402,n21510);
  nand U26531(G8511,n25217,n25218,n25219,n25220);
  nor U26532(n25220,n25221,n25222,n25223);
  nor U26533(n25223,G59568,n25224,n22394);
  nor U26534(n25222,n25225,n25226);
  nor U26535(n25225,n25227,n22399);
  nor U26536(n25221,n21130,n22401);
  nand U26537(n25218,n22403,n21522);
  xor U26538(n21522,n25216,n25228);
  and U26539(n25228,n25215,n25213);
  or U26540(n25213,n25229,n25230);
  nand U26541(n25215,n25230,n25229);
  xor U26542(n25229,n25231,n22414);
  nand U26543(n25231,n25232,n25233,n25234,n25235);
  nor U26544(n25235,n25236,n25237,n25238,n25239);
  nor U26545(n25239,n25240,n21935);
  nor U26546(n25240,n25241,n25242,n25243,n25244);
  nand U26547(n25244,n25245,n25246,n25247,n25248);
  nand U26548(n25248,n25008,G59435);
  nand U26549(n25247,n25009,G59443);
  nand U26550(n25246,n25010,G59451);
  nand U26551(n25245,n25011,G59459);
  nand U26552(n25243,n25249,n25250,n25251,n25252);
  nand U26553(n25252,n25016,G59467);
  nand U26554(n25251,n25017,G59475);
  nand U26555(n25250,n25018,G59483);
  nand U26556(n25249,n25019,G59491);
  nand U26557(n25242,n25253,n25254,n25255,n25256);
  nand U26558(n25256,n25024,G59499);
  nand U26559(n25255,n25025,G59507);
  nand U26560(n25254,n25026,G59515);
  nand U26561(n25253,n25027,G59523);
  nand U26562(n25241,n25257,n25258,n25259,n25260);
  nand U26563(n25260,n25032,G59531);
  nand U26564(n25259,n25033,G59539);
  nand U26565(n25258,n25034,G59547);
  nand U26566(n25257,n25035,G59555);
  nor U26567(n25238,n25261,n25262,n25263,n25264);
  nand U26568(n25264,n22406,n25265,n25266,n25267);
  nand U26569(n25267,n25268,G59523);
  nand U26570(n25266,n25269,G59491);
  nand U26571(n25265,n25270,G59459);
  nand U26572(n25263,n25271,n25272,n25273,n25274);
  nand U26573(n25274,n24433,G59451);
  nand U26574(n25273,n24434,G59443);
  nand U26575(n25272,n25275,G59435);
  nand U26576(n25271,n25276,G59555);
  nand U26577(n25262,n25277,n25278,n25279,n25280);
  nand U26578(n25280,n25281,G59499);
  nand U26579(n25279,n25282,G59483);
  nand U26580(n25278,n25283,G59475);
  nand U26581(n25277,n25284,G59467);
  nand U26582(n25261,n25285,n25286,n25287,n25288);
  nor U26583(n25288,n25289,n25290);
  nor U26584(n25290,n23048,n24454);
  nor U26585(n25289,n23049,n24455);
  nand U26586(n25287,n25291,G59531);
  nand U26587(n25286,n25292,G59507);
  nand U26588(n25285,n25293,G59515);
  nand U26589(n25234,G59560,n21849);
  nand U26590(n25233,n24531,n25294);
  nand U26591(n25294,n25295,n25296,n25297,n25298);
  nor U26592(n25298,n25299,n25300,n25301,n25302);
  nor U26593(n25302,n23048,n24640);
  nor U26594(n25301,n23047,n24641);
  nor U26595(n25300,n23042,n24642);
  nor U26596(n25299,n23040,n24643);
  nor U26597(n25297,n25303,n25304,n25305,n25306);
  nor U26598(n25306,n23039,n24648);
  nor U26599(n25305,n23034,n24649);
  nor U26600(n25304,n23032,n24650);
  nor U26601(n25303,n23031,n24651);
  nor U26602(n25296,n25307,n25308,n25309,n25310);
  nor U26603(n25310,n23026,n24656);
  nor U26604(n25309,n23024,n24657);
  nor U26605(n25308,n23023,n24658);
  nor U26606(n25307,n23050,n24659);
  nor U26607(n25295,n25311,n25312,n25313,n25314);
  nor U26608(n25314,n23049,n24664);
  nor U26609(n25313,n23041,n24665);
  nor U26610(n25312,n23033,n24666);
  nor U26611(n25311,n23025,n24667);
  nand U26612(n25232,n24457,n23640);
  nand U26613(n23640,n25315,n25316,n25317,n25318);
  nor U26614(n25318,n25319,n25320,n25321,n25322);
  nor U26615(n25322,n23049,n24466);
  nor U26616(n25321,n23048,n24467);
  nor U26617(n25320,n23047,n24468);
  nor U26618(n25319,n23041,n24469);
  nor U26619(n25317,n25323,n25324,n25325,n25326);
  nor U26620(n25326,n23040,n24474);
  nor U26621(n25325,n23039,n24475);
  nor U26622(n25324,n23033,n24476);
  nor U26623(n25323,n23032,n24477);
  nor U26624(n25316,n25327,n25328,n25329,n25330);
  nor U26625(n25330,n23031,n24482);
  nor U26626(n25329,n23025,n24483);
  nor U26627(n25328,n23024,n24484);
  nor U26628(n25327,n23023,n24485);
  nor U26629(n25315,n25331,n25332,n25333,n25334);
  nor U26630(n25334,n23050,n24490);
  nor U26631(n25333,n23042,n24491);
  nor U26632(n25332,n23034,n24492);
  nor U26633(n25331,n23026,n24493);
  and U26634(n25230,n25335,n25336,n25337,n25338);
  nand U26635(n25338,n21015,n22473);
  nor U26636(n25337,n25339,n25340);
  nor U26637(n25340,n21130,n22469);
  nor U26638(n25339,n22470,n25226);
  nand U26639(n25336,n22406,n21521);
  nand U26640(n25335,n21015,n22423);
  nand U26641(n25216,n25341,n25342);
  nand U26642(n25342,n22406,n25343);
  nand U26643(n25343,n25344,n25345);
  not U26644(n25344,n25346);
  nand U26645(n25217,n22402,n21521);
  nand U26646(G8510,n25347,n25348,n25349,n25350);
  nor U26647(n25350,n25351,n25227,n25352);
  nor U26648(n25352,n25224,n22456);
  nor U26649(n25227,G59567,n22394);
  nand U26650(n22394,n25353,n25354);
  nor U26651(n25351,n21122,n22401);
  nand U26652(n25349,n22403,n21546);
  xnor U26653(n21546,n22414,n25355);
  nor U26654(n25355,n25356,n25357);
  not U26655(n25357,n25341);
  nand U26656(n25341,n25358,n25346);
  nor U26657(n25356,n25358,n25346);
  nand U26658(n25346,n25359,n25360,n24879,n25361);
  nor U26659(n25361,n25362,n25363,n25364);
  nor U26660(n25364,n21122,n22469);
  nand U26661(n22469,n25365,n21846,n25366);
  nor U26662(n25363,n21532,n21935);
  nor U26663(n25362,n22470,n25224);
  nand U26664(n25360,n22406,n21084);
  nand U26665(n25359,n21030,n22423);
  not U26666(n22423,n22750);
  nor U26667(n22750,n24531,n24457);
  xnor U26668(n25358,n25345,n22414);
  nand U26669(n25345,n25369,n25370,n25371,n25372);
  nor U26670(n25372,n25367,n25368,n25373,n25374);
  nor U26671(n25374,n25375,n21935);
  nor U26672(n25375,n25376,n25377,n25378,n25379);
  nand U26673(n25379,n25380,n25381,n25382,n25383);
  nand U26674(n25383,n25008,G59436);
  not U26675(n25008,n24530);
  nand U26676(n24530,n25384,n25385);
  nand U26677(n25382,n25009,G59444);
  not U26678(n25009,n24529);
  nand U26679(n24529,n25384,n25386);
  nand U26680(n25381,n25010,G59452);
  not U26681(n25010,n24528);
  nand U26682(n24528,n25387,n25385);
  nand U26683(n25380,n25011,G59460);
  not U26684(n25011,n24527);
  nand U26685(n24527,n25387,n25386);
  nand U26686(n25378,n25388,n25389,n25390,n25391);
  nand U26687(n25391,n25016,G59468);
  not U26688(n25016,n24522);
  nand U26689(n24522,n25384,n25392);
  nand U26690(n25390,n25017,G59476);
  not U26691(n25017,n24521);
  nand U26692(n24521,n25384,n25393);
  nor U26693(n25384,n25394,n25395);
  nand U26694(n25389,n25018,G59484);
  not U26695(n25018,n24520);
  nand U26696(n24520,n25387,n25392);
  nand U26697(n25388,n25019,G59492);
  not U26698(n25019,n24519);
  nand U26699(n24519,n25387,n25393);
  nor U26700(n25387,n25396,n25394);
  nand U26701(n25377,n25397,n25398,n25399,n25400);
  nand U26702(n25400,n25024,G59500);
  not U26703(n25024,n24514);
  nand U26704(n24514,n25385,n25401);
  nand U26705(n25399,n25025,G59508);
  not U26706(n25025,n24513);
  nand U26707(n24513,n25386,n25401);
  nand U26708(n25398,n25026,G59516);
  not U26709(n25026,n24512);
  nand U26710(n24512,n25385,n25402);
  nor U26711(n25385,n25403,G59561);
  nand U26712(n25397,n25027,G59524);
  not U26713(n25027,n24511);
  nand U26714(n24511,n25386,n25402);
  nor U26715(n25386,n25403,n23142);
  nand U26716(n25376,n25404,n25405,n25406,n25407);
  nand U26717(n25407,n25032,G59532);
  not U26718(n25032,n24506);
  nand U26719(n24506,n25392,n25401);
  nand U26720(n25406,n25033,G59540);
  not U26721(n25033,n24505);
  nand U26722(n24505,n25393,n25401);
  and U26723(n25401,n25396,n25394);
  not U26724(n25396,n25395);
  nand U26725(n25405,n25034,G59548);
  not U26726(n25034,n24504);
  nand U26727(n24504,n25402,n25392);
  and U26728(n25392,n25403,n23142);
  nand U26729(n25404,n25035,G59556);
  not U26730(n25035,n24503);
  nand U26731(n24503,n25402,n25393);
  and U26732(n25393,G59561,n25403);
  and U26733(n25402,n25395,n25394);
  nor U26734(n25373,n25408,n25409,n25410,n25411);
  nand U26735(n25411,n22406,n25412,n25413,n25414);
  nand U26736(n25414,n25268,G59524);
  not U26737(n25268,n24429);
  nand U26738(n24429,n25415,n25416);
  nand U26739(n25413,n25269,G59492);
  not U26740(n25269,n24428);
  nand U26741(n24428,n25417,n25418);
  nand U26742(n25412,n25270,G59460);
  not U26743(n25270,n24430);
  nand U26744(n24430,n25418,n25416);
  nand U26745(n25410,n25419,n25420,n25421,n25422);
  nand U26746(n25422,n24433,G59452);
  not U26747(n24433,n25131);
  nand U26748(n25131,n25423,n25418);
  nand U26749(n25421,n24434,G59444);
  not U26750(n24434,n25136);
  nand U26751(n25136,n25424,n25416);
  nand U26752(n25420,n25275,G59436);
  not U26753(n25275,n24442);
  nand U26754(n24442,n25424,n25423);
  nand U26755(n25419,n25276,G59556);
  not U26756(n25276,n24441);
  nand U26757(n24441,n25417,n25415);
  nand U26758(n25409,n25425,n25426,n25427,n25428);
  nand U26759(n25428,n25281,G59500);
  not U26760(n25281,n24440);
  nand U26761(n24440,n25429,n25423);
  nand U26762(n25427,n25282,G59484);
  not U26763(n25282,n24439);
  nand U26764(n24439,n25430,n25418);
  nor U26765(n25418,n21496,n21015);
  nand U26766(n25426,n25283,G59476);
  not U26767(n25283,n24450);
  nand U26768(n24450,n25424,n25417);
  nand U26769(n25425,n25284,G59468);
  not U26770(n25284,n24449);
  nand U26771(n24449,n25430,n25424);
  nor U26772(n25424,n21520,n21496);
  not U26773(n21496,n20996);
  nand U26774(n25408,n25431,n25432,n25433,n25434);
  nor U26775(n25434,n25435,n25436);
  nor U26776(n25436,n23144,n24454);
  nand U26777(n24454,n25429,n25417);
  nor U26778(n25417,n21030,n21006);
  nor U26779(n25435,n23145,n24455);
  nand U26780(n24455,n25430,n25415);
  nand U26781(n25433,n25291,G59532);
  not U26782(n25291,n24456);
  nand U26783(n24456,n25430,n25429);
  nor U26784(n25430,n21532,n21006);
  nand U26785(n25432,n25292,G59508);
  not U26786(n25292,n24448);
  nand U26787(n24448,n25429,n25416);
  nor U26788(n25416,n21030,n21508);
  nor U26789(n25429,n21520,n20996);
  nand U26790(n25431,n25293,G59516);
  not U26791(n25293,n24447);
  nand U26792(n24447,n25423,n25415);
  nor U26793(n25415,n21015,n20996);
  nor U26794(n25423,n21508,n21532);
  not U26795(n21532,n21030);
  nand U26796(n25371,G59561,n21849);
  nand U26797(n25370,n24531,n25437);
  nand U26798(n25437,n25438,n25439,n25440,n25441);
  nor U26799(n25441,n25442,n25443,n25444,n25445);
  nor U26800(n25445,n23144,n24640);
  nor U26801(n25444,n23140,n24641);
  nor U26802(n25443,n23135,n24642);
  nor U26803(n25442,n23133,n24643);
  nor U26804(n25440,n25446,n25447,n25448,n25449);
  nor U26805(n25449,n23131,n24648);
  nor U26806(n25448,n23125,n24649);
  nor U26807(n25447,n23123,n24650);
  nor U26808(n25446,n23121,n24651);
  nor U26809(n25439,n25450,n25451,n25452,n25453);
  nor U26810(n25453,n23113,n24656);
  nor U26811(n25452,n23109,n24657);
  nor U26812(n25451,n23106,n24658);
  nor U26813(n25450,n23147,n24659);
  nor U26814(n25438,n25454,n25455,n25456,n25457);
  nor U26815(n25457,n23145,n24664);
  nor U26816(n25456,n23134,n24665);
  nor U26817(n25455,n23124,n24666);
  nor U26818(n25454,n23111,n24667);
  nand U26819(n25369,n24457,n23720);
  nand U26820(n23720,n25458,n25459,n25460,n25461);
  nor U26821(n25461,n25462,n25463,n25464,n25465);
  nor U26822(n25465,n23145,n24466);
  nand U26823(n24466,n25466,n25467);
  nor U26824(n25464,n23144,n24467);
  nand U26825(n24467,n25468,n25466);
  nor U26826(n25463,n23140,n24468);
  nand U26827(n24468,n25466,n25469);
  nor U26828(n25462,n23134,n24469);
  nand U26829(n24469,n25470,n25467);
  nor U26830(n25460,n25471,n25472,n25473,n25474);
  nor U26831(n25474,n23133,n24474);
  nand U26832(n24474,n25468,n25470);
  nor U26833(n25473,n23131,n24475);
  nand U26834(n24475,n25469,n25470);
  nor U26835(n25472,n23124,n24476);
  nand U26836(n24476,n25475,n25467);
  nor U26837(n25471,n23123,n24477);
  nand U26838(n24477,n25475,n25468);
  nor U26839(n25459,n25476,n25477,n25478,n25479);
  nor U26840(n25479,n23121,n24482);
  nand U26841(n24482,n25475,n25469);
  nor U26842(n25478,n23111,n24483);
  nand U26843(n24483,n25480,n25467);
  nor U26844(n25467,n25481,n21521);
  nor U26845(n25477,n23109,n24484);
  nand U26846(n24484,n25480,n25468);
  nor U26847(n25468,n21084,n22375);
  nor U26848(n25476,n23106,n24485);
  nand U26849(n24485,n25480,n25469);
  nor U26850(n25469,n22375,n25481);
  nor U26851(n25458,n25482,n25483,n25484,n25485);
  nor U26852(n25485,n23147,n24490);
  nand U26853(n24490,n25486,n25466);
  nor U26854(n25466,n21510,n21498);
  nor U26855(n25484,n23135,n24491);
  nand U26856(n24491,n25486,n25470);
  nor U26857(n25470,n22368,n21498);
  nor U26858(n25483,n23125,n24492);
  nand U26859(n24492,n25486,n25475);
  nor U26860(n25475,n22361,n21510);
  nor U26861(n25482,n23113,n24493);
  nand U26862(n24493,n25486,n25480);
  nor U26863(n25480,n22368,n22361);
  nor U26864(n25486,n21084,n21521);
  nor U26865(n24457,n21031,n22163,n25487);
  nand U26866(n25488,n25489,n25490,n25491,n25492);
  nand U26867(n25348,n22402,n21084);
  not U26868(n22402,n22975);
  nand U26869(n22975,n25353,n25493);
  nand U26870(n25493,n25494,n25495,n25496,n25497);
  nand U26871(n25347,n22440,n21030);
  not U26872(n22440,n23868);
  nand U26873(n23868,n25353,n25498);
  nand U26874(n25498,n25499,n25500,n25501,n25502);
  nor U26875(n25502,n25503,n25504);
  not U26876(n25500,n25505);
  nor U26877(n25353,n21044,n22399);
  not U26878(n22399,n22456);
  nand U26879(n22456,n21553,n25506);
  nand U26880(n25506,n21022,n25507);
  nand U26881(n25507,n25508,n25509,n25510,n25511);
  nand U26882(n25511,n24879,n21534,n25512);
  nand U26883(n25510,n25513,n21045);
  nand U26884(n25513,n25514,n25515);
  nand U26885(n25515,n25512,n25516,n25517);
  nand U26886(n25514,n25518,n21080);
  nand U26887(n25518,n25519,n25520);
  nand U26888(n25520,n25521,n21849);
  nand U26889(n25521,n21057,n21059);
  nand U26890(n25519,n25366,n21060);
  nand U26891(n25509,n21080,n25522);
  nand U26892(n21553,n21043,n21531,n21075);
  nand U26893(G8509,n25523,n25524,n25525);
  nand U26894(n25525,n21082,G59565);
  nand U26895(n25524,n21083,n21521);
  nand U26896(n25523,n21085,n21014);
  nand U26897(G8508,n25526,n25527,n25528);
  nand U26898(n25528,n21082,G59564);
  nand U26899(n25527,n21083,n21510);
  nand U26900(n25526,n21085,n21005);
  nand U26901(G8507,n25529,n25530,n25531);
  nand U26902(n25531,n21082,G59563);
  nand U26903(n25530,n21083,n21498);
  and U26904(n21083,n25532,n21081);
  nand U26905(n25532,n25533,n25534);
  nand U26906(n25534,n22383,n21044);
  nand U26907(n25529,n21085,n25535);
  nor U26908(n21085,n21082,G59426,n22383);
  not U26909(n21082,n21081);
  nor U26910(G8506,n25536,n21081);
  nand U26911(n21081,n25537,n21020,n25538);
  nand U26912(n21020,G59795,n25539);
  nand U26913(n25537,n21031,n25539);
  nand U26914(G8505,n25540,n25541,n25542,n25543);
  nor U26915(n25543,n25544,n25545,n25546);
  nor U26916(n25546,n21848,n25547);
  nor U26917(n25545,n25548,n25549);
  nor U26918(n25544,n23169,n25550);
  nand U26919(n25542,n25551,G59556);
  nand U26920(n25541,n25552,n25553);
  nand U26921(n25540,n21932,n25554);
  nand U26922(G8504,n25555,n25556,n25557,n25558);
  nor U26923(n25558,n25559,n25560,n25561);
  nor U26924(n25561,n21838,n25547);
  nor U26925(n25560,n25562,n25549);
  nor U26926(n25559,n23169,n25563);
  nand U26927(n25557,n25551,G59555);
  nand U26928(n25556,n25564,n25553);
  nand U26929(n25555,n21927,n25554);
  nand U26930(G8503,n25565,n25566,n25567,n25568);
  nor U26931(n25568,n25569,n25570,n25571);
  nor U26932(n25571,n21830,n25547);
  nor U26933(n25570,n25572,n25549);
  nor U26934(n25569,n23169,n25573);
  nand U26935(n25567,n25551,G59554);
  nand U26936(n25566,n25574,n25553);
  nand U26937(n25565,n21922,n25554);
  nand U26938(G8502,n25575,n25576,n25577,n25578);
  nor U26939(n25578,n25579,n25580,n25581);
  nor U26940(n25581,n21822,n25547);
  nor U26941(n25580,n25582,n25549);
  nor U26942(n25579,n23169,n25583);
  nand U26943(n25577,n25551,G59553);
  nand U26944(n25576,n25584,n25553);
  nand U26945(n25575,n21917,n25554);
  nand U26946(G8501,n25585,n25586,n25587,n25588);
  nor U26947(n25588,n25589,n25590,n25591);
  nor U26948(n25591,n21813,n25547);
  nor U26949(n25590,n25592,n25549);
  nor U26950(n25589,n23169,n25593);
  nand U26951(n25587,n25551,G59552);
  nand U26952(n25586,n25594,n25553);
  nand U26953(n25585,n21912,n25554);
  nand U26954(G8500,n25595,n25596,n25597,n25598);
  nor U26955(n25598,n25599,n25600,n25601);
  nor U26956(n25601,n21804,n25547);
  nor U26957(n25600,n25602,n25549);
  nor U26958(n25599,n23169,n25603);
  nand U26959(n25597,n25551,G59551);
  nand U26960(n25596,n25604,n25553);
  nand U26961(n25595,n21907,n25554);
  nand U26962(G8499,n25605,n25606,n25607,n25608);
  nor U26963(n25608,n25609,n25610,n25611);
  nor U26964(n25611,n21795,n25547);
  nor U26965(n25610,n25612,n25549);
  nor U26966(n25609,n23169,n25613);
  nand U26967(n25607,n25551,G59550);
  nand U26968(n25606,n25614,n25553);
  nand U26969(n25605,n21901,n25554);
  nand U26970(G8498,n25615,n25616,n25617,n25618);
  nor U26971(n25618,n25619,n25620,n25621);
  nor U26972(n25621,n21785,n25547);
  nand U26973(n25547,n25622,n23169,n25623);
  nor U26974(n25620,n25624,n25549);
  nor U26975(n25619,n23169,n25625);
  nand U26976(n25617,n25551,G59549);
  and U26977(n25551,n25626,n25627);
  nand U26978(n25627,n25628,n25629,n25630);
  nand U26979(n25630,G59426,n24659);
  nand U26980(n25628,n25631,n25632);
  nand U26981(n25626,n25633,n25634);
  nand U26982(n25616,n25635,n25553);
  nand U26983(n25553,n25636,n25637);
  or U26984(n25637,n25632,n22383);
  nand U26985(n25636,n25622,G59426);
  not U26986(n25622,n24659);
  nand U26987(n25615,n21896,n25554);
  nand U26988(n25554,n25638,n25639);
  nand U26989(n25639,n25633,n25631);
  nand U26990(n25631,n25640,n25641);
  not U26991(n25633,n25549);
  nand U26992(n25549,n25642,n25643);
  or U26993(n25638,n25641,n25632);
  nand U26994(n25632,n25644,n25645);
  nand U26995(n25641,n23169,n24659,n25623);
  nand U26996(n23169,n25646,n25647);
  nand U26997(G8497,n25648,n25649,n25650,n25651);
  nor U26998(n25651,n25652,n25653,n25654);
  nor U26999(n25654,n25655,n21845);
  nor U27000(n25653,n25656,n25657);
  nor U27001(n25652,n23145,n25658);
  nand U27002(n25650,n25659,n25660);
  nand U27003(n25649,n25661,n25662);
  nand U27004(n25648,n25663,n25664);
  nand U27005(G8496,n25665,n25666,n25667,n25668);
  nor U27006(n25668,n25669,n25670,n25671);
  nor U27007(n25671,n25655,n21837);
  nor U27008(n25670,n25656,n25672);
  nor U27009(n25669,n23049,n25658);
  nand U27010(n25667,n25659,n25673);
  nand U27011(n25666,n25674,n25662);
  nand U27012(n25665,n25663,n25675);
  nand U27013(G8495,n25676,n25677,n25678,n25679);
  nor U27014(n25679,n25680,n25681,n25682);
  nor U27015(n25682,n25655,n21829);
  nor U27016(n25681,n25656,n25683);
  nor U27017(n25680,n23587,n25658);
  nand U27018(n25678,n25659,n25684);
  nand U27019(n25677,n25685,n25662);
  nand U27020(n25676,n25663,n25686);
  nand U27021(G8494,n25687,n25688,n25689,n25690);
  nor U27022(n25690,n25691,n25692,n25693);
  nor U27023(n25693,n25655,n21821);
  nor U27024(n25692,n25656,n25694);
  nor U27025(n25691,n23502,n25658);
  nand U27026(n25689,n25659,n25695);
  nand U27027(n25688,n25696,n25662);
  nand U27028(n25687,n25663,n25697);
  nand U27029(G8493,n25698,n25699,n25700,n25701);
  nor U27030(n25701,n25702,n25703,n25704);
  nor U27031(n25704,n25655,n21812);
  nor U27032(n25703,n25656,n25705);
  nor U27033(n25702,n23418,n25658);
  nand U27034(n25700,n25659,n25706);
  nand U27035(n25699,n25707,n25662);
  nand U27036(n25698,n25663,n25708);
  nand U27037(G8492,n25709,n25710,n25711,n25712);
  nor U27038(n25712,n25713,n25714,n25715);
  nor U27039(n25715,n25655,n21803);
  nor U27040(n25714,n25656,n25716);
  nor U27041(n25713,n23337,n25658);
  nand U27042(n25711,n25659,n25717);
  nand U27043(n25710,n25718,n25662);
  nand U27044(n25709,n25663,n25719);
  nand U27045(G8491,n25720,n25721,n25722,n25723);
  nor U27046(n25723,n25724,n25725,n25726);
  nor U27047(n25726,n25655,n21794);
  nor U27048(n25725,n25656,n25727);
  nor U27049(n25724,n23257,n25658);
  nand U27050(n25722,n25659,n25728);
  nand U27051(n25721,n25729,n25662);
  nand U27052(n25720,n25663,n25730);
  nand U27053(G8490,n25731,n25732,n25733,n25734);
  nor U27054(n25734,n25735,n25736,n25737);
  nor U27055(n25737,n25655,n21784);
  and U27056(n25655,n25738,n25739);
  nand U27057(n25739,n25623,n25740,n23183,n24664);
  nand U27058(n25740,n25741,n25742);
  nand U27059(n25738,n25663,n25743);
  nor U27060(n25736,n25656,n25744);
  and U27061(n25656,n25745,n25746);
  or U27062(n25746,n25742,n22383);
  nand U27063(n25745,n25747,G59426);
  nor U27064(n25735,n22563,n25658);
  nand U27065(n25658,n25748,n25749);
  nand U27066(n25749,n25750,n25629,n25751);
  nand U27067(n25751,n25743,n25742);
  nand U27068(n25750,n25752,n24664);
  nand U27069(n25752,n25753,n21044);
  nand U27070(n25753,n25742,n23183);
  nand U27071(n25742,n25754,n25645);
  nand U27072(n25748,n25663,n25634);
  nand U27073(n25733,n25659,n25755);
  and U27074(n25659,n25623,n25747);
  not U27075(n25747,n24664);
  nand U27076(n25732,n25756,n25662);
  not U27077(n25662,n23183);
  nand U27078(n23183,n25757,n25646);
  nand U27079(n25731,n25663,n25758);
  not U27080(n25663,n25741);
  nand U27081(n25741,n25759,n25643);
  nand U27082(G8489,n25760,n25761,n25762,n25763);
  nor U27083(n25763,n25764,n25765,n25766);
  nor U27084(n25766,n21848,n25767);
  nor U27085(n25765,n25548,n25768);
  nor U27086(n25764,n23184,n25550);
  nand U27087(n25762,n25769,G59540);
  nand U27088(n25761,n25552,n25770);
  nand U27089(n25760,n21932,n25771);
  nand U27090(G8488,n25772,n25773,n25774,n25775);
  nor U27091(n25775,n25776,n25777,n25778);
  nor U27092(n25778,n21838,n25767);
  nor U27093(n25777,n25562,n25768);
  nor U27094(n25776,n23184,n25563);
  nand U27095(n25774,n25769,G59539);
  nand U27096(n25773,n25564,n25770);
  nand U27097(n25772,n21927,n25771);
  nand U27098(G8487,n25779,n25780,n25781,n25782);
  nor U27099(n25782,n25783,n25784,n25785);
  nor U27100(n25785,n21830,n25767);
  nor U27101(n25784,n25572,n25768);
  nor U27102(n25783,n23184,n25573);
  nand U27103(n25781,n25769,G59538);
  nand U27104(n25780,n25574,n25770);
  nand U27105(n25779,n21922,n25771);
  nand U27106(G8486,n25786,n25787,n25788,n25789);
  nor U27107(n25789,n25790,n25791,n25792);
  nor U27108(n25792,n21822,n25767);
  nor U27109(n25791,n25582,n25768);
  nor U27110(n25790,n23184,n25583);
  nand U27111(n25788,n25769,G59537);
  nand U27112(n25787,n25584,n25770);
  nand U27113(n25786,n21917,n25771);
  nand U27114(G8485,n25793,n25794,n25795,n25796);
  nor U27115(n25796,n25797,n25798,n25799);
  nor U27116(n25799,n21813,n25767);
  nor U27117(n25798,n25592,n25768);
  nor U27118(n25797,n23184,n25593);
  nand U27119(n25795,n25769,G59536);
  nand U27120(n25794,n25594,n25770);
  nand U27121(n25793,n21912,n25771);
  nand U27122(G8484,n25800,n25801,n25802,n25803);
  nor U27123(n25803,n25804,n25805,n25806);
  nor U27124(n25806,n21804,n25767);
  nor U27125(n25805,n25602,n25768);
  nor U27126(n25804,n23184,n25603);
  nand U27127(n25802,n25769,G59535);
  nand U27128(n25801,n25604,n25770);
  nand U27129(n25800,n21907,n25771);
  nand U27130(G8483,n25807,n25808,n25809,n25810);
  nor U27131(n25810,n25811,n25812,n25813);
  nor U27132(n25813,n21795,n25767);
  nor U27133(n25812,n25612,n25768);
  nor U27134(n25811,n23184,n25613);
  nand U27135(n25809,n25769,G59534);
  nand U27136(n25808,n25614,n25770);
  nand U27137(n25807,n21901,n25771);
  nand U27138(G8482,n25814,n25815,n25816,n25817);
  nor U27139(n25817,n25818,n25819,n25820);
  nor U27140(n25820,n21785,n25767);
  nand U27141(n25767,n25821,n23184,n25623);
  nor U27142(n25819,n25624,n25768);
  nor U27143(n25818,n23184,n25625);
  nand U27144(n25816,n25769,G59533);
  and U27145(n25769,n25822,n25823);
  nand U27146(n25823,n25824,n25629,n25825);
  nand U27147(n25825,G59426,n24640);
  nand U27148(n25824,n25826,n25827);
  nand U27149(n25822,n25828,n25634);
  nand U27150(n25815,n25635,n25770);
  nand U27151(n25770,n25829,n25830);
  or U27152(n25830,n25827,n22383);
  nand U27153(n25829,n25821,G59426);
  not U27154(n25821,n24640);
  nand U27155(n25814,n21896,n25771);
  nand U27156(n25771,n25831,n25832);
  nand U27157(n25832,n25828,n25826);
  nand U27158(n25826,n25640,n25833);
  not U27159(n25828,n25768);
  nand U27160(n25768,n25834,n25643);
  or U27161(n25831,n25833,n25827);
  nand U27162(n25827,n25835,n25645);
  nand U27163(n25833,n23184,n24640,n25623);
  nand U27164(n23184,n25836,n25647);
  nand U27165(G8481,n25837,n25838,n25839,n25840);
  nor U27166(n25840,n25841,n25842,n25843);
  nor U27167(n25843,n25548,n25844);
  nor U27168(n25842,n23177,n25550);
  nor U27169(n25841,n21848,n25845);
  nand U27170(n25839,n25846,G59532);
  nand U27171(n25838,n25552,n25847);
  nand U27172(n25837,n21932,n25848);
  nand U27173(G8480,n25849,n25850,n25851,n25852);
  nor U27174(n25852,n25853,n25854,n25855);
  nor U27175(n25855,n25562,n25844);
  nor U27176(n25854,n23177,n25563);
  nor U27177(n25853,n21838,n25845);
  nand U27178(n25851,n25846,G59531);
  nand U27179(n25850,n25564,n25847);
  nand U27180(n25849,n21927,n25848);
  nand U27181(G8479,n25856,n25857,n25858,n25859);
  nor U27182(n25859,n25860,n25861,n25862);
  nor U27183(n25862,n25572,n25844);
  nor U27184(n25861,n23177,n25573);
  nor U27185(n25860,n21830,n25845);
  nand U27186(n25858,n25846,G59530);
  nand U27187(n25857,n25574,n25847);
  nand U27188(n25856,n21922,n25848);
  nand U27189(G8478,n25863,n25864,n25865,n25866);
  nor U27190(n25866,n25867,n25868,n25869);
  nor U27191(n25869,n25582,n25844);
  nor U27192(n25868,n23177,n25583);
  nor U27193(n25867,n21822,n25845);
  nand U27194(n25865,n25846,G59529);
  nand U27195(n25864,n25584,n25847);
  nand U27196(n25863,n21917,n25848);
  nand U27197(G8477,n25870,n25871,n25872,n25873);
  nor U27198(n25873,n25874,n25875,n25876);
  nor U27199(n25876,n25592,n25844);
  nor U27200(n25875,n23177,n25593);
  nor U27201(n25874,n21813,n25845);
  nand U27202(n25872,n25846,G59528);
  nand U27203(n25871,n25594,n25847);
  nand U27204(n25870,n21912,n25848);
  nand U27205(G8476,n25877,n25878,n25879,n25880);
  nor U27206(n25880,n25881,n25882,n25883);
  nor U27207(n25883,n25602,n25844);
  nor U27208(n25882,n23177,n25603);
  nor U27209(n25881,n21804,n25845);
  nand U27210(n25879,n25846,G59527);
  nand U27211(n25878,n25604,n25847);
  nand U27212(n25877,n21907,n25848);
  nand U27213(G8475,n25884,n25885,n25886,n25887);
  nor U27214(n25887,n25888,n25889,n25890);
  nor U27215(n25890,n25612,n25844);
  nor U27216(n25889,n23177,n25613);
  nor U27217(n25888,n21795,n25845);
  nand U27218(n25886,n25846,G59526);
  nand U27219(n25885,n25614,n25847);
  nand U27220(n25884,n21901,n25848);
  nand U27221(G8474,n25891,n25892,n25893,n25894);
  nor U27222(n25894,n25895,n25896,n25897);
  nor U27223(n25897,n25624,n25844);
  nor U27224(n25896,n23177,n25625);
  nor U27225(n25895,n21785,n25845);
  nand U27226(n25845,n25623,n25898);
  nand U27227(n25893,n25846,G59525);
  and U27228(n25846,n25899,n25900);
  nand U27229(n25900,n25901,n25629,n25902);
  nand U27230(n25902,G59426,n24641);
  nand U27231(n25901,n25903,n25904);
  nand U27232(n25899,n25905,n25634);
  nand U27233(n25892,n25635,n25847);
  nand U27234(n25847,n25906,n25907);
  nand U27235(n25907,n25908,n22435);
  nand U27236(n25906,n25898,G59426);
  not U27237(n25898,n24641);
  nand U27238(n25891,n21896,n25848);
  nand U27239(n25848,n25909,n25910);
  nand U27240(n25910,n25623,n23177,n25908);
  not U27241(n25908,n25904);
  nand U27242(n25904,n25911,n25645);
  nor U27243(n25645,n25912,n25913);
  nand U27244(n25909,n25905,n25903);
  nand U27245(n25903,n25640,n25914);
  nand U27246(n25914,n23177,n24641,n25623);
  nand U27247(n23177,n25836,n25757);
  not U27248(n25905,n25844);
  nand U27249(n25844,n25643,n25915);
  nor U27250(n25643,G59564,G59563);
  nand U27251(G8473,n25916,n25917,n25918,n25919);
  nor U27252(n25919,n25920,n25921,n25922);
  nor U27253(n25922,n21848,n25923);
  nor U27254(n25921,n25548,n25924);
  nor U27255(n25920,n23176,n25550);
  nand U27256(n25918,n25925,G59524);
  nand U27257(n25917,n25552,n25926);
  nand U27258(n25916,n21932,n25927);
  nand U27259(G8472,n25928,n25929,n25930,n25931);
  nor U27260(n25931,n25932,n25933,n25934);
  nor U27261(n25934,n21838,n25923);
  nor U27262(n25933,n25562,n25924);
  nor U27263(n25932,n23176,n25563);
  nand U27264(n25930,n25925,G59523);
  nand U27265(n25929,n25564,n25926);
  nand U27266(n25928,n21927,n25927);
  nand U27267(G8471,n25935,n25936,n25937,n25938);
  nor U27268(n25938,n25939,n25940,n25941);
  nor U27269(n25941,n21830,n25923);
  nor U27270(n25940,n25572,n25924);
  nor U27271(n25939,n23176,n25573);
  nand U27272(n25937,n25925,G59522);
  nand U27273(n25936,n25574,n25926);
  nand U27274(n25935,n21922,n25927);
  nand U27275(G8470,n25942,n25943,n25944,n25945);
  nor U27276(n25945,n25946,n25947,n25948);
  nor U27277(n25948,n21822,n25923);
  nor U27278(n25947,n25582,n25924);
  nor U27279(n25946,n23176,n25583);
  nand U27280(n25944,n25925,G59521);
  nand U27281(n25943,n25584,n25926);
  nand U27282(n25942,n21917,n25927);
  nand U27283(G8469,n25949,n25950,n25951,n25952);
  nor U27284(n25952,n25953,n25954,n25955);
  nor U27285(n25955,n21813,n25923);
  nor U27286(n25954,n25592,n25924);
  nor U27287(n25953,n23176,n25593);
  nand U27288(n25951,n25925,G59520);
  nand U27289(n25950,n25594,n25926);
  nand U27290(n25949,n21912,n25927);
  nand U27291(G8468,n25956,n25957,n25958,n25959);
  nor U27292(n25959,n25960,n25961,n25962);
  nor U27293(n25962,n21804,n25923);
  nor U27294(n25961,n25602,n25924);
  nor U27295(n25960,n23176,n25603);
  nand U27296(n25958,n25925,G59519);
  nand U27297(n25957,n25604,n25926);
  nand U27298(n25956,n21907,n25927);
  nand U27299(G8467,n25963,n25964,n25965,n25966);
  nor U27300(n25966,n25967,n25968,n25969);
  nor U27301(n25969,n21795,n25923);
  nor U27302(n25968,n25612,n25924);
  nor U27303(n25967,n23176,n25613);
  nand U27304(n25965,n25925,G59518);
  nand U27305(n25964,n25614,n25926);
  nand U27306(n25963,n21901,n25927);
  nand U27307(G8466,n25970,n25971,n25972,n25973);
  nor U27308(n25973,n25974,n25975,n25976);
  nor U27309(n25976,n21785,n25923);
  nand U27310(n25923,n25977,n23176,n25623);
  nor U27311(n25975,n25624,n25924);
  nor U27312(n25974,n23176,n25625);
  nand U27313(n25972,n25925,G59517);
  and U27314(n25925,n25978,n25979);
  nand U27315(n25979,n25980,n25629,n25981);
  nand U27316(n25981,G59426,n24642);
  nand U27317(n25980,n25982,n25983);
  nand U27318(n25978,n25984,n25634);
  nand U27319(n25971,n25635,n25926);
  nand U27320(n25926,n25985,n25986);
  or U27321(n25986,n25983,n22383);
  nand U27322(n25985,n25977,G59426);
  not U27323(n25977,n24642);
  nand U27324(n25970,n21896,n25927);
  nand U27325(n25927,n25987,n25988);
  nand U27326(n25988,n25984,n25982);
  nand U27327(n25982,n25640,n25989);
  not U27328(n25984,n25924);
  nand U27329(n25924,n25642,n25990);
  or U27330(n25987,n25989,n25983);
  nand U27331(n25983,n25991,n25644);
  nand U27332(n25989,n23176,n24642,n25623);
  nand U27333(n23176,n25992,n25646);
  nand U27334(G8465,n25993,n25994,n25995,n25996);
  nor U27335(n25996,n25997,n25998,n25999);
  nor U27336(n25999,n25548,n26000);
  nor U27337(n25998,n23162,n25550);
  nor U27338(n25997,n21848,n26001);
  nand U27339(n25995,n26002,G59516);
  nand U27340(n25994,n25552,n26003);
  nand U27341(n25993,n21932,n26004);
  nand U27342(G8464,n26005,n26006,n26007,n26008);
  nor U27343(n26008,n26009,n26010,n26011);
  nor U27344(n26011,n25562,n26000);
  nor U27345(n26010,n23162,n25563);
  nor U27346(n26009,n21838,n26001);
  nand U27347(n26007,n26002,G59515);
  nand U27348(n26006,n25564,n26003);
  nand U27349(n26005,n21927,n26004);
  nand U27350(G8463,n26012,n26013,n26014,n26015);
  nor U27351(n26015,n26016,n26017,n26018);
  nor U27352(n26018,n25572,n26000);
  nor U27353(n26017,n23162,n25573);
  nor U27354(n26016,n21830,n26001);
  nand U27355(n26014,n26002,G59514);
  nand U27356(n26013,n25574,n26003);
  nand U27357(n26012,n21922,n26004);
  nand U27358(G8462,n26019,n26020,n26021,n26022);
  nor U27359(n26022,n26023,n26024,n26025);
  nor U27360(n26025,n25582,n26000);
  nor U27361(n26024,n23162,n25583);
  nor U27362(n26023,n21822,n26001);
  nand U27363(n26021,n26002,G59513);
  nand U27364(n26020,n25584,n26003);
  nand U27365(n26019,n21917,n26004);
  nand U27366(G8461,n26026,n26027,n26028,n26029);
  nor U27367(n26029,n26030,n26031,n26032);
  nor U27368(n26032,n25592,n26000);
  nor U27369(n26031,n23162,n25593);
  nor U27370(n26030,n21813,n26001);
  nand U27371(n26028,n26002,G59512);
  nand U27372(n26027,n25594,n26003);
  nand U27373(n26026,n21912,n26004);
  nand U27374(G8460,n26033,n26034,n26035,n26036);
  nor U27375(n26036,n26037,n26038,n26039);
  nor U27376(n26039,n25602,n26000);
  nor U27377(n26038,n23162,n25603);
  nor U27378(n26037,n21804,n26001);
  nand U27379(n26035,n26002,G59511);
  nand U27380(n26034,n25604,n26003);
  nand U27381(n26033,n21907,n26004);
  nand U27382(G8459,n26040,n26041,n26042,n26043);
  nor U27383(n26043,n26044,n26045,n26046);
  nor U27384(n26046,n25612,n26000);
  nor U27385(n26045,n23162,n25613);
  nor U27386(n26044,n21795,n26001);
  nand U27387(n26042,n26002,G59510);
  nand U27388(n26041,n25614,n26003);
  nand U27389(n26040,n21901,n26004);
  nand U27390(G8458,n26047,n26048,n26049,n26050);
  nor U27391(n26050,n26051,n26052,n26053);
  nor U27392(n26053,n25624,n26000);
  nor U27393(n26052,n23162,n25625);
  nor U27394(n26051,n21785,n26001);
  nand U27395(n26001,n25623,n26054);
  nand U27396(n26049,n26002,G59509);
  and U27397(n26002,n26055,n26056);
  nand U27398(n26056,n26057,n25629,n26058);
  nand U27399(n26058,G59426,n24665);
  nand U27400(n26057,n26059,n26060);
  nand U27401(n26055,n26061,n25634);
  nand U27402(n26048,n25635,n26003);
  nand U27403(n26003,n26062,n26063);
  nand U27404(n26063,n26064,n22435);
  nand U27405(n26062,n26054,G59426);
  not U27406(n26054,n24665);
  nand U27407(n26047,n21896,n26004);
  nand U27408(n26004,n26065,n26066);
  nand U27409(n26066,n25623,n23162,n26064);
  not U27410(n26064,n26060);
  nand U27411(n26060,n25991,n25754);
  nand U27412(n26065,n26061,n26059);
  nand U27413(n26059,n25640,n26067);
  nand U27414(n26067,n23162,n24665,n25623);
  nand U27415(n23162,n26068,n25646);
  nor U27416(n25646,n26069,n26070);
  not U27417(n26061,n26000);
  nand U27418(n26000,n25759,n25990);
  nand U27419(G8457,n26071,n26072,n26073,n26074);
  nor U27420(n26074,n26075,n26076,n26077);
  nor U27421(n26077,n21848,n26078);
  nor U27422(n26076,n25548,n26079);
  nor U27423(n26075,n23175,n25550);
  nand U27424(n26073,n26080,G59508);
  nand U27425(n26072,n25552,n26081);
  nand U27426(n26071,n21932,n26082);
  nand U27427(G8456,n26083,n26084,n26085,n26086);
  nor U27428(n26086,n26087,n26088,n26089);
  nor U27429(n26089,n21838,n26078);
  nor U27430(n26088,n25562,n26079);
  nor U27431(n26087,n23175,n25563);
  nand U27432(n26085,n26080,G59507);
  nand U27433(n26084,n25564,n26081);
  nand U27434(n26083,n21927,n26082);
  nand U27435(G8455,n26090,n26091,n26092,n26093);
  nor U27436(n26093,n26094,n26095,n26096);
  nor U27437(n26096,n21830,n26078);
  nor U27438(n26095,n25572,n26079);
  nor U27439(n26094,n23175,n25573);
  nand U27440(n26092,n26080,G59506);
  nand U27441(n26091,n25574,n26081);
  nand U27442(n26090,n21922,n26082);
  nand U27443(G8454,n26097,n26098,n26099,n26100);
  nor U27444(n26100,n26101,n26102,n26103);
  nor U27445(n26103,n21822,n26078);
  nor U27446(n26102,n25582,n26079);
  nor U27447(n26101,n23175,n25583);
  nand U27448(n26099,n26080,G59505);
  nand U27449(n26098,n25584,n26081);
  nand U27450(n26097,n21917,n26082);
  nand U27451(G8453,n26104,n26105,n26106,n26107);
  nor U27452(n26107,n26108,n26109,n26110);
  nor U27453(n26110,n21813,n26078);
  nor U27454(n26109,n25592,n26079);
  nor U27455(n26108,n23175,n25593);
  nand U27456(n26106,n26080,G59504);
  nand U27457(n26105,n25594,n26081);
  nand U27458(n26104,n21912,n26082);
  nand U27459(G8452,n26111,n26112,n26113,n26114);
  nor U27460(n26114,n26115,n26116,n26117);
  nor U27461(n26117,n21804,n26078);
  nor U27462(n26116,n25602,n26079);
  nor U27463(n26115,n23175,n25603);
  nand U27464(n26113,n26080,G59503);
  nand U27465(n26112,n25604,n26081);
  nand U27466(n26111,n21907,n26082);
  nand U27467(G8451,n26118,n26119,n26120,n26121);
  nor U27468(n26121,n26122,n26123,n26124);
  nor U27469(n26124,n21795,n26078);
  nor U27470(n26123,n25612,n26079);
  nor U27471(n26122,n23175,n25613);
  nand U27472(n26120,n26080,G59502);
  nand U27473(n26119,n25614,n26081);
  nand U27474(n26118,n21901,n26082);
  nand U27475(G8450,n26125,n26126,n26127,n26128);
  nor U27476(n26128,n26129,n26130,n26131);
  nor U27477(n26131,n21785,n26078);
  nand U27478(n26078,n26132,n23175,n25623);
  nor U27479(n26130,n25624,n26079);
  nor U27480(n26129,n23175,n25625);
  nand U27481(n26127,n26080,G59501);
  and U27482(n26080,n26133,n26134);
  nand U27483(n26134,n26135,n25629,n26136);
  nand U27484(n26136,G59426,n24643);
  nand U27485(n26135,n26137,n26138);
  nand U27486(n26133,n26139,n25634);
  nand U27487(n26126,n25635,n26081);
  nand U27488(n26081,n26140,n26141);
  or U27489(n26141,n26138,n22383);
  nand U27490(n26140,n26132,G59426);
  not U27491(n26132,n24643);
  nand U27492(n26125,n21896,n26082);
  nand U27493(n26082,n26142,n26143);
  nand U27494(n26143,n26139,n26137);
  nand U27495(n26137,n25640,n26144);
  not U27496(n26139,n26079);
  nand U27497(n26079,n25834,n25990);
  or U27498(n26142,n26144,n26138);
  nand U27499(n26138,n25991,n25835);
  nand U27500(n26144,n23175,n24643,n25623);
  nand U27501(n23175,n25992,n25836);
  nand U27502(G8449,n26145,n26146,n26147,n26148);
  nor U27503(n26148,n26149,n26150,n26151);
  nor U27504(n26151,n21848,n26152);
  nor U27505(n26150,n23185,n25550);
  nor U27506(n26149,n25548,n26153);
  nand U27507(n26147,n26154,G59500);
  nand U27508(n26146,n25552,n26155);
  nand U27509(n26145,n21932,n26156);
  nand U27510(G8448,n26157,n26158,n26159,n26160);
  nor U27511(n26160,n26161,n26162,n26163);
  nor U27512(n26163,n21838,n26152);
  nor U27513(n26162,n23185,n25563);
  nor U27514(n26161,n25562,n26153);
  nand U27515(n26159,n26154,G59499);
  nand U27516(n26158,n25564,n26155);
  nand U27517(n26157,n21927,n26156);
  nand U27518(G8447,n26164,n26165,n26166,n26167);
  nor U27519(n26167,n26168,n26169,n26170);
  nor U27520(n26170,n21830,n26152);
  nor U27521(n26169,n23185,n25573);
  nor U27522(n26168,n25572,n26153);
  nand U27523(n26166,n26154,G59498);
  nand U27524(n26165,n25574,n26155);
  nand U27525(n26164,n21922,n26156);
  nand U27526(G8446,n26171,n26172,n26173,n26174);
  nor U27527(n26174,n26175,n26176,n26177);
  nor U27528(n26177,n21822,n26152);
  nor U27529(n26176,n23185,n25583);
  nor U27530(n26175,n25582,n26153);
  nand U27531(n26173,n26154,G59497);
  nand U27532(n26172,n25584,n26155);
  nand U27533(n26171,n21917,n26156);
  nand U27534(G8445,n26178,n26179,n26180,n26181);
  nor U27535(n26181,n26182,n26183,n26184);
  nor U27536(n26184,n21813,n26152);
  nor U27537(n26183,n23185,n25593);
  nor U27538(n26182,n25592,n26153);
  nand U27539(n26180,n26154,G59496);
  nand U27540(n26179,n25594,n26155);
  nand U27541(n26178,n21912,n26156);
  nand U27542(G8444,n26185,n26186,n26187,n26188);
  nor U27543(n26188,n26189,n26190,n26191);
  nor U27544(n26191,n21804,n26152);
  nor U27545(n26190,n23185,n25603);
  nor U27546(n26189,n25602,n26153);
  nand U27547(n26187,n26154,G59495);
  nand U27548(n26186,n25604,n26155);
  nand U27549(n26185,n21907,n26156);
  nand U27550(G8443,n26192,n26193,n26194,n26195);
  nor U27551(n26195,n26196,n26197,n26198);
  nor U27552(n26198,n21795,n26152);
  nor U27553(n26197,n23185,n25613);
  nor U27554(n26196,n25612,n26153);
  nand U27555(n26194,n26154,G59494);
  nand U27556(n26193,n25614,n26155);
  nand U27557(n26192,n21901,n26156);
  nand U27558(G8442,n26199,n26200,n26201,n26202);
  nor U27559(n26202,n26203,n26204,n26205);
  nor U27560(n26205,n21785,n26152);
  nand U27561(n26152,n25623,n26206);
  nor U27562(n26204,n23185,n25625);
  nor U27563(n26203,n25624,n26153);
  nand U27564(n26201,n26154,G59493);
  and U27565(n26154,n26207,n26208);
  nand U27566(n26208,n26209,n25629,n26210);
  nand U27567(n26210,G59426,n24648);
  nand U27568(n26209,n26211,n26212);
  nand U27569(n26207,n26213,n25634);
  nand U27570(n26200,n25635,n26155);
  nand U27571(n26155,n26214,n26215);
  nand U27572(n26215,n26216,n22435);
  nand U27573(n26214,n26206,G59426);
  not U27574(n26206,n24648);
  nand U27575(n26199,n21896,n26156);
  nand U27576(n26156,n26217,n26218);
  nand U27577(n26218,n25623,n23185,n26216);
  not U27578(n26216,n26212);
  nand U27579(n26212,n25991,n25911);
  nor U27580(n25991,n25912,n26219);
  nand U27581(n26217,n26213,n26211);
  nand U27582(n26211,n25640,n26220);
  nand U27583(n26220,n23185,n24648,n25623);
  nand U27584(n23185,n26068,n25836);
  nor U27585(n25836,n26070,n26221);
  nand U27586(G8441,n26222,n26223,n26224,n26225);
  nor U27587(n26225,n26226,n26227,n26228);
  nor U27588(n26228,n21848,n26229);
  nor U27589(n26227,n25548,n26230);
  nor U27590(n26226,n23168,n25550);
  nand U27591(n26224,n26231,G59492);
  nand U27592(n26223,n25552,n26232);
  nand U27593(n26222,n21932,n26233);
  nand U27594(G8440,n26234,n26235,n26236,n26237);
  nor U27595(n26237,n26238,n26239,n26240);
  nor U27596(n26240,n21838,n26229);
  nor U27597(n26239,n25562,n26230);
  nor U27598(n26238,n23168,n25563);
  nand U27599(n26236,n26231,G59491);
  nand U27600(n26235,n25564,n26232);
  nand U27601(n26234,n21927,n26233);
  nand U27602(G8439,n26241,n26242,n26243,n26244);
  nor U27603(n26244,n26245,n26246,n26247);
  nor U27604(n26247,n21830,n26229);
  nor U27605(n26246,n25572,n26230);
  nor U27606(n26245,n23168,n25573);
  nand U27607(n26243,n26231,G59490);
  nand U27608(n26242,n25574,n26232);
  nand U27609(n26241,n21922,n26233);
  nand U27610(G8438,n26248,n26249,n26250,n26251);
  nor U27611(n26251,n26252,n26253,n26254);
  nor U27612(n26254,n21822,n26229);
  nor U27613(n26253,n25582,n26230);
  nor U27614(n26252,n23168,n25583);
  nand U27615(n26250,n26231,G59489);
  nand U27616(n26249,n25584,n26232);
  nand U27617(n26248,n21917,n26233);
  nand U27618(G8437,n26255,n26256,n26257,n26258);
  nor U27619(n26258,n26259,n26260,n26261);
  nor U27620(n26261,n21813,n26229);
  nor U27621(n26260,n25592,n26230);
  nor U27622(n26259,n23168,n25593);
  nand U27623(n26257,n26231,G59488);
  nand U27624(n26256,n25594,n26232);
  nand U27625(n26255,n21912,n26233);
  nand U27626(G8436,n26262,n26263,n26264,n26265);
  nor U27627(n26265,n26266,n26267,n26268);
  nor U27628(n26268,n21804,n26229);
  nor U27629(n26267,n25602,n26230);
  nor U27630(n26266,n23168,n25603);
  nand U27631(n26264,n26231,G59487);
  nand U27632(n26263,n25604,n26232);
  nand U27633(n26262,n21907,n26233);
  nand U27634(G8435,n26269,n26270,n26271,n26272);
  nor U27635(n26272,n26273,n26274,n26275);
  nor U27636(n26275,n21795,n26229);
  nor U27637(n26274,n25612,n26230);
  nor U27638(n26273,n23168,n25613);
  nand U27639(n26271,n26231,G59486);
  nand U27640(n26270,n25614,n26232);
  nand U27641(n26269,n21901,n26233);
  nand U27642(G8434,n26276,n26277,n26278,n26279);
  nor U27643(n26279,n26280,n26281,n26282);
  nor U27644(n26282,n21785,n26229);
  nand U27645(n26229,n26283,n23168,n25623);
  nor U27646(n26281,n25624,n26230);
  nor U27647(n26280,n23168,n25625);
  nand U27648(n26278,n26231,G59485);
  and U27649(n26231,n26284,n26285);
  nand U27650(n26285,n26286,n25629,n26287);
  nand U27651(n26287,G59426,n24649);
  nand U27652(n26286,n26288,n26289);
  nand U27653(n26284,n26290,n25634);
  nand U27654(n26277,n25635,n26232);
  nand U27655(n26232,n26291,n26292);
  or U27656(n26292,n26289,n22383);
  nand U27657(n26291,n26283,G59426);
  not U27658(n26283,n24649);
  nand U27659(n26276,n21896,n26233);
  nand U27660(n26233,n26293,n26294);
  nand U27661(n26294,n26290,n26288);
  nand U27662(n26288,n25640,n26295);
  not U27663(n26290,n26230);
  nand U27664(n26230,n26296,n25642);
  or U27665(n26293,n26295,n26289);
  nand U27666(n26289,n26297,n25644);
  nand U27667(n26295,n23168,n24649,n25623);
  nand U27668(n23168,n26298,n25647);
  nand U27669(G8433,n26299,n26300,n26301,n26302);
  nor U27670(n26302,n26303,n26304,n26305);
  nor U27671(n26305,n26306,n21845);
  nor U27672(n26304,n26307,n25657);
  nor U27673(n26303,n23124,n26308);
  nand U27674(n26301,n26309,n25660);
  nand U27675(n26300,n25661,n26310);
  nand U27676(n26299,n26311,n25664);
  nand U27677(G8432,n26312,n26313,n26314,n26315);
  nor U27678(n26315,n26316,n26317,n26318);
  nor U27679(n26318,n26306,n21837);
  nor U27680(n26317,n26307,n25672);
  nor U27681(n26316,n23033,n26308);
  nand U27682(n26314,n26309,n25673);
  nand U27683(n26313,n25674,n26310);
  nand U27684(n26312,n26311,n25675);
  nand U27685(G8431,n26319,n26320,n26321,n26322);
  nor U27686(n26322,n26323,n26324,n26325);
  nor U27687(n26325,n26306,n21829);
  nor U27688(n26324,n26307,n25683);
  nor U27689(n26323,n22963,n26308);
  nand U27690(n26321,n26309,n25684);
  nand U27691(n26320,n25685,n26310);
  nand U27692(n26319,n26311,n25686);
  nand U27693(G8430,n26326,n26327,n26328,n26329);
  nor U27694(n26329,n26330,n26331,n26332);
  nor U27695(n26332,n26306,n21821);
  nor U27696(n26331,n26307,n25694);
  nor U27697(n26330,n22884,n26308);
  nand U27698(n26328,n26309,n25695);
  nand U27699(n26327,n25696,n26310);
  nand U27700(n26326,n26311,n25697);
  nand U27701(G8429,n26333,n26334,n26335,n26336);
  nor U27702(n26336,n26337,n26338,n26339);
  nor U27703(n26339,n26306,n21812);
  nor U27704(n26338,n26307,n25705);
  nor U27705(n26337,n22810,n26308);
  nand U27706(n26335,n26309,n25706);
  nand U27707(n26334,n25707,n26310);
  nand U27708(n26333,n26311,n25708);
  nand U27709(G8428,n26340,n26341,n26342,n26343);
  nor U27710(n26343,n26344,n26345,n26346);
  nor U27711(n26346,n26306,n21803);
  nor U27712(n26345,n26307,n25716);
  nor U27713(n26344,n22729,n26308);
  nand U27714(n26342,n26309,n25717);
  nand U27715(n26341,n25718,n26310);
  nand U27716(n26340,n26311,n25719);
  nand U27717(G8427,n26347,n26348,n26349,n26350);
  nor U27718(n26350,n26351,n26352,n26353);
  nor U27719(n26353,n26306,n21794);
  nor U27720(n26352,n26307,n25727);
  nor U27721(n26351,n22653,n26308);
  nand U27722(n26349,n26309,n25728);
  nand U27723(n26348,n25729,n26310);
  nand U27724(n26347,n26311,n25730);
  nand U27725(G8426,n26354,n26355,n26356,n26357);
  nor U27726(n26357,n26358,n26359,n26360);
  nor U27727(n26360,n26306,n21784);
  and U27728(n26306,n26361,n26362);
  nand U27729(n26362,n25623,n26363,n23161,n24666);
  nand U27730(n26363,n26364,n26365);
  nand U27731(n26361,n26311,n25743);
  nor U27732(n26359,n26307,n25744);
  and U27733(n26307,n26366,n26367);
  or U27734(n26367,n26365,n22383);
  nand U27735(n26366,n26368,G59426);
  nor U27736(n26358,n22539,n26308);
  nand U27737(n26308,n26369,n26370);
  nand U27738(n26370,n26371,n25629,n26372);
  nand U27739(n26372,n25743,n26365);
  nand U27740(n26371,n26373,n24666);
  nand U27741(n26373,n26374,n21044);
  nand U27742(n26374,n26365,n23161);
  nand U27743(n26365,n26297,n25754);
  nand U27744(n26369,n26311,n25634);
  nand U27745(n26356,n26309,n25755);
  and U27746(n26309,n25623,n26368);
  not U27747(n26368,n24666);
  nand U27748(n26355,n25756,n26310);
  not U27749(n26310,n23161);
  nand U27750(n23161,n26298,n25757);
  nand U27751(n26354,n26311,n25758);
  not U27752(n26311,n26364);
  nand U27753(n26364,n26296,n25759);
  nand U27754(G8425,n26375,n26376,n26377,n26378);
  nor U27755(n26378,n26379,n26380,n26381);
  nor U27756(n26381,n21848,n26382);
  nor U27757(n26380,n25548,n26383);
  nor U27758(n26379,n23167,n25550);
  nand U27759(n26377,n26384,G59476);
  nand U27760(n26376,n25552,n26385);
  nand U27761(n26375,n21932,n26386);
  nand U27762(G8424,n26387,n26388,n26389,n26390);
  nor U27763(n26390,n26391,n26392,n26393);
  nor U27764(n26393,n21838,n26382);
  nor U27765(n26392,n25562,n26383);
  nor U27766(n26391,n23167,n25563);
  nand U27767(n26389,n26384,G59475);
  nand U27768(n26388,n25564,n26385);
  nand U27769(n26387,n21927,n26386);
  nand U27770(G8423,n26394,n26395,n26396,n26397);
  nor U27771(n26397,n26398,n26399,n26400);
  nor U27772(n26400,n21830,n26382);
  nor U27773(n26399,n25572,n26383);
  nor U27774(n26398,n23167,n25573);
  nand U27775(n26396,n26384,G59474);
  nand U27776(n26395,n25574,n26385);
  nand U27777(n26394,n21922,n26386);
  nand U27778(G8422,n26401,n26402,n26403,n26404);
  nor U27779(n26404,n26405,n26406,n26407);
  nor U27780(n26407,n21822,n26382);
  nor U27781(n26406,n25582,n26383);
  nor U27782(n26405,n23167,n25583);
  nand U27783(n26403,n26384,G59473);
  nand U27784(n26402,n25584,n26385);
  nand U27785(n26401,n21917,n26386);
  nand U27786(G8421,n26408,n26409,n26410,n26411);
  nor U27787(n26411,n26412,n26413,n26414);
  nor U27788(n26414,n21813,n26382);
  nor U27789(n26413,n25592,n26383);
  nor U27790(n26412,n23167,n25593);
  nand U27791(n26410,n26384,G59472);
  nand U27792(n26409,n25594,n26385);
  nand U27793(n26408,n21912,n26386);
  nand U27794(G8420,n26415,n26416,n26417,n26418);
  nor U27795(n26418,n26419,n26420,n26421);
  nor U27796(n26421,n21804,n26382);
  nor U27797(n26420,n25602,n26383);
  nor U27798(n26419,n23167,n25603);
  nand U27799(n26417,n26384,G59471);
  nand U27800(n26416,n25604,n26385);
  nand U27801(n26415,n21907,n26386);
  nand U27802(G8419,n26422,n26423,n26424,n26425);
  nor U27803(n26425,n26426,n26427,n26428);
  nor U27804(n26428,n21795,n26382);
  nor U27805(n26427,n25612,n26383);
  nor U27806(n26426,n23167,n25613);
  nand U27807(n26424,n26384,G59470);
  nand U27808(n26423,n25614,n26385);
  nand U27809(n26422,n21901,n26386);
  nand U27810(G8418,n26429,n26430,n26431,n26432);
  nor U27811(n26432,n26433,n26434,n26435);
  nor U27812(n26435,n21785,n26382);
  nand U27813(n26382,n26436,n23167,n25623);
  nor U27814(n26434,n25624,n26383);
  nor U27815(n26433,n23167,n25625);
  nand U27816(n26431,n26384,G59469);
  and U27817(n26384,n26437,n26438);
  nand U27818(n26438,n26439,n25629,n26440);
  nand U27819(n26440,G59426,n24650);
  nand U27820(n26439,n26441,n26442);
  nand U27821(n26437,n26443,n25634);
  nand U27822(n26430,n25635,n26385);
  nand U27823(n26385,n26444,n26445);
  or U27824(n26445,n26442,n22383);
  nand U27825(n26444,n26436,G59426);
  not U27826(n26436,n24650);
  nand U27827(n26429,n21896,n26386);
  nand U27828(n26386,n26446,n26447);
  nand U27829(n26447,n26443,n26441);
  nand U27830(n26441,n25640,n26448);
  not U27831(n26443,n26383);
  nand U27832(n26383,n26296,n25834);
  or U27833(n26446,n26448,n26442);
  nand U27834(n26442,n26297,n25835);
  nand U27835(n26448,n23167,n24650,n25623);
  nand U27836(n23167,n26449,n25647);
  and U27837(n25647,n26450,n26451);
  nand U27838(G8417,n26452,n26453,n26454,n26455);
  nor U27839(n26455,n26456,n26457,n26458);
  nor U27840(n26458,n25548,n26459);
  nor U27841(n26457,n23178,n25550);
  nor U27842(n26456,n21848,n26460);
  nand U27843(n26454,n26461,G59468);
  nand U27844(n26453,n25552,n26462);
  nand U27845(n26452,n21932,n26463);
  nand U27846(G8416,n26464,n26465,n26466,n26467);
  nor U27847(n26467,n26468,n26469,n26470);
  nor U27848(n26470,n25562,n26459);
  nor U27849(n26469,n23178,n25563);
  nor U27850(n26468,n21838,n26460);
  nand U27851(n26466,n26461,G59467);
  nand U27852(n26465,n25564,n26462);
  nand U27853(n26464,n21927,n26463);
  nand U27854(G8415,n26471,n26472,n26473,n26474);
  nor U27855(n26474,n26475,n26476,n26477);
  nor U27856(n26477,n25572,n26459);
  nor U27857(n26476,n23178,n25573);
  nor U27858(n26475,n21830,n26460);
  nand U27859(n26473,n26461,G59466);
  nand U27860(n26472,n25574,n26462);
  nand U27861(n26471,n21922,n26463);
  nand U27862(G8414,n26478,n26479,n26480,n26481);
  nor U27863(n26481,n26482,n26483,n26484);
  nor U27864(n26484,n25582,n26459);
  nor U27865(n26483,n23178,n25583);
  nor U27866(n26482,n21822,n26460);
  nand U27867(n26480,n26461,G59465);
  nand U27868(n26479,n25584,n26462);
  nand U27869(n26478,n21917,n26463);
  nand U27870(G8413,n26485,n26486,n26487,n26488);
  nor U27871(n26488,n26489,n26490,n26491);
  nor U27872(n26491,n25592,n26459);
  nor U27873(n26490,n23178,n25593);
  nor U27874(n26489,n21813,n26460);
  nand U27875(n26487,n26461,G59464);
  nand U27876(n26486,n25594,n26462);
  nand U27877(n26485,n21912,n26463);
  nand U27878(G8412,n26492,n26493,n26494,n26495);
  nor U27879(n26495,n26496,n26497,n26498);
  nor U27880(n26498,n25602,n26459);
  nor U27881(n26497,n23178,n25603);
  nor U27882(n26496,n21804,n26460);
  nand U27883(n26494,n26461,G59463);
  nand U27884(n26493,n25604,n26462);
  nand U27885(n26492,n21907,n26463);
  nand U27886(G8411,n26499,n26500,n26501,n26502);
  nor U27887(n26502,n26503,n26504,n26505);
  nor U27888(n26505,n25612,n26459);
  nor U27889(n26504,n23178,n25613);
  nor U27890(n26503,n21795,n26460);
  nand U27891(n26501,n26461,G59462);
  nand U27892(n26500,n25614,n26462);
  nand U27893(n26499,n21901,n26463);
  nand U27894(G8410,n26506,n26507,n26508,n26509);
  nor U27895(n26509,n26510,n26511,n26512);
  nor U27896(n26512,n25624,n26459);
  nor U27897(n26511,n23178,n25625);
  nor U27898(n26510,n21785,n26460);
  nand U27899(n26460,n25623,n26513);
  nand U27900(n26508,n26461,G59461);
  and U27901(n26461,n26514,n26515);
  nand U27902(n26515,n26516,n25629,n26517);
  nand U27903(n26517,G59426,n24651);
  nand U27904(n26516,n26518,n26519);
  nand U27905(n26514,n26520,n25634);
  nand U27906(n26507,n25635,n26462);
  nand U27907(n26462,n26521,n26522);
  nand U27908(n26522,n26523,n22435);
  nand U27909(n26521,n26513,G59426);
  not U27910(n26513,n24651);
  nand U27911(n26506,n21896,n26463);
  nand U27912(n26463,n26524,n26525);
  nand U27913(n26525,n25623,n23178,n26523);
  not U27914(n26523,n26519);
  nand U27915(n26519,n26297,n25911);
  nor U27916(n26297,n25913,n26526);
  nand U27917(n26524,n26520,n26518);
  nand U27918(n26518,n25640,n26527);
  nand U27919(n26527,n23178,n24651,n25623);
  nand U27920(n23178,n26449,n25757);
  and U27921(n25757,n26528,n26450);
  not U27922(n26520,n26459);
  nand U27923(n26459,n26296,n25915);
  nand U27924(G8409,n26529,n26530,n26531,n26532);
  nor U27925(n26532,n26533,n26534,n26535);
  nor U27926(n26535,n21848,n26536);
  nor U27927(n26534,n25548,n26537);
  nor U27928(n26533,n23186,n25550);
  nand U27929(n26531,n26538,G59460);
  nand U27930(n26530,n25552,n26539);
  nand U27931(n26529,n21932,n26540);
  nand U27932(G8408,n26541,n26542,n26543,n26544);
  nor U27933(n26544,n26545,n26546,n26547);
  nor U27934(n26547,n21838,n26536);
  nor U27935(n26546,n25562,n26537);
  nor U27936(n26545,n23186,n25563);
  nand U27937(n26543,n26538,G59459);
  nand U27938(n26542,n25564,n26539);
  nand U27939(n26541,n21927,n26540);
  nand U27940(G8407,n26548,n26549,n26550,n26551);
  nor U27941(n26551,n26552,n26553,n26554);
  nor U27942(n26554,n21830,n26536);
  nor U27943(n26553,n25572,n26537);
  nor U27944(n26552,n23186,n25573);
  nand U27945(n26550,n26538,G59458);
  nand U27946(n26549,n25574,n26539);
  nand U27947(n26548,n21922,n26540);
  nand U27948(G8406,n26555,n26556,n26557,n26558);
  nor U27949(n26558,n26559,n26560,n26561);
  nor U27950(n26561,n21822,n26536);
  nor U27951(n26560,n25582,n26537);
  nor U27952(n26559,n23186,n25583);
  nand U27953(n26557,n26538,G59457);
  nand U27954(n26556,n25584,n26539);
  nand U27955(n26555,n21917,n26540);
  nand U27956(G8405,n26562,n26563,n26564,n26565);
  nor U27957(n26565,n26566,n26567,n26568);
  nor U27958(n26568,n21813,n26536);
  nor U27959(n26567,n25592,n26537);
  nor U27960(n26566,n23186,n25593);
  nand U27961(n26564,n26538,G59456);
  nand U27962(n26563,n25594,n26539);
  nand U27963(n26562,n21912,n26540);
  nand U27964(G8404,n26569,n26570,n26571,n26572);
  nor U27965(n26572,n26573,n26574,n26575);
  nor U27966(n26575,n21804,n26536);
  nor U27967(n26574,n25602,n26537);
  nor U27968(n26573,n23186,n25603);
  nand U27969(n26571,n26538,G59455);
  nand U27970(n26570,n25604,n26539);
  nand U27971(n26569,n21907,n26540);
  nand U27972(G8403,n26576,n26577,n26578,n26579);
  nor U27973(n26579,n26580,n26581,n26582);
  nor U27974(n26582,n21795,n26536);
  nor U27975(n26581,n25612,n26537);
  nor U27976(n26580,n23186,n25613);
  nand U27977(n26578,n26538,G59454);
  nand U27978(n26577,n25614,n26539);
  nand U27979(n26576,n21901,n26540);
  nand U27980(G8402,n26583,n26584,n26585,n26586);
  nor U27981(n26586,n26587,n26588,n26589);
  nor U27982(n26589,n21785,n26536);
  nand U27983(n26536,n26590,n23186,n25623);
  nor U27984(n26588,n25624,n26537);
  nor U27985(n26587,n23186,n25625);
  nand U27986(n26585,n26538,G59453);
  and U27987(n26538,n26591,n26592);
  nand U27988(n26592,n26593,n25629,n26594);
  nand U27989(n26594,G59426,n24656);
  nand U27990(n26593,n26595,n26596);
  nand U27991(n26591,n26597,n25634);
  nand U27992(n26584,n25635,n26539);
  nand U27993(n26539,n26598,n26599);
  or U27994(n26599,n26596,n22383);
  nand U27995(n26598,n26590,G59426);
  not U27996(n26590,n24656);
  nand U27997(n26583,n21896,n26540);
  nand U27998(n26540,n26600,n26601);
  nand U27999(n26601,n26597,n26595);
  nand U28000(n26595,n25640,n26602);
  not U28001(n26597,n26537);
  nand U28002(n26537,n26603,n25642);
  nor U28003(n25642,G59566,G59565);
  or U28004(n26600,n26602,n26596);
  nand U28005(n26596,n26604,n25644);
  nor U28006(n25644,n26605,n26606);
  nand U28007(n26602,n23186,n24656,n25623);
  nand U28008(n23186,n26298,n25992);
  nand U28009(G8401,n26607,n26608,n26609,n26610);
  nor U28010(n26610,n26611,n26612,n26613);
  nor U28011(n26613,n26614,n21845);
  nor U28012(n26612,n26615,n25657);
  nor U28013(n26611,n23111,n26616);
  nand U28014(n26609,n26617,n25660);
  not U28015(n25660,n21848);
  nand U28016(n26608,n25661,n26618);
  nand U28017(n26607,n26619,n25664);
  nand U28018(G8400,n26620,n26621,n26622,n26623);
  nor U28019(n26623,n26624,n26625,n26626);
  nor U28020(n26626,n26614,n21837);
  nor U28021(n26625,n26615,n25672);
  nor U28022(n26624,n23025,n26616);
  nand U28023(n26622,n26617,n25673);
  not U28024(n25673,n21838);
  nand U28025(n26621,n25674,n26618);
  nand U28026(n26620,n26619,n25675);
  nand U28027(G8399,n26627,n26628,n26629,n26630);
  nor U28028(n26630,n26631,n26632,n26633);
  nor U28029(n26633,n26614,n21829);
  nor U28030(n26632,n26615,n25683);
  nor U28031(n26631,n22955,n26616);
  nand U28032(n26629,n26617,n25684);
  not U28033(n25684,n21830);
  nand U28034(n26628,n25685,n26618);
  nand U28035(n26627,n26619,n25686);
  nand U28036(G8398,n26634,n26635,n26636,n26637);
  nor U28037(n26637,n26638,n26639,n26640);
  nor U28038(n26640,n26614,n21821);
  nor U28039(n26639,n26615,n25694);
  nor U28040(n26638,n22876,n26616);
  nand U28041(n26636,n26617,n25695);
  not U28042(n25695,n21822);
  nand U28043(n26635,n25696,n26618);
  nand U28044(n26634,n26619,n25697);
  nand U28045(G8397,n26641,n26642,n26643,n26644);
  nor U28046(n26644,n26645,n26646,n26647);
  nor U28047(n26647,n26614,n21812);
  nor U28048(n26646,n26615,n25705);
  nor U28049(n26645,n22802,n26616);
  nand U28050(n26643,n26617,n25706);
  not U28051(n25706,n21813);
  nand U28052(n26642,n25707,n26618);
  nand U28053(n26641,n26619,n25708);
  nand U28054(G8396,n26648,n26649,n26650,n26651);
  nor U28055(n26651,n26652,n26653,n26654);
  nor U28056(n26654,n26614,n21803);
  nor U28057(n26653,n26615,n25716);
  nor U28058(n26652,n22721,n26616);
  nand U28059(n26650,n26617,n25717);
  not U28060(n25717,n21804);
  nand U28061(n26649,n25718,n26618);
  nand U28062(n26648,n26619,n25719);
  nand U28063(G8395,n26655,n26656,n26657,n26658);
  nor U28064(n26658,n26659,n26660,n26661);
  nor U28065(n26661,n26614,n21794);
  nor U28066(n26660,n26615,n25727);
  nor U28067(n26659,n22645,n26616);
  nand U28068(n26657,n26617,n25728);
  not U28069(n25728,n21795);
  nand U28070(n26656,n25729,n26618);
  nand U28071(n26655,n26619,n25730);
  nand U28072(G8394,n26662,n26663,n26664,n26665);
  nor U28073(n26665,n26666,n26667,n26668);
  nor U28074(n26668,n26614,n21784);
  and U28075(n26614,n26669,n26670);
  nand U28076(n26670,n25623,n26671,n23160,n24667);
  nand U28077(n26671,n26672,n26673);
  nand U28078(n26669,n26619,n25743);
  nor U28079(n26667,n26615,n25744);
  and U28080(n26615,n26674,n26675);
  or U28081(n26675,n26673,n22383);
  nand U28082(n26674,n26676,G59426);
  nor U28083(n26666,n22527,n26616);
  nand U28084(n26616,n26677,n26678);
  nand U28085(n26678,n26679,n25629,n26680);
  nand U28086(n26680,n25743,n26673);
  nand U28087(n26679,n26681,n24667);
  nand U28088(n26681,n26682,n21044);
  nand U28089(n26682,n26673,n23160);
  nand U28090(n26673,n26604,n25754);
  nor U28091(n25754,n26605,G59566);
  nand U28092(n26677,n26619,n25634);
  nand U28093(n26664,n26617,n25755);
  not U28094(n25755,n21785);
  and U28095(n26617,n25623,n26676);
  not U28096(n26676,n24667);
  nand U28097(n26663,n25756,n26618);
  not U28098(n26618,n23160);
  nand U28099(n23160,n26298,n26068);
  nor U28100(n26298,n26069,n26683);
  not U28101(n25756,n25625);
  nand U28102(n26662,n26619,n25758);
  not U28103(n26619,n26672);
  nand U28104(n26672,n26603,n25759);
  nand U28105(G8393,n26684,n26685,n26686,n26687);
  nor U28106(n26687,n26688,n26689,n26690);
  nor U28107(n26690,n21848,n26691);
  nor U28108(n26689,n25548,n26692);
  nor U28109(n26688,n23159,n25550);
  nand U28110(n26686,n26693,G59444);
  nand U28111(n26685,n25552,n26694);
  nand U28112(n26684,n21932,n26695);
  nand U28113(G8392,n26696,n26697,n26698,n26699);
  nor U28114(n26699,n26700,n26701,n26702);
  nor U28115(n26702,n21838,n26691);
  nor U28116(n26701,n25562,n26692);
  nor U28117(n26700,n23159,n25563);
  nand U28118(n26698,n26693,G59443);
  nand U28119(n26697,n25564,n26694);
  nand U28120(n26696,n21927,n26695);
  nand U28121(G8391,n26703,n26704,n26705,n26706);
  nor U28122(n26706,n26707,n26708,n26709);
  nor U28123(n26709,n21830,n26691);
  nor U28124(n26708,n25572,n26692);
  nor U28125(n26707,n23159,n25573);
  nand U28126(n26705,n26693,G59442);
  nand U28127(n26704,n25574,n26694);
  nand U28128(n26703,n21922,n26695);
  nand U28129(G8390,n26710,n26711,n26712,n26713);
  nor U28130(n26713,n26714,n26715,n26716);
  nor U28131(n26716,n21822,n26691);
  nor U28132(n26715,n25582,n26692);
  nor U28133(n26714,n23159,n25583);
  nand U28134(n26712,n26693,G59441);
  nand U28135(n26711,n25584,n26694);
  nand U28136(n26710,n21917,n26695);
  nand U28137(G8389,n26717,n26718,n26719,n26720);
  nor U28138(n26720,n26721,n26722,n26723);
  nor U28139(n26723,n21813,n26691);
  nor U28140(n26722,n25592,n26692);
  nor U28141(n26721,n23159,n25593);
  nand U28142(n26719,n26693,G59440);
  nand U28143(n26718,n25594,n26694);
  nand U28144(n26717,n21912,n26695);
  nand U28145(G8388,n26724,n26725,n26726,n26727);
  nor U28146(n26727,n26728,n26729,n26730);
  nor U28147(n26730,n21804,n26691);
  nor U28148(n26729,n25602,n26692);
  nor U28149(n26728,n23159,n25603);
  nand U28150(n26726,n26693,G59439);
  nand U28151(n26725,n25604,n26694);
  nand U28152(n26724,n21907,n26695);
  nand U28153(G8387,n26731,n26732,n26733,n26734);
  nor U28154(n26734,n26735,n26736,n26737);
  nor U28155(n26737,n21795,n26691);
  nor U28156(n26736,n25612,n26692);
  nor U28157(n26735,n23159,n25613);
  nand U28158(n26733,n26693,G59438);
  nand U28159(n26732,n25614,n26694);
  nand U28160(n26731,n21901,n26695);
  nand U28161(G8386,n26738,n26739,n26740,n26741);
  nor U28162(n26741,n26742,n26743,n26744);
  nor U28163(n26744,n21785,n26691);
  nand U28164(n26691,n26745,n23159,n25623);
  nor U28165(n26743,n25624,n26692);
  nor U28166(n26742,n23159,n25625);
  nand U28167(n26740,n26693,G59437);
  and U28168(n26693,n26746,n26747);
  nand U28169(n26747,n26748,n25629,n26749);
  nand U28170(n26749,G59426,n24657);
  nand U28171(n26748,n26750,n26751);
  nand U28172(n26746,n26752,n25634);
  nand U28173(n26739,n25635,n26694);
  nand U28174(n26694,n26753,n26754);
  or U28175(n26754,n26751,n22383);
  nand U28176(n26753,n26745,G59426);
  not U28177(n26745,n24657);
  nand U28178(n26738,n21896,n26695);
  nand U28179(n26695,n26755,n26756);
  nand U28180(n26756,n26752,n26750);
  nand U28181(n26750,n25640,n26757);
  not U28182(n26752,n26692);
  nand U28183(n26692,n26603,n25834);
  or U28184(n26755,n26757,n26751);
  nand U28185(n26751,n26604,n25835);
  nor U28186(n25835,n26606,n26758);
  nand U28187(n26757,n23159,n24657,n25623);
  nand U28188(n23159,n26449,n25992);
  nor U28189(n25992,n26450,n26528);
  nand U28190(G8385,n26759,n26760,n26761,n26762);
  nor U28191(n26762,n26763,n26764,n26765);
  nor U28192(n26765,n21848,n26766);
  nand U28193(n21848,n26767,n26768);
  or U28194(n26768,n21776,G58855);
  nand U28195(n26767,n21776,n26769);
  nor U28196(n26764,n25548,n26770);
  not U28197(n25548,n25664);
  nand U28198(n25664,n26771,n26772);
  nand U28199(n26772,n26773,n21846);
  nand U28200(n26771,n25552,G59426);
  nor U28201(n26763,n26774,n25657);
  not U28202(n25657,n25552);
  nor U28203(n25552,n21845,n25538);
  nand U28204(n26761,n26775,G59436);
  nand U28205(n26760,n21932,n26776);
  not U28206(n21932,n21845);
  nand U28207(n21845,n26777,n26778);
  or U28208(n26778,n21776,G58839);
  nand U28209(n26777,n21776,n26779);
  nand U28210(n26759,n25661,n26780);
  not U28211(n25661,n25550);
  nand U28212(n25550,n26781,n26782,n25623);
  nand U28213(n26782,n21774,n21775);
  nand U28214(n26781,n21776,n21772);
  nand U28215(G8384,n26783,n26784,n26785,n26786);
  nor U28216(n26786,n26787,n26788,n26789);
  nor U28217(n26789,n21838,n26766);
  nand U28218(n21838,n26790,n26791);
  or U28219(n26791,n21776,G58856);
  nand U28220(n26790,n21776,n26792);
  nor U28221(n26788,n25562,n26770);
  not U28222(n25562,n25675);
  nand U28223(n25675,n26793,n26794);
  nand U28224(n26794,n26773,n21057);
  nand U28225(n26793,n25564,G59426);
  nor U28226(n26787,n26774,n25672);
  not U28227(n25672,n25564);
  nor U28228(n25564,n21837,n25538);
  nand U28229(n26785,n26775,G59435);
  nand U28230(n26784,n21927,n26776);
  not U28231(n21927,n21837);
  nand U28232(n21837,n26795,n26796);
  or U28233(n26796,n21776,G58840);
  nand U28234(n26795,n21776,n26797);
  nand U28235(n26783,n25674,n26780);
  not U28236(n25674,n25563);
  nand U28237(n25563,n26798,n26799,n25623);
  nand U28238(n26799,n21774,n21763);
  nand U28239(n26798,n21776,n21762);
  nand U28240(G8383,n26800,n26801,n26802,n26803);
  nor U28241(n26803,n26804,n26805,n26806);
  nor U28242(n26806,n21830,n26766);
  nand U28243(n21830,n26807,n26808);
  or U28244(n26808,n21776,G58857);
  nand U28245(n26807,n21776,n26809);
  nor U28246(n26805,n25572,n26770);
  not U28247(n25572,n25686);
  nand U28248(n25686,n26810,n26811);
  nand U28249(n26811,n26773,n21849);
  nand U28250(n26810,n25574,G59426);
  nor U28251(n26804,n26774,n25683);
  not U28252(n25683,n25574);
  nor U28253(n25574,n21829,n25538);
  nand U28254(n26802,n26775,G59434);
  nand U28255(n26801,n21922,n26776);
  not U28256(n21922,n21829);
  nand U28257(n21829,n26812,n26813);
  or U28258(n26813,n21776,G58841);
  nand U28259(n26812,n21776,n26814);
  nand U28260(n26800,n25685,n26780);
  not U28261(n25685,n25573);
  nand U28262(n25573,n26815,n26816,n25623);
  nand U28263(n26816,n21774,n21753);
  nand U28264(n26815,n21776,n21752);
  nand U28265(G8382,n26817,n26818,n26819,n26820);
  nor U28266(n26820,n26821,n26822,n26823);
  nor U28267(n26823,n21822,n26766);
  nand U28268(n21822,n26824,n26825);
  or U28269(n26825,n21776,G58858);
  nand U28270(n26824,n21776,n26826);
  nor U28271(n26822,n25582,n26770);
  not U28272(n25582,n25697);
  nand U28273(n25697,n26827,n26828);
  nand U28274(n26828,n26773,n21687);
  nand U28275(n26827,n25584,G59426);
  nor U28276(n26821,n26774,n25694);
  not U28277(n25694,n25584);
  nor U28278(n25584,n21821,n25538);
  nand U28279(n26819,n26775,G59433);
  nand U28280(n26818,n21917,n26776);
  not U28281(n21917,n21821);
  nand U28282(n21821,n26829,n26830);
  or U28283(n26830,n21776,G58842);
  nand U28284(n26829,n21776,n26831);
  nand U28285(n26817,n25696,n26780);
  not U28286(n25696,n25583);
  nand U28287(n25583,n26832,n26833,n25623);
  nand U28288(n26833,n21774,n21743);
  nand U28289(n26832,n21776,n21742);
  nand U28290(G8381,n26834,n26835,n26836,n26837);
  nor U28291(n26837,n26838,n26839,n26840);
  nor U28292(n26840,n21813,n26766);
  nand U28293(n21813,n26841,n26842);
  or U28294(n26842,n21776,G58859);
  nand U28295(n26841,n21776,n26843);
  nor U28296(n26839,n25592,n26770);
  not U28297(n25592,n25708);
  nand U28298(n25708,n26844,n26845);
  nand U28299(n26845,n26773,n25522);
  nand U28300(n26844,n25594,G59426);
  nor U28301(n26838,n26774,n25705);
  not U28302(n25705,n25594);
  nor U28303(n25594,n21812,n25538);
  nand U28304(n26836,n26775,G59432);
  nand U28305(n26835,n21912,n26776);
  not U28306(n21912,n21812);
  nand U28307(n21812,n26846,n26847);
  or U28308(n26847,n21776,G58843);
  nand U28309(n26846,n21776,n26848);
  nand U28310(n26834,n25707,n26780);
  not U28311(n25707,n25593);
  nand U28312(n25593,n26849,n26850,n25623);
  nand U28313(n26850,n21774,n21733);
  nand U28314(n26849,n21776,n21732);
  nand U28315(G8380,n26851,n26852,n26853,n26854);
  nor U28316(n26854,n26855,n26856,n26857);
  nor U28317(n26857,n21804,n26766);
  nand U28318(n21804,n26858,n26859);
  or U28319(n26859,n21776,G58860);
  nand U28320(n26858,n21776,n26860);
  nor U28321(n26856,n25602,n26770);
  not U28322(n25602,n25719);
  nand U28323(n25719,n26861,n26862);
  nand U28324(n26862,n26773,n26863);
  nand U28325(n26861,n25604,G59426);
  nor U28326(n26855,n26774,n25716);
  not U28327(n25716,n25604);
  nor U28328(n25604,n21803,n25538);
  nand U28329(n26853,n26775,G59431);
  nand U28330(n26852,n21907,n26776);
  not U28331(n21907,n21803);
  nand U28332(n21803,n26864,n26865);
  or U28333(n26865,n21776,G58844);
  nand U28334(n26864,n21776,n26866);
  nand U28335(n26851,n25718,n26780);
  not U28336(n25718,n25603);
  nand U28337(n25603,n26867,n26868,n25623);
  nand U28338(n26868,n21774,n21723);
  nand U28339(n26867,n21776,n21722);
  nand U28340(G8379,n26869,n26870,n26871,n26872);
  nor U28341(n26872,n26873,n26874,n26875);
  nor U28342(n26875,n21795,n26766);
  nand U28343(n21795,n26876,n26877);
  or U28344(n26877,n21776,G58861);
  nand U28345(n26876,n21776,n26878);
  nor U28346(n26874,n25612,n26770);
  not U28347(n25612,n25730);
  nand U28348(n25730,n26879,n26880);
  nand U28349(n26880,n26773,n21534);
  nand U28350(n26879,n25614,G59426);
  nor U28351(n26873,n26774,n25727);
  not U28352(n25727,n25614);
  nor U28353(n25614,n21794,n25538);
  nand U28354(n26871,n26775,G59430);
  nand U28355(n26870,n21901,n26776);
  not U28356(n21901,n21794);
  nand U28357(n21794,n26881,n26882);
  or U28358(n26882,n21776,G58845);
  nand U28359(n26881,n21776,n26883);
  nand U28360(n26869,n25729,n26780);
  not U28361(n26780,n23170);
  not U28362(n25729,n25613);
  nand U28363(n25613,n26884,n26885,n25623);
  nand U28364(n26885,n21774,n21711);
  nand U28365(n26884,n21776,n21709);
  nand U28366(G8378,n26886,n26887,n26888,n26889);
  nor U28367(n26889,n26890,n26891,n26892);
  nor U28368(n26892,n25624,n26770);
  not U28369(n25624,n25758);
  nand U28370(n25758,n26893,n26894);
  nand U28371(n26894,n26773,n26895);
  nor U28372(n26773,n21047,n25538);
  nand U28373(n26893,n25635,G59426);
  nor U28374(n26891,n26774,n25744);
  not U28375(n25744,n25635);
  nor U28376(n25635,n21784,n25538);
  and U28377(n26774,n26896,n26897);
  nand U28378(n26897,n26898,n22435);
  nand U28379(n26896,n26899,G59426);
  nor U28380(n26890,n23170,n25625);
  nand U28381(n25625,n26900,n26901,n25623);
  nand U28382(n26901,n21774,n26902);
  or U28383(n26900,n21774,G58902);
  not U28384(n21774,n21776);
  or U28385(n26888,n26766,n21785);
  nand U28386(n21785,n26903,n26904);
  or U28387(n26904,n21776,G58862);
  nand U28388(n26903,n21776,n26905);
  nand U28389(n26766,n25623,n26899);
  not U28390(n26899,n24658);
  nand U28391(n26887,n21896,n26776);
  nand U28392(n26776,n26906,n26907);
  nand U28393(n26907,n25623,n23170,n26898);
  not U28394(n26898,n26908);
  nand U28395(n26906,n26909,n26910);
  not U28396(n21896,n21784);
  nand U28397(n21784,n26911,n26912);
  or U28398(n26912,n21776,G58846);
  nand U28399(n26911,n21776,n26913);
  nand U28400(n26886,n26775,G59429);
  and U28401(n26775,n26914,n26915);
  nand U28402(n26915,n26916,n25629,n26917);
  nand U28403(n26917,G59426,n24658);
  nor U28404(n25629,n25538,n21075);
  nand U28405(n26916,n26910,n26908);
  nand U28406(n26908,n26604,n25911);
  nor U28407(n25911,G59566,n26758);
  nor U28408(n26604,n26219,n26526);
  not U28409(n26219,n25913);
  nand U28410(n26910,n25640,n26918);
  nand U28411(n26918,n23170,n24658,n25623);
  nand U28412(n23170,n26449,n26068);
  nor U28413(n26068,n26450,n26451);
  nor U28414(n26449,n26683,n26221);
  not U28415(n25640,n25743);
  nor U28416(n25743,n22383,n25538);
  nand U28417(n26914,n26909,n25634);
  nand U28418(n25634,n26920,n26921,n26922);
  or U28419(n26922,n21019,n21031);
  nand U28420(n26921,n21046,n26923);
  nand U28421(n26920,n21044,n21531,G59427);
  not U28422(n26909,n26770);
  nand U28423(n26770,n26603,n25915);
  nor U28424(n26603,n26924,n26925);
  nand U28425(G8377,n21555,n26926,n26927,n26928);
  nand U28426(n26928,n26929,G59428);
  nand U28427(n26927,n26930,n26931);
  nand U28428(n26930,n26932,n26933,n26934);
  nand U28429(n26934,n26935,n21080);
  nand U28430(n26933,n26936,n21531);
  nand U28431(n26936,G59425,n21080,n21075);
  nand U28432(n26932,n20985,n26937);
  nand U28433(n21555,G59425,G59428,n21075);
  nand U28434(G8376,n26938,n21554,n26939);
  nand U28435(n26939,G59427,n26940);
  nand U28436(n26940,n26931,n26926);
  nand U28437(n26926,G59428,n21044,n21944);
  nand U28438(n21554,n21044,n21531,n22435);
  nand U28439(n26938,n26941,n26931);
  nand U28440(n26941,n21563,n26942);
  nand U28441(n26942,n21045,n21043,n22385);
  not U28442(n21563,n21022);
  nor U28443(n21022,n22166,n21531);
  nand U28444(G8375,n22166,n25533,n26943,n26944);
  or U28445(n26944,n26919,G59428);
  nand U28446(n26943,n21045,n21044,G59427,G59428);
  nand U28447(G8374,n26945,n21019,n26946);
  nand U28448(n26946,n26929,G59425);
  not U28449(n26929,n26931);
  nand U28450(n26931,n26947,n26948,n26949);
  nand U28451(n26949,n26950,n21531);
  nand U28452(n26950,n21944,G59427);
  nand U28453(n26948,n22165,n21060,n21538);
  nor U28454(n21538,G59797,n21944);
  nand U28455(n26947,n26951,n25533);
  or U28456(n26951,n26937,n22166);
  not U28457(n22166,n20985);
  nor U28458(n20985,n21044,G59427);
  nand U28459(n26937,n26952,n26953,n26954,n26955);
  nor U28460(n26955,n26956,n26957,n26958,n26959);
  and U28461(n26959,n20986,n20987);
  xnor U28462(n20986,n26960,n24857);
  and U28463(n24857,n26961,n26962);
  nand U28464(n26961,n26963,n26964);
  nand U28465(n26960,n24858,n24855);
  nand U28466(n24855,n26965,n26966);
  or U28467(n24858,n26966,n26965);
  nor U28468(n26965,n21114,n23419);
  xor U28469(n26966,n26967,n22435);
  nand U28470(n26967,n26968,n26969,n26970,n26971);
  nor U28471(n26971,n26972,n26973);
  nor U28472(n26973,n22382,n22354);
  nor U28473(n26972,n22167,n24870);
  not U28474(n24870,G59762);
  nand U28475(n26970,G59571,n22496);
  nand U28476(n26969,G59557,n26974);
  nand U28477(n26974,n21943,n26975);
  nand U28478(n26975,n22049,G59428);
  nand U28479(n26968,n21674,n22497);
  not U28480(n21674,n21484);
  xnor U28481(n21484,n24851,n24850);
  xnor U28482(n24851,n21108,n26976);
  nor U28483(n26976,n26977,n26978,n26979,n26980);
  and U28484(n26980,n22437,G59698);
  and U28485(n26979,n22436,G59571);
  nor U28486(n26978,n22383,n22354);
  not U28487(n22354,G59603);
  nor U28488(n26977,n24241,n21485);
  not U28489(n21485,G59730);
  not U28490(n24241,n22434);
  nor U28491(n26958,n24880,n21023);
  nor U28492(n26957,n25512,n25492);
  nor U28493(n26956,n26981,n26982);
  nor U28494(n26954,n22386,n26983);
  nor U28495(n26983,n26984,n21101);
  nand U28496(n21101,n21091,n26985);
  nand U28497(n26985,n26986,n21045);
  nand U28498(n26986,n26987,n21059,n26988);
  nand U28499(n26988,n22163,n21849);
  and U28500(n21091,n26989,n26990,n26991,n26992);
  nand U28501(n26991,n24879,n26993);
  nand U28502(n26993,n26994,n26995);
  nor U28503(n26989,n26996,n26997);
  nor U28504(n26997,n25517,n21080);
  nor U28505(n26996,n25512,n26987);
  not U28506(n25512,n21105);
  nor U28507(n26984,G59795,G59796);
  nand U28508(n26953,n26998,n25536);
  nand U28509(n26998,n26999,n27000);
  nand U28510(n27000,n27001,n26924,n27002);
  not U28511(n27002,n26982);
  nand U28512(n26999,n27003,n26925);
  nand U28513(n27003,n26982,n27004);
  nand U28514(n27004,n27005,n27001);
  nand U28515(n27001,n27006,n27007,n27008,n27009);
  nand U28516(n27009,n27010,n27011);
  nand U28517(n27011,n27012,n27013);
  nand U28518(n27013,G59560,n27014);
  nand U28519(n27008,n27015,n21013,n21023);
  nand U28520(n21013,n27016,n27017,n27018,n27019);
  nor U28521(n27019,n27020,n27021,n27022);
  nor U28522(n27022,n27023,n26221);
  nor U28523(n27021,n27024,n27025);
  nor U28524(n27024,n24369,n23146);
  not U28525(n23146,n23143);
  nor U28526(n23143,n27026,n24362);
  nor U28527(n27026,n24388,n21058);
  nor U28528(n27020,n25395,n25491);
  nor U28529(n25395,n24362,n24369);
  nand U28530(n27018,n21521,n27027);
  nand U28531(n27017,n21015,n27028);
  not U28532(n21015,n21520);
  xnor U28533(n21520,n27029,n27030);
  and U28534(n27030,n27031,n27032);
  nand U28535(n27016,n21014,n27033);
  or U28536(n27015,n21027,n27014);
  not U28537(n27014,n25915);
  nand U28538(n27007,n27034,n27035);
  nand U28539(n27034,n27036,n27037,G59566);
  nand U28540(n27037,n27010,G59561);
  nand U28541(n27036,n21027,n21023);
  nand U28542(n21027,n27038,n27039,n27040,n27041);
  nor U28543(n27041,n27042,n27043);
  nor U28544(n27043,n27044,n25481);
  not U28545(n25481,n21084);
  nor U28546(n27042,n27045,n21029);
  nand U28547(n27040,n21030,n27028);
  xor U28548(n21030,n27046,n22383);
  nand U28549(n27046,n27047,n27048);
  nand U28550(n27039,n27049,n23142);
  nand U28551(n27038,n26528,n27050);
  or U28552(n27006,n26981,G59564);
  nand U28553(n27005,G59564,n26981);
  nand U28554(n26981,n27051,n27052);
  nand U28555(n27052,n27010,n27053);
  or U28556(n27051,n21004,n27010);
  nand U28557(n21004,n27054,n27055,n27056,n27057);
  nor U28558(n27057,n27058,n27059,n27060);
  nor U28559(n27060,n25491,n25403);
  xor U28560(n25403,n27061,n27012);
  not U28561(n27012,n24361);
  nor U28562(n27059,n27023,n26450);
  nor U28563(n27058,n27045,n27062);
  nand U28564(n27056,n23115,n25354);
  xor U28565(n23115,G59559,n27063);
  nand U28566(n27055,n21510,n27027);
  nand U28567(n27054,n21006,n27028);
  not U28568(n21006,n21508);
  nand U28569(n21508,n27064,n27065);
  nand U28570(n27065,n27066,n27067);
  not U28571(n27066,n27068);
  nand U28572(n27064,n27069,n27032,n27070);
  nand U28573(n27069,n27071,n27067);
  nand U28574(n26982,n27072,n27073);
  nand U28575(n27073,n27010,n24998);
  or U28576(n27072,n20997,n27010);
  not U28577(n27010,n21023);
  nand U28578(n21023,n27074,n27075,n25508);
  and U28579(n25508,n27076,n27077,n27078,n27079);
  nor U28580(n27079,n27080,n27081);
  xnor U28581(n27081,n26995,n27082);
  not U28582(n27080,n26990);
  nor U28583(n26990,n27083,n27084,n25368,n27085);
  and U28584(n27083,n27086,n21849);
  nand U28585(n27086,n27087,n21534,n21058);
  not U28586(n27077,n27088);
  nand U28587(n27076,n21933,n27089);
  nand U28588(n27089,n22163,n25522);
  nand U28589(n27075,n27090,n21045);
  nand U28590(n27090,n27091,n27092);
  nand U28591(n27092,n27093,n21080);
  nand U28592(n27093,n25497,n27094);
  nand U28593(n27094,n21060,n27095);
  nand U28594(n27095,n21562,n25496);
  not U28595(n25496,n22049);
  not U28596(n21060,n21059);
  nand U28597(n21059,n22050,n25365);
  or U28598(n27091,n25492,n21105);
  nand U28599(n21105,n27096,n27097);
  nand U28600(n27097,n27098,n27099,n27100,n27101);
  nand U28601(n27101,n27102,n27103,n27104);
  or U28602(n27104,n27105,n21057);
  nand U28603(n27103,n27106,n27107,n27108);
  not U28604(n27108,n27109);
  not U28605(n27107,n25237);
  nand U28606(n27106,n27110,n27111);
  or U28607(n27102,n27111,n27110);
  nand U28608(n27100,n27105,n21057);
  not U28609(n27098,n27112);
  nand U28610(n27074,n27049,n21080);
  nand U28611(n20997,n27113,n27114,n27115,n27116);
  nor U28612(n27116,n27117,n27118,n27119);
  nor U28613(n27119,n25491,n25394);
  nand U28614(n25394,n27120,n27121,n27122);
  nand U28615(n27122,n27123,n21846);
  or U28616(n27121,n27124,n24998);
  nand U28617(n27120,n27125,n27124);
  nand U28618(n27124,n27061,n24361);
  xnor U28619(n27061,n21058,G59559);
  nand U28620(n27125,n27126,n27127);
  nand U28621(n27127,n21058,n24998);
  nor U28622(n27118,n27044,n22361);
  not U28623(n22361,n21498);
  not U28624(n27044,n27027);
  nand U28625(n27027,n27128,n25501,n27129,n25499);
  nand U28626(n25499,n27130,n25522);
  nor U28627(n27129,n25505,n27131);
  nor U28628(n27131,n22163,n27132);
  nor U28629(n25505,n21935,n25522);
  not U28630(n21935,n22473);
  not U28631(n27128,n25503);
  nand U28632(n25503,n21562,n27133,n27134,n27135);
  nand U28633(n27135,n25237,n21058);
  nand U28634(n27134,n27136,n21846);
  nand U28635(n27136,n27137,n27138);
  nand U28636(n27138,n21688,n27139);
  nand U28637(n27139,n27085,n27140);
  nand U28638(n27140,n26987,n21057);
  nand U28639(n27137,n25368,n26987);
  not U28640(n26987,n25517);
  nor U28641(n25517,n21849,n22163);
  nand U28642(n27133,n25368,n27141);
  nand U28643(n27141,n25487,n27082);
  nor U28644(n27117,n27045,n27142);
  not U28645(n27045,n27033);
  nand U28646(n27033,n27143,n25492);
  nand U28647(n27115,n20996,n27028);
  nand U28648(n27028,n25494,n25495,n25490,n25497);
  not U28649(n25497,n20987);
  not U28650(n25495,n27144);
  xnor U28651(n20996,n26963,n27145);
  and U28652(n27145,n26964,n26962);
  nand U28653(n26962,n27146,n27147,n27148);
  nand U28654(n27148,n21691,G59553);
  nand U28655(n26964,G59553,n27149,n21691);
  nand U28656(n27149,n27146,n27147);
  or U28657(n27147,n27150,n22383);
  nand U28658(n27146,n27150,n22383);
  nand U28659(n27150,n27151,n27152,n27153,n27154);
  nor U28660(n27154,n27155,n27156);
  nor U28661(n27156,n22382,n21494);
  nor U28662(n27155,n22167,n21497);
  not U28663(n21497,G59761);
  nand U28664(n27153,G59558,n27157);
  nand U28665(n27152,n21498,n22497);
  nor U28666(n21498,n27158,n24850);
  nor U28667(n24850,n27159,n27160);
  and U28668(n27158,n27160,n27159);
  xor U28669(n27160,n27161,n22167);
  nand U28670(n27161,n27162,n27163,n27164,n27165);
  nor U28671(n27165,n27166,n27167,n27168,n27169);
  nor U28672(n27169,n22383,n21494);
  not U28673(n21494,G59602);
  and U28674(n27168,n22434,G59729);
  nor U28675(n27167,n27170,n24998);
  nor U28676(n27166,n26683,n26919);
  not U28677(n26683,n26070);
  nor U28678(n27164,n27171,n27172);
  and U28679(n27172,n22437,G59697);
  nor U28680(n27171,n22508,n24866);
  not U28681(n24866,G59570);
  nand U28682(n27163,n21075,G59563);
  nand U28683(n27162,n25535,n21046);
  nand U28684(n27151,G59570,n22496);
  and U28685(n26963,n27067,n27068);
  nand U28686(n27068,n27071,n27173);
  nand U28687(n27173,n27070,n27032);
  nand U28688(n27032,n27174,n27175);
  nand U28689(n27175,n27176,n27177);
  nand U28690(n27070,n27029,n27031);
  nand U28691(n27031,n27176,n27177,n27178);
  not U28692(n27178,n27174);
  nand U28693(n27174,n22167,n25533,n27179,n27180);
  nor U28694(n27180,n27181,n27182,n27183);
  nor U28695(n27183,n22163,n27184);
  nor U28696(n27182,n23050,n21114);
  nand U28697(n27179,n25236,n27185,n26994,G59428);
  and U28698(n25236,n25365,n21846,n26995);
  or U28699(n27177,n27186,n22383);
  nand U28700(n27176,n22383,n27186);
  nand U28701(n27186,n27187,n27188,n27189,n27190);
  nor U28702(n27190,n27191,n27192);
  nor U28703(n27192,n22382,n21519);
  nor U28704(n27191,n22167,n21130);
  not U28705(n21130,G59759);
  nand U28706(n27189,n21521,n22497);
  not U28707(n21521,n22375);
  xor U28708(n22375,n27193,n27194);
  nand U28709(n27193,n27195,n27196);
  nand U28710(n27188,G59568,n22496);
  nand U28711(n27187,G59560,n27157);
  nand U28712(n27029,n27048,n27197);
  nand U28713(n27197,n22435,n27047);
  nand U28714(n27047,n27198,n27199,n27200);
  not U28715(n27200,n27201);
  nand U28716(n27048,n27201,n27202);
  nand U28717(n27202,n27198,n27199);
  or U28718(n27199,n27203,n22383);
  nand U28719(n27198,n27203,n22383);
  nand U28720(n27203,n27204,n27205,n27206,n27207);
  nor U28721(n27207,n27208,n27209);
  nor U28722(n27209,n22382,n21530);
  nor U28723(n27208,n22167,n21122);
  not U28724(n21122,G59758);
  nand U28725(n27206,G59561,n27157);
  nand U28726(n27205,n21084,n22497);
  nand U28727(n21084,n27210,n27211);
  nand U28728(n27211,n27212,n27213);
  nand U28729(n27212,n27214,n27215);
  nand U28730(n27215,n27216,n22167);
  or U28731(n27210,n27213,n22167);
  nand U28732(n27204,G59567,n22496);
  nand U28733(n27201,n27217,n27218,n27219,n21047);
  nand U28734(n27218,G59428,n27220);
  nand U28735(n27220,n27221,n26895,n27222,n27223);
  nor U28736(n27223,n27224,n27225,n27226,n27227);
  nor U28737(n27225,n27228,n27229);
  nor U28738(n27229,n27230,n27231);
  nor U28739(n27231,n21688,n26863);
  nor U28740(n27230,n22163,n21080);
  nor U28741(n27224,n21687,n21534);
  nand U28742(n27222,n21933,n27087);
  not U28743(n27221,n27130);
  nand U28744(n27217,n21691,G59556);
  nand U28745(n27071,n27232,n27233,n27219,n26919);
  xnor U28746(n27232,n22435,n27234);
  nand U28747(n27067,n27235,n27236);
  nand U28748(n27236,n27219,n26919,n27233);
  nand U28749(n27233,n21691,G59554);
  xnor U28750(n27235,n27234,n22383);
  nand U28751(n27234,n27237,n27238,n27239,n27240);
  nand U28752(n27240,G59559,n27157);
  nand U28753(n27157,n21943,n21939,n21047,n27241);
  nor U28754(n27241,n27242,n27243,n27244);
  nor U28755(n27244,n22163,n21531,n25489,n21080);
  not U28756(n25489,n22386);
  nor U28757(n27243,n27245,n21531);
  nor U28758(n27245,n22049,n27144);
  nor U28759(n27144,n27246,n21846);
  nor U28760(n27242,n21531,n25494);
  not U28761(n21939,n22437);
  nor U28762(n27239,n27247,n27248);
  nor U28763(n27248,n22446,n24982);
  not U28764(n22446,n22496);
  and U28765(n27250,n27251,n27252,n27219);
  nand U28766(n27219,G59428,n21534,n25516,n27253);
  and U28767(n27253,n27185,n24531);
  nor U28768(n24531,n21069,n21058);
  nand U28769(n27249,G59428,n25504);
  nand U28770(n25504,n27143,n27254);
  and U28771(n27143,n27255,n27256);
  nand U28772(n27256,n27130,n27257,n27085);
  or U28773(n27255,n27246,n21058);
  and U28774(n27247,n22497,n21510);
  not U28775(n21510,n22368);
  nand U28776(n22368,n27258,n27159);
  nand U28777(n27159,n27259,n27260);
  nand U28778(n27260,n27261,n27195);
  xnor U28779(n27259,n27262,n22167);
  nand U28780(n27258,n27261,n27195,n27263);
  xnor U28781(n27263,n21108,n27262);
  nand U28782(n27262,n27264,n27265,n27266,n27267);
  nor U28783(n27267,n27268,n27269,n27270,n27271);
  nor U28784(n27271,n27062,n25533);
  nor U28785(n27270,n26919,n26450);
  nand U28786(n26450,n27272,n27273);
  nand U28787(n27273,n27274,n27275);
  nand U28788(n27274,n27276,n27277);
  nand U28789(n27272,n27278,n21061);
  xor U28790(n27278,n27279,n27280);
  nor U28791(n27269,n26924,n21047);
  and U28792(n27268,n22437,G59696);
  nor U28793(n27266,n27281,n27282);
  nor U28794(n27282,n22508,n24982);
  not U28795(n24982,G59569);
  nor U28796(n27281,n22383,n21507);
  not U28797(n21507,G59601);
  nand U28798(n27265,G59559,n27283);
  nand U28799(n27264,G59728,n22434);
  nand U28800(n27195,n27284,n27285);
  nand U28801(n27285,n27252,n22383,n21113,n27286);
  and U28802(n27286,n27287,n27288);
  xnor U28803(n27284,n27289,n22167);
  nand U28804(n27261,n27196,n27194);
  nand U28805(n27194,n27213,n27290);
  nand U28806(n27290,n21108,n27214);
  nand U28807(n27214,n27291,n27292);
  not U28808(n27291,n27216);
  nand U28809(n27213,n27293,n27216);
  nand U28810(n27216,n22382,n27294,n21113,n21047);
  nand U28811(n27294,G59428,n27295);
  nand U28812(n27295,n27296,n27297,n27298,n27299);
  nor U28813(n27299,n27300,n27301,n27302);
  nor U28814(n27302,n21688,n27303);
  nor U28815(n27301,n25516,n27304,n27305);
  nor U28816(n27305,n21688,n26995);
  nor U28817(n27304,n27228,n26863);
  nor U28818(n27300,n21849,n25487);
  not U28819(n27298,n27226);
  nand U28820(n27226,n27306,n27307,n27308,n27309);
  nor U28821(n27309,n27088,n27084);
  nand U28822(n27308,n26995,n21849);
  nand U28823(n27307,n21688,n21846);
  nand U28824(n27306,n26994,n21058);
  nand U28825(n27297,n21933,n21057);
  nand U28826(n27296,n27085,n22163);
  not U28827(n22382,n23278);
  xnor U28828(n27293,n27292,n22167);
  nand U28829(n27292,n27310,n27311);
  nor U28830(n27311,n27312,n27313,n27314,n27315);
  nor U28831(n27315,n26919,n26451);
  not U28832(n26451,n26528);
  nor U28833(n26528,n27316,n27317);
  nor U28834(n27317,n21073,n27318);
  and U28835(n27318,G59561,n27319);
  nor U28836(n27314,n22383,n21530);
  not U28837(n21530,G59599);
  and U28838(n27313,n22434,G59726);
  nor U28839(n27312,n27170,n23142);
  nor U28840(n27310,n27320,n27321,n27322,n27323);
  nor U28841(n27323,n25533,n21029);
  nor U28842(n27322,n26606,n21047);
  and U28843(n27321,n22437,G59694);
  nor U28844(n27320,n22508,n25224);
  nand U28845(n27196,n27324,n27287,n27288,n27325);
  not U28846(n22051,n27252);
  not U28847(n27288,n27181);
  nand U28848(n27181,n21943,n27326);
  nand U28849(n27326,G59428,n21534,n27327);
  nand U28850(n27287,n27130,n27257,G59428,n25365);
  xnor U28851(n27324,n21108,n27289);
  nand U28852(n27289,n27328,n27329);
  nor U28853(n27329,n27330,n27331,n27332,n27333);
  nor U28854(n27333,n22383,n21519);
  not U28855(n21519,G59600);
  and U28856(n27332,n22434,G59727);
  nand U28857(n22434,n22167,n27334);
  nand U28858(n27334,n21692,G59428);
  nor U28859(n27331,n27170,n24388);
  not U28860(n27170,n27283);
  nand U28861(n27283,n21113,n27251,n27252,n27184);
  nand U28862(n27184,G59428,n21080,n22386);
  nand U28863(n27252,G59428,n25365,n22165);
  not U28864(n22165,n21562);
  nand U28865(n27251,G59428,n27335);
  nand U28866(n27335,n27336,n27337,n25501,n27338);
  nor U28867(n27338,n27339,n27340,n27341);
  nor U28868(n27341,n21058,n27342);
  nor U28869(n27342,n27343,n27344,n27345);
  nor U28870(n27345,n26863,n27085,n27228);
  nor U28871(n27344,n26995,n21687);
  nor U28872(n27343,n21057,n21934);
  nor U28873(n27340,n27346,n26992);
  not U28874(n26992,n21933);
  nor U28875(n21933,n21846,n21849);
  nor U28876(n27346,n27347,n26994);
  nor U28877(n27347,n27228,n21069);
  nor U28878(n27339,n27348,n27349);
  and U28879(n25501,n27350,n27351,n27352,n27353);
  nor U28880(n27353,n27084,n27354,n27088);
  nor U28881(n27088,n21057,n25148);
  not U28882(n25148,n25367);
  and U28883(n27354,n21849,n27303);
  nor U28884(n27084,n21688,n24879);
  not U28885(n27352,n27227);
  nand U28886(n27227,n27355,n27356);
  nand U28887(n27356,n27357,n26863);
  nand U28888(n27357,n27082,n27078);
  nand U28889(n27078,n25522,n21534);
  not U28890(n27082,n26994);
  nand U28891(n27355,n25522,n21687,n26995);
  nand U28892(n27351,n21934,n21534,n26995);
  nand U28893(n27350,n27358,n27359);
  nand U28894(n27359,n25516,n21688,n27360,n21069);
  nand U28895(n27358,n27361,n26895);
  nand U28896(n27361,n27327,n25516);
  not U28897(n27327,n27360);
  nand U28898(n27337,n27362,n22473);
  nand U28899(n27336,n27130,n25368);
  not U28900(n21113,n22567);
  nor U28901(n22567,n27025,n21531);
  nor U28902(n27330,n26221,n26919);
  not U28903(n26221,n26069);
  xor U28904(n26069,n27363,n27364);
  xnor U28905(n27363,n27316,n27365);
  nor U28906(n27328,n27366,n27367,n27368,n27369);
  nor U28907(n27369,n27370,n25533);
  nor U28908(n27368,n27035,n21047);
  not U28909(n21047,n21075);
  nor U28910(n21075,G59427,G59426);
  and U28911(n27367,n22437,G59695);
  nor U28912(n22437,n25490,n21531);
  nand U28913(n25490,n25366,n21058,n27371);
  nor U28914(n27366,n22508,n25226);
  not U28915(n22508,n22436);
  nand U28916(n22436,n21943,n27372);
  nand U28917(n27372,G59428,n27373);
  nand U28918(n27373,n27374,n27375,n25494,n27246);
  nand U28919(n27246,n21548,n26995,n27085,n27376);
  nor U28920(n27376,n25522,n24879,n21687);
  nand U28921(n25494,n25522,n27377);
  nand U28922(n27377,n27378,n27360);
  nand U28923(n27360,n25366,n27379);
  nor U28924(n25366,n26863,n21057);
  nand U28925(n27378,n27379,n21548);
  nor U28926(n27379,n21846,n27085,n21934);
  nand U28927(n27375,n27257,n25365,n27130);
  nand U28928(n27374,n21031,n22386);
  nor U28929(n22386,n27132,n27380);
  not U28930(n27132,n27362);
  nor U28931(n27362,n25487,n21849,n27228,n27085);
  nand U28932(n21943,n20987,G59428);
  nor U28933(n20987,n21561,n21057);
  nand U28934(n22497,n22383,n21114);
  not U28935(n21114,n21691);
  nand U28936(n27238,G59760,n21108);
  nand U28937(n25492,n27185,n25237,n26994,n21846);
  nor U28938(n26994,n21534,n25522);
  nand U28939(n27237,G59601,n23278);
  nand U28940(n23278,n25533,n26919);
  nand U28941(n26919,G59797,G59427);
  not U28942(n25533,n21046);
  nand U28943(n27114,n26070,n27050);
  not U28944(n27050,n27023);
  nor U28945(n27023,n22049,n21692);
  not U28946(n21692,n27254);
  nand U28947(n27254,n25237,n21846,n27371);
  nor U28948(n27371,n26895,n21934,n25522,n27228);
  not U28949(n21934,n25368);
  nor U28950(n25368,n21687,n21849);
  nor U28951(n22049,n21561,n22163);
  nand U28952(n26070,n27381,n27382);
  nand U28953(n27382,n27383,n27384);
  nand U28954(n27383,n27276,n27385);
  nand U28955(n27385,n27277,n27275);
  nand U28956(n27381,n27386,n27387);
  nand U28957(n27387,n27277,n27388);
  nand U28958(n27388,n21061,n27276);
  or U28959(n27276,n27280,n27279);
  nand U28960(n27277,n27279,n27280);
  nand U28961(n27280,n27389,n27390);
  nand U28962(n27390,G59559,n27319);
  nand U28963(n27389,n21005,n21044);
  nand U28964(n27279,n27391,n27392);
  nand U28965(n27392,n27393,n27394);
  or U28966(n27394,n27364,n27316);
  not U28967(n27393,n27365);
  nand U28968(n27391,n27364,n27316);
  nand U28969(n27316,n27395,n27396);
  nand U28970(n27396,n21073,n27319,G59561);
  nand U28971(n21073,n21058,G59426);
  nand U28972(n27395,n21086,n21044);
  nand U28973(n27364,n27397,n27398);
  nand U28974(n27398,G59560,n27319);
  nand U28975(n27397,n21014,n21044);
  not U28976(n27386,n27384);
  nand U28977(n27384,n27399,n27400);
  nand U28978(n27400,G59558,n27319);
  nand U28979(n27319,n27365,n27275,n27401);
  nand U28980(n27401,G59426,n21846);
  not U28981(n27275,n21061);
  nor U28982(n21061,n21057,n21044);
  nand U28983(n27365,G59426,n27402);
  nand U28984(n27402,n27380,n27403);
  nand U28985(n27403,n27130,n25365);
  nand U28986(n25365,n27404,n27405);
  nand U28987(n27405,G59390,n21097);
  nor U28988(n27130,n21846,n22163);
  not U28989(n27380,n27348);
  nor U28990(n27348,n21688,n21058);
  nand U28991(n27399,n25535,n21044);
  nand U28992(n27113,n25354,n23116);
  nand U28993(n23116,n27406,n27407);
  nand U28994(n27407,n27126,n27053,n27063);
  not U28995(n27126,n27408);
  nand U28996(n27406,n27409,n24998);
  nand U28997(n27409,n27408,n27063);
  nand U28998(n27063,n21058,n24361);
  not U28999(n25354,n27025);
  nand U29000(n26952,n21031,n27410);
  nand U29001(n27410,n21562,n21561,n27411);
  not U29002(n27411,n27049);
  nand U29003(n27049,n25491,n27025);
  nand U29004(n27025,n22473,n27303,n27412);
  nor U29005(n27412,n21069,n25516,n21849);
  not U29006(n21069,n27110);
  nor U29007(n27303,n21534,n27085);
  nand U29008(n25491,n21539,n27185,n25367,n26863);
  nand U29009(n21561,n21058,n26895,n27257);
  nor U29010(n27257,n25487,n21687,n24879,n27228);
  not U29011(n25487,n27087);
  nor U29012(n27087,n25522,n26995);
  nand U29013(n21562,n25516,n21846,n26995,n27413);
  and U29014(n27413,n27185,n21548);
  nor U29015(n21548,n21534,n21057);
  nor U29016(n27185,n21688,n27085,n21849);
  not U29017(n27085,n26895);
  nand U29018(n26895,n27414,n27415,n27416,n27417);
  nor U29019(n27417,n27418,n27419,n27420,n27421);
  nor U29020(n27421,n27422,n22561);
  nor U29021(n27420,n27423,n22559);
  nor U29022(n27419,n27424,n22553);
  nor U29023(n27418,n27425,n22549);
  nor U29024(n27416,n27426,n27427,n27428,n27429);
  nor U29025(n27429,n27430,n22547);
  nor U29026(n27428,n27431,n22541);
  nor U29027(n27427,n27432,n22537);
  nor U29028(n27426,n27433,n22535);
  nor U29029(n27415,n27434,n27435,n27436,n27437);
  nor U29030(n27437,n27438,n22529);
  nor U29031(n27436,n27439,n22525);
  nor U29032(n27435,n27440,n22523);
  nor U29033(n27434,n27441,n22565);
  nor U29034(n27414,n27442,n27443,n27444,n27445);
  nor U29035(n27445,n27446,n22563);
  nor U29036(n27444,n27447,n22551);
  nor U29037(n27443,n27448,n22539);
  nor U29038(n27442,n27449,n22527);
  not U29039(n25516,n25522);
  nand U29040(n25522,n27450,n27451,n27452,n27453);
  nor U29041(n27453,n27454,n27455,n27456,n27457);
  nor U29042(n27457,n27422,n23417);
  not U29043(n23417,G59536);
  nor U29044(n27456,n27423,n23416);
  not U29045(n23416,G59528);
  nor U29046(n27455,n27424,n23427);
  not U29047(n23427,G59520);
  nor U29048(n27454,n27425,n23425);
  not U29049(n23425,G59504);
  nor U29050(n27452,n27458,n27459,n27460,n27461);
  nor U29051(n27461,n27430,n23424);
  not U29052(n23424,G59496);
  nor U29053(n27460,n27431,n22811);
  not U29054(n22811,G59488);
  nor U29055(n27459,n27432,n22809);
  not U29056(n22809,G59472);
  nor U29057(n27458,n27433,n22808);
  not U29058(n22808,G59464);
  nor U29059(n27451,n27462,n27463,n27464,n27465);
  nor U29060(n27465,n27438,n22803);
  not U29061(n22803,G59456);
  nor U29062(n27464,n27439,n22801);
  not U29063(n22801,G59440);
  nor U29064(n27463,n27440,n22800);
  not U29065(n22800,G59432);
  nor U29066(n27462,n27441,n23419);
  not U29067(n23419,G59552);
  nor U29068(n27450,n27466,n27467,n27468,n27469);
  nor U29069(n27469,n27446,n23418);
  not U29070(n23418,G59544);
  nor U29071(n27468,n27447,n23426);
  not U29072(n23426,G59512);
  nor U29073(n27467,n27448,n22810);
  not U29074(n22810,G59480);
  nor U29075(n27466,n27449,n22802);
  not U29076(n22802,G59448);
  not U29077(n21031,n21080);
  nand U29078(n21080,n27470,n27471);
  or U29079(n27471,n27472,n27473);
  nand U29080(n27470,n27474,n27472,n27475,n27476);
  nor U29081(n27476,n27477,n27478);
  nor U29082(n27478,n27479,n27096);
  nand U29083(n27096,n27480,n27481);
  nand U29084(n27481,G59562,n27482);
  nand U29085(n27482,G59557,n27483);
  or U29086(n27480,n27483,G59557);
  nor U29087(n27477,n24880,G59795,n26923);
  not U29088(n24880,G59557);
  nand U29089(n27475,n27484,n27485,n27486,n27487);
  nor U29090(n27487,n27488,n27489);
  nor U29091(n27489,n27479,n27099);
  xnor U29092(n27099,n27483,n27490);
  xnor U29093(n27490,n25536,G59557);
  not U29094(n25536,G59562);
  nand U29095(n27483,n27491,n27492);
  nand U29096(n27492,n27493,n26925);
  nand U29097(n27493,n27494,n24998);
  nand U29098(n27491,G59558,n27495);
  nor U29099(n27488,G59558,n27496);
  nand U29100(n27486,n27497,n27112);
  nand U29101(n27112,n27498,n27499);
  nand U29102(n27499,n27500,n27495);
  xnor U29103(n27500,G59563,G59558);
  nand U29104(n27498,n27501,n27494);
  not U29105(n27494,n27495);
  nand U29106(n27495,n27502,n27503);
  nand U29107(n27503,n27504,n26924);
  nand U29108(n27504,n27053,n27505);
  or U29109(n27502,n27505,n27053);
  xnor U29110(n27501,n26925,G59558);
  nand U29111(n27485,n27506,n27507);
  nand U29112(n27507,n27508,n27509);
  nand U29113(n27509,n27510,n27511);
  nand U29114(n27511,n21043,n27512,G59559);
  nand U29115(n27506,n27496,n27513);
  nand U29116(n27484,n27514,n27515,n27516);
  nand U29117(n27516,n27517,n27518);
  nand U29118(n27518,n27496,n27519);
  not U29119(n27517,n27520);
  nand U29120(n27515,n27513,n27508,n27496);
  nand U29121(n27508,n27497,n27105);
  xor U29122(n27105,n27521,n27505);
  nand U29123(n27505,n27522,n27523);
  nand U29124(n27523,G59565,n27524);
  or U29125(n27524,n27525,n24388);
  nand U29126(n27522,n27525,n24388);
  xnor U29127(n27521,G59564,G59559);
  nand U29128(n27514,n27526,n27527,n27528);
  nand U29129(n27528,n27510,n23142);
  nand U29130(n27527,n27529,n26923);
  nand U29131(n27529,n27530,n27513);
  nand U29132(n27513,n27349,n27531);
  nand U29133(n27531,n27228,n26863);
  nand U29134(n27530,n27519,n27520);
  nand U29135(n27520,n27532,n27533,n27534);
  nand U29136(n27534,n27497,n27111);
  xnor U29137(n27111,n27525,n27535);
  xnor U29138(n27535,n27035,G59560);
  not U29139(n27533,n27536);
  nand U29140(n27532,n27537,n27510);
  nand U29141(n27537,n27538,n27539,n21043);
  not U29142(n21043,G59425);
  nand U29143(n27539,n24388,n27512);
  not U29144(n27512,G59795);
  nand U29145(n27538,G59795,n27540);
  nand U29146(n27540,G59567,n21014);
  nand U29147(n27519,n27541,n27542);
  nand U29148(n27542,n27110,n27228);
  nor U29149(n27110,n21057,n26995);
  not U29150(n27541,n27473);
  nand U29151(n27526,n27497,n27109);
  nand U29152(n27109,n27525,n27543);
  nand U29153(n27543,G59566,n23142);
  nand U29154(n27525,G59561,n26606);
  not U29155(n27497,n27479);
  nand U29156(n27479,n27496,n27544);
  nand U29157(n27544,n27473,n27349);
  not U29158(n27349,n21539);
  nor U29159(n21539,n21534,n22163);
  nor U29160(n27473,n21688,n22163,n26995);
  not U29161(n26995,n26863);
  nand U29162(n27472,n27536,n24532);
  nand U29163(n24532,n27545,n27546,n27547,n27548);
  nor U29164(n27548,n27549,n27550,n27551,n27552);
  nor U29165(n27552,n22561,n24640);
  nand U29166(n24640,n27553,n27554);
  not U29167(n22561,G59533);
  nor U29168(n27551,n22559,n24641);
  nand U29169(n24641,n27553,n27555);
  not U29170(n22559,G59525);
  nor U29171(n27550,n22553,n24642);
  nand U29172(n24642,n27556,n27557);
  not U29173(n22553,G59517);
  nor U29174(n27549,n22549,n24643);
  nand U29175(n24643,n27557,n27554);
  not U29176(n22549,G59501);
  nor U29177(n27547,n27558,n27559,n27560,n27561);
  nor U29178(n27561,n22547,n24648);
  nand U29179(n24648,n27555,n27557);
  not U29180(n22547,G59493);
  nor U29181(n27560,n22541,n24649);
  nand U29182(n24649,n27562,n27556);
  not U29183(n22541,G59485);
  nor U29184(n27559,n22537,n24650);
  nand U29185(n24650,n27562,n27554);
  not U29186(n22537,G59469);
  nor U29187(n27558,n22535,n24651);
  nand U29188(n24651,n27562,n27555);
  not U29189(n22535,G59461);
  nor U29190(n27546,n27563,n27564,n27565,n27566);
  nor U29191(n27566,n22529,n24656);
  nand U29192(n24656,n27567,n27556);
  not U29193(n22529,G59453);
  nor U29194(n27565,n22525,n24657);
  nand U29195(n24657,n27567,n27554);
  nor U29196(n27554,n27370,n21086);
  not U29197(n22525,G59437);
  nor U29198(n27564,n22523,n24658);
  nand U29199(n24658,n27567,n27555);
  nor U29200(n27555,n21029,n27370);
  not U29201(n27370,n21014);
  not U29202(n22523,G59429);
  nor U29203(n27563,n22565,n24659);
  nand U29204(n24659,n27553,n27556);
  nor U29205(n27556,n21014,n21086);
  not U29206(n21086,n21029);
  not U29207(n22565,G59549);
  nor U29208(n27545,n27568,n27569,n27570,n27571);
  nor U29209(n27571,n22563,n24664);
  nand U29210(n24664,n27572,n27553);
  nor U29211(n27553,n21005,n25535);
  not U29212(n22563,G59541);
  nor U29213(n27570,n22551,n24665);
  nand U29214(n24665,n27572,n27557);
  nor U29215(n27557,n27062,n25535);
  not U29216(n25535,n27142);
  not U29217(n22551,G59509);
  nor U29218(n27569,n22539,n24666);
  nand U29219(n24666,n27572,n27562);
  nor U29220(n27562,n27142,n21005);
  not U29221(n22539,G59477);
  nor U29222(n27568,n22527,n24667);
  nand U29223(n24667,n27572,n27567);
  nor U29224(n27567,n27142,n27062);
  not U29225(n27062,n21005);
  xor U29226(n21005,n27573,n27574);
  xnor U29227(n27142,n27575,n27576);
  nor U29228(n27576,n27573,n27574);
  and U29229(n27574,n27577,n27578);
  nand U29230(n27578,n27579,n27580);
  or U29231(n27580,n27581,n27582);
  not U29232(n27579,n27583);
  nand U29233(n27577,n27582,n27581);
  and U29234(n27573,n27584,n27585,n27586);
  nand U29235(n27586,G59564,n21046);
  nand U29236(n27585,n25913,n21044);
  xnor U29237(n25913,n25915,n26924);
  nand U29238(n27584,n22385,G59559);
  nand U29239(n27575,n27587,n27588,n27589);
  nand U29240(n27589,n21044,n25912);
  not U29241(n25912,n26526);
  nor U29242(n26526,n26213,n26296,n27590);
  nor U29243(n27590,n26925,n25915);
  nor U29244(n26296,n26925,G59564);
  not U29245(n26925,G59563);
  not U29246(n26213,n26153);
  nand U29247(n26153,n25915,n25990);
  nor U29248(n25990,n26924,G59563);
  not U29249(n26924,G59564);
  nor U29250(n25915,n26606,n27035);
  nand U29251(n27588,G59563,n21046);
  nand U29252(n27587,n22385,G59558);
  nor U29253(n27572,n21029,n21014);
  xor U29254(n21014,n27591,n27582);
  nand U29255(n27582,n27592,n27593);
  nand U29256(n27593,n26935,n27594);
  xnor U29257(n27594,n25226,n27595);
  nor U29258(n27595,n21544,n25224);
  nand U29259(n21544,n27596,n27597);
  nand U29260(n27597,G59427,n22397);
  not U29261(n22397,G59598);
  or U29262(n27596,G59427,G59757);
  not U29263(n25226,G59568);
  nand U29264(n27592,n25237,n22385);
  xnor U29265(n27591,n27583,n27581);
  nand U29266(n27581,n27598,n27599,n27600);
  nand U29267(n27600,G59565,n21046);
  nand U29268(n27599,n26605,n21044);
  not U29269(n26605,n26758);
  nor U29270(n26758,n25834,n25759);
  nor U29271(n25759,n26606,G59565);
  nor U29272(n25834,n27035,G59566);
  not U29273(n27035,G59565);
  nand U29274(n27598,n22385,G59560);
  nand U29275(n21029,n27601,n27583);
  nand U29276(n27583,n27602,n27603);
  or U29277(n27601,n27603,n27602);
  nand U29278(n27602,n27604,n27605,G59426);
  nand U29279(n27605,n26923,n21070);
  nand U29280(n21070,n24879,n21846,n25237);
  nor U29281(n25237,n26863,n22163);
  not U29282(n22163,n21057);
  nand U29283(n21057,n27606,n27607,n27608,n27609);
  nor U29284(n27609,n27610,n27611,n27612,n27613);
  nor U29285(n27613,n27422,n23048);
  not U29286(n23048,G59539);
  nor U29287(n27612,n27423,n23047);
  not U29288(n23047,G59531);
  nor U29289(n27611,n27424,n23042);
  not U29290(n23042,G59523);
  nor U29291(n27610,n27425,n23040);
  not U29292(n23040,G59507);
  nor U29293(n27608,n27614,n27615,n27616,n27617);
  nor U29294(n27617,n27430,n23039);
  not U29295(n23039,G59499);
  nor U29296(n27616,n27431,n23034);
  not U29297(n23034,G59491);
  nor U29298(n27615,n27432,n23032);
  not U29299(n23032,G59475);
  nor U29300(n27614,n27433,n23031);
  not U29301(n23031,G59467);
  nor U29302(n27607,n27618,n27619,n27620,n27621);
  nor U29303(n27621,n27438,n23026);
  not U29304(n23026,G59459);
  nor U29305(n27620,n27439,n23024);
  not U29306(n23024,G59443);
  nor U29307(n27619,n27440,n23023);
  not U29308(n23023,G59435);
  nor U29309(n27618,n27441,n23050);
  not U29310(n23050,G59555);
  nor U29311(n27606,n27622,n27623,n27624,n27625);
  nor U29312(n27625,n27446,n23049);
  not U29313(n23049,G59547);
  nor U29314(n27624,n27447,n23041);
  not U29315(n23041,G59515);
  nor U29316(n27623,n27448,n23033);
  not U29317(n23033,G59483);
  nor U29318(n27622,n27449,n23025);
  not U29319(n23025,G59451);
  nand U29320(n26863,n27626,n27627,n27628,n27629);
  nor U29321(n27629,n27630,n27631,n27632,n27633);
  nor U29322(n27633,n27422,n23336);
  not U29323(n23336,G59535);
  nor U29324(n27632,n27423,n23335);
  not U29325(n23335,G59527);
  nor U29326(n27631,n27424,n23346);
  not U29327(n23346,G59519);
  nor U29328(n27630,n27425,n23344);
  not U29329(n23344,G59503);
  nor U29330(n27628,n27634,n27635,n27636,n27637);
  nor U29331(n27637,n27430,n23343);
  not U29332(n23343,G59495);
  nor U29333(n27636,n27431,n22730);
  not U29334(n22730,G59487);
  nor U29335(n27635,n27432,n22728);
  not U29336(n22728,G59471);
  nor U29337(n27634,n27433,n22727);
  not U29338(n22727,G59463);
  nor U29339(n27627,n27638,n27639,n27640,n27641);
  nor U29340(n27641,n27438,n22722);
  not U29341(n22722,G59455);
  nor U29342(n27640,n27439,n22720);
  not U29343(n22720,G59439);
  nor U29344(n27639,n27440,n22719);
  not U29345(n22719,G59431);
  nor U29346(n27638,n27441,n23338);
  not U29347(n23338,G59551);
  nor U29348(n27626,n27642,n27643,n27644,n27645);
  nor U29349(n27645,n27446,n23337);
  not U29350(n23337,G59543);
  nor U29351(n27644,n27447,n23345);
  not U29352(n23345,G59511);
  nor U29353(n27643,n27448,n22729);
  not U29354(n22729,G59479);
  nor U29355(n27642,n27449,n22721);
  not U29356(n22721,G59447);
  nor U29357(n27649,n27650,n27651,n27652,n27653);
  nor U29358(n27653,n27422,n23144);
  not U29359(n23144,G59540);
  nor U29360(n27652,n27423,n23140);
  not U29361(n23140,G59532);
  nor U29362(n27651,n27424,n23135);
  not U29363(n23135,G59524);
  nor U29364(n27650,n27425,n23133);
  not U29365(n23133,G59508);
  nor U29366(n27648,n27654,n27655,n27656,n27657);
  nor U29367(n27657,n27430,n23131);
  not U29368(n23131,G59500);
  nor U29369(n27656,n27431,n23125);
  not U29370(n23125,G59492);
  nor U29371(n27655,n27432,n23123);
  not U29372(n23123,G59476);
  nor U29373(n27654,n27433,n23121);
  not U29374(n23121,G59468);
  nor U29375(n27647,n27658,n27659,n27660,n27661);
  nor U29376(n27661,n27438,n23113);
  not U29377(n23113,G59460);
  nor U29378(n27660,n27439,n23109);
  not U29379(n23109,G59444);
  nor U29380(n27659,n27440,n23106);
  not U29381(n23106,G59436);
  nor U29382(n27658,n27441,n23147);
  not U29383(n23147,G59556);
  nor U29384(n27646,n27662,n27663,n27664,n27665);
  nor U29385(n27665,n27446,n23145);
  not U29386(n23145,G59548);
  nor U29387(n27664,n27447,n23134);
  not U29388(n23134,G59516);
  nor U29389(n27663,n27448,n23124);
  not U29390(n23124,G59484);
  nor U29391(n27662,n27449,n23111);
  not U29392(n23111,G59452);
  not U29393(n24879,n21849);
  nand U29394(n21849,n27666,n27667,n27668,n27669);
  nor U29395(n27669,n27670,n27671,n27672,n27673);
  nor U29396(n27673,n27422,n23586);
  not U29397(n23586,G59538);
  nor U29398(n27672,n27423,n23585);
  not U29399(n23585,G59530);
  nor U29400(n27671,n27424,n23596);
  not U29401(n23596,G59522);
  nor U29402(n27670,n27425,n23594);
  not U29403(n23594,G59506);
  nor U29404(n27668,n27674,n27675,n27676,n27677);
  nor U29405(n27677,n27430,n23593);
  not U29406(n23593,G59498);
  nor U29407(n27676,n27431,n22964);
  not U29408(n22964,G59490);
  nor U29409(n27675,n27432,n22962);
  not U29410(n22962,G59474);
  nor U29411(n27674,n27433,n22961);
  not U29412(n22961,G59466);
  nor U29413(n27667,n27678,n27679,n27680,n27681);
  nor U29414(n27681,n27438,n22956);
  not U29415(n22956,G59458);
  nor U29416(n27680,n27439,n22954);
  not U29417(n22954,G59442);
  nor U29418(n27679,n27440,n22953);
  not U29419(n22953,G59434);
  nor U29420(n27678,n27441,n23588);
  not U29421(n23588,G59554);
  nor U29422(n27666,n27682,n27683,n27684,n27685);
  nor U29423(n27685,n27446,n23587);
  not U29424(n23587,G59546);
  nor U29425(n27684,n27447,n23595);
  not U29426(n23595,G59514);
  nor U29427(n27683,n27448,n22963);
  not U29428(n22963,G59482);
  nor U29429(n27682,n27449,n22955);
  not U29430(n22955,G59450);
  nand U29431(n27604,n21560,n27686);
  nand U29432(n27686,G59428,n25224);
  not U29433(n25224,G59567);
  not U29434(n21560,n22385);
  nand U29435(n27603,n22384,n27687,n27688,n27689);
  nand U29436(n27689,n21044,n26606);
  not U29437(n26606,G59566);
  nand U29438(n27688,G59566,n21046);
  nor U29439(n21046,n21044,G59428);
  nand U29440(n27687,n22385,G59561);
  nor U29441(n22385,n21531,G59427);
  not U29442(n22527,G59445);
  nor U29443(n27536,n21688,n27228,n27510);
  not U29444(n27510,n27496);
  nor U29445(n27496,G59427,G59425);
  not U29446(n27228,n21534);
  nand U29447(n21534,n27690,n27691,n27692,n27693);
  nor U29448(n27693,n27694,n27695,n27696,n27697);
  nor U29449(n27697,n27422,n23256);
  not U29450(n23256,G59534);
  nor U29451(n27696,n27423,n23255);
  not U29452(n23255,G59526);
  nor U29453(n27695,n27424,n23266);
  not U29454(n23266,G59518);
  nor U29455(n27694,n27425,n23264);
  not U29456(n23264,G59502);
  nor U29457(n27692,n27698,n27699,n27700,n27701);
  nor U29458(n27701,n27430,n23263);
  not U29459(n23263,G59494);
  nor U29460(n27700,n27431,n22654);
  not U29461(n22654,G59486);
  nor U29462(n27699,n27432,n22652);
  not U29463(n22652,G59470);
  nor U29464(n27698,n27433,n22651);
  not U29465(n22651,G59462);
  nor U29466(n27691,n27702,n27703,n27704,n27705);
  nor U29467(n27705,n27438,n22646);
  not U29468(n22646,G59454);
  nor U29469(n27704,n27439,n22644);
  not U29470(n22644,G59438);
  nor U29471(n27703,n27440,n22643);
  not U29472(n22643,G59430);
  nor U29473(n27702,n27441,n23258);
  not U29474(n23258,G59550);
  nor U29475(n27690,n27706,n27707,n27708,n27709);
  nor U29476(n27709,n27446,n23257);
  not U29477(n23257,G59542);
  nor U29478(n27708,n27447,n23265);
  not U29479(n23265,G59510);
  nor U29480(n27707,n27448,n22653);
  not U29481(n22653,G59478);
  nor U29482(n27706,n27449,n22645);
  not U29483(n22645,G59446);
  not U29484(n21688,n21687);
  nand U29485(n21687,n27710,n27711,n27712,n27713);
  nor U29486(n27713,n27714,n27715,n27716,n27717);
  nor U29487(n27717,n27422,n23501);
  not U29488(n23501,G59537);
  nand U29489(n27422,n27408,n24362);
  nor U29490(n27716,n27423,n23500);
  not U29491(n23500,G59529);
  nand U29492(n27423,n24361,n27408);
  nor U29493(n27715,n27424,n23511);
  not U29494(n23511,G59521);
  nand U29495(n27424,n24370,n24389);
  nor U29496(n27714,n27425,n23509);
  not U29497(n23509,G59505);
  nand U29498(n27425,n24389,n24362);
  nor U29499(n27712,n27718,n27719,n27720,n27721);
  nor U29500(n27721,n27430,n23508);
  not U29501(n23508,G59497);
  nand U29502(n27430,n24361,n24389);
  nor U29503(n27720,n27431,n22885);
  not U29504(n22885,G59489);
  nand U29505(n27431,n24387,n24370);
  nor U29506(n27719,n27432,n22883);
  not U29507(n22883,G59473);
  nand U29508(n27432,n24387,n24362);
  nor U29509(n27718,n27433,n22882);
  not U29510(n22882,G59465);
  nand U29511(n27433,n24387,n24361);
  nor U29512(n27711,n27722,n27723,n27724,n27725);
  nor U29513(n27725,n27438,n22877);
  not U29514(n22877,G59457);
  nand U29515(n27438,n27123,n24370);
  nor U29516(n27724,n27439,n22875);
  not U29517(n22875,G59441);
  nand U29518(n27439,n27123,n24362);
  nor U29519(n24362,n24388,G59561);
  nor U29520(n27723,n27440,n22874);
  not U29521(n22874,G59433);
  nand U29522(n27440,n27123,n24361);
  nor U29523(n24361,n23142,n24388);
  not U29524(n24388,G59560);
  nor U29525(n27722,n27441,n23503);
  not U29526(n23503,G59553);
  nand U29527(n27441,n27408,n24370);
  nor U29528(n24370,G59560,G59561);
  nor U29529(n27710,n27726,n27727,n27728,n27729);
  nor U29530(n27729,n27446,n23502);
  not U29531(n23502,G59545);
  nand U29532(n27446,n24369,n27408);
  nor U29533(n27408,G59559,G59558);
  nor U29534(n27728,n27447,n23510);
  not U29535(n23510,G59513);
  nand U29536(n27447,n24369,n24389);
  nor U29537(n24389,n27053,G59558);
  nor U29538(n27727,n27448,n22884);
  not U29539(n22884,G59481);
  nand U29540(n27448,n24369,n24387);
  nor U29541(n24387,n24998,G59559);
  nor U29542(n27726,n27449,n22876);
  not U29543(n22876,G59449);
  nand U29544(n27449,n24369,n27123);
  nor U29545(n27123,n24998,n27053);
  not U29546(n27053,G59559);
  not U29547(n24998,G59558);
  nor U29548(n24369,n23142,G59560);
  not U29549(n23142,G59561);
  nand U29550(n27474,G59557,G59425);
  nand U29551(n21019,G59425,n21531);
  not U29552(n26945,n25539);
  nor U29553(n25539,n21531,n22384);
  not U29554(n22384,n26935);
  nor U29555(n26935,n26923,n21044);
  not U29556(n21044,G59426);
  not U29557(n26923,G59427);
  not U29558(n21531,G59428);
  nor U29559(G8373,n20977,n21158);
  not U29560(n21158,G59424);
  nor U29561(G8372,n20977,n21157);
  not U29562(n21157,G59423);
  nor U29563(G8371,n20977,n21156);
  not U29564(n21156,G59422);
  nor U29565(G8370,n20977,n21155);
  not U29566(n21155,G59421);
  nor U29567(G8369,n20977,n21154);
  not U29568(n21154,G59420);
  nor U29569(G8368,n20977,n21153);
  not U29570(n21153,G59419);
  nor U29571(G8367,n20977,n21152);
  not U29572(n21152,G59418);
  nor U29573(G8366,n20977,n21151);
  not U29574(n21151,G59417);
  nor U29575(G8365,n20977,n21150);
  not U29576(n21150,G59416);
  nor U29577(G8364,n20977,n21149);
  not U29578(n21149,G59415);
  nor U29579(G8363,n20977,n21148);
  not U29580(n21148,G59414);
  nor U29581(G8362,n20977,n21147);
  not U29582(n21147,G59413);
  nor U29583(G8361,n20977,n21146);
  not U29584(n21146,G59412);
  nor U29585(G8360,n20977,n21145);
  not U29586(n21145,G59411);
  nor U29587(G8359,n20977,n21144);
  not U29588(n21144,G59410);
  nor U29589(G8358,n20977,n21143);
  not U29590(n21143,G59409);
  and U29591(G8357,n20978,G59408);
  and U29592(G8356,n20978,G59407);
  and U29593(G8355,n20978,G59406);
  and U29594(G8354,n20978,G59405);
  and U29595(G8353,n20978,G59404);
  and U29596(G8352,n20978,G59403);
  and U29597(G8351,n20978,G59402);
  and U29598(G8350,n20978,G59401);
  nor U29599(G8349,n20977,n21164);
  not U29600(n21164,G59400);
  nor U29601(G8348,n20977,n21163);
  not U29602(n21163,G59399);
  nor U29603(G8347,n20977,n21162);
  not U29604(n21162,G59398);
  nor U29605(G8346,n20977,n21161);
  not U29606(n21161,G59397);
  and U29607(G8345,n20978,G59396);
  and U29608(G8344,n20978,G59395);
  not U29609(n20978,n20977);
  nand U29610(n20977,n27730,n27731);
  nand U29611(n27731,G59392,n27732);
  nand U29612(G8343,n27733,n27734,n27735,n27736);
  nor U29613(n27736,n27737,n20982,n27738);
  nor U29614(n27738,n27404,n21045);
  not U29615(n27404,n27732);
  nor U29616(n20982,G59392,G59390);
  nor U29617(n27737,n27730,n27739);
  nand U29618(n27735,n20965,n21037);
  nand U29619(n27734,n27740,n21097);
  nand U29620(n27733,G33,G59392,G59391);
  nand U29621(G8342,n27741,n27742,n27743,n27744);
  nand U29622(n27744,G33,n27732);
  nor U29623(n27732,n21097,G59390);
  nor U29624(n27743,n27745,n27746);
  nor U29625(n27746,n21037,n27740,n22050);
  nor U29626(n27740,n27747,n27748);
  or U29627(n27742,n27730,n27748);
  nand U29628(n27730,n21097,n22050);
  nand U29629(n27741,n21944,G59391);
  nand U29630(G8341,n27749,n27750,n27751,n27752);
  nand U29631(n27752,G59390,n27739,n22050);
  not U29632(n22050,G59392);
  nand U29633(n27751,G33,n27753,G59392);
  nand U29634(n27753,n27748,n27754);
  nand U29635(n27754,n21097,n21037);
  not U29636(n27750,n27755);
  nand U29637(n27749,G59391,n27756,n21944);
  not U29638(n21944,n21045);
  nand U29639(n21045,G58904,G58903);
  nand U29640(n27756,n27748,n27757);
  nand U29641(n27757,n27758,n27739,G59392);
  nand U29642(n27758,n21037,n27747);
  not U29643(n21037,G59798);
  nand U29644(G8340,n27759,n27760,n27761);
  nand U29645(n27761,G59389,n20965);
  nand U29646(n27760,n27755,G59759);
  nand U29647(n27759,n27745,G59760);
  nand U29648(G8339,n27762,n27763,n27764);
  nand U29649(n27764,G59388,n20965);
  nand U29650(n27763,n27755,G59760);
  nand U29651(n27762,n27745,G59761);
  nand U29652(G8338,n27765,n27766,n27767);
  nand U29653(n27767,G59387,n20965);
  nand U29654(n27766,n27755,G59761);
  nand U29655(n27765,n27745,G59762);
  nand U29656(G8337,n27768,n27769,n27770);
  nand U29657(n27770,G59386,n20965);
  nand U29658(n27769,n27755,G59762);
  nand U29659(n27768,n27745,G59763);
  nand U29660(G8336,n27771,n27772,n27773);
  nand U29661(n27773,G59385,n20965);
  nand U29662(n27772,n27755,G59763);
  nand U29663(n27771,n27745,G59764);
  nand U29664(G8335,n27774,n27775,n27776);
  nand U29665(n27776,G59384,n20965);
  nand U29666(n27775,n27755,G59764);
  nand U29667(n27774,n27745,G59765);
  nand U29668(G8334,n27777,n27778,n27779);
  nand U29669(n27779,G59383,n20965);
  nand U29670(n27778,n27755,G59765);
  nand U29671(n27777,n27745,G59766);
  nand U29672(G8333,n27780,n27781,n27782);
  nand U29673(n27782,G59382,n20965);
  nand U29674(n27781,n27755,G59766);
  nand U29675(n27780,n27745,G59767);
  nand U29676(G8332,n27783,n27784,n27785);
  nand U29677(n27785,G59381,n20965);
  nand U29678(n27784,n27755,G59767);
  nand U29679(n27783,n27745,G59768);
  nand U29680(G8331,n27786,n27787,n27788);
  nand U29681(n27788,G59380,n20965);
  nand U29682(n27787,n27755,G59768);
  nand U29683(n27786,n27745,G59769);
  nand U29684(G8330,n27789,n27790,n27791);
  nand U29685(n27791,G59379,n20965);
  nand U29686(n27790,n27755,G59769);
  nand U29687(n27789,n27745,G59770);
  nand U29688(G8329,n27792,n27793,n27794);
  nand U29689(n27794,G59378,n20965);
  nand U29690(n27793,n27755,G59770);
  nand U29691(n27792,n27745,G59771);
  nand U29692(G8328,n27795,n27796,n27797);
  nand U29693(n27797,G59377,n20965);
  nand U29694(n27796,n27755,G59771);
  nand U29695(n27795,n27745,G59772);
  nand U29696(G8327,n27798,n27799,n27800);
  nand U29697(n27800,G59376,n20965);
  nand U29698(n27799,n27755,G59772);
  nand U29699(n27798,n27745,G59773);
  nand U29700(G8326,n27801,n27802,n27803);
  nand U29701(n27803,G59375,n20965);
  nand U29702(n27802,n27755,G59773);
  nand U29703(n27801,n27745,G59774);
  nand U29704(G8325,n27804,n27805,n27806);
  nand U29705(n27806,G59374,n20965);
  nand U29706(n27805,n27755,G59774);
  nand U29707(n27804,n27745,G59775);
  nand U29708(G8324,n27807,n27808,n27809);
  nand U29709(n27809,G59373,n20965);
  nand U29710(n27808,n27755,G59775);
  nand U29711(n27807,n27745,G59776);
  nand U29712(G8323,n27810,n27811,n27812);
  nand U29713(n27812,G59372,n20965);
  nand U29714(n27811,n27755,G59776);
  nand U29715(n27810,n27745,G59777);
  nand U29716(G8322,n27813,n27814,n27815);
  nand U29717(n27815,G59371,n20965);
  nand U29718(n27814,n27755,G59777);
  nand U29719(n27813,n27745,G59778);
  nand U29720(G8321,n27816,n27817,n27818);
  nand U29721(n27818,G59370,n20965);
  nand U29722(n27817,n27755,G59778);
  nand U29723(n27816,n27745,G59779);
  nand U29724(G8320,n27819,n27820,n27821);
  nand U29725(n27821,G59369,n20965);
  nand U29726(n27820,n27755,G59779);
  nand U29727(n27819,n27745,G59780);
  nand U29728(G8319,n27822,n27823,n27824);
  nand U29729(n27824,G59368,n20965);
  nand U29730(n27823,n27755,G59780);
  nand U29731(n27822,n27745,G59781);
  nand U29732(G8318,n27825,n27826,n27827);
  nand U29733(n27827,G59367,n20965);
  nand U29734(n27826,n27755,G59781);
  nand U29735(n27825,n27745,G59782);
  nand U29736(G8317,n27828,n27829,n27830);
  nand U29737(n27830,G59366,n20965);
  nand U29738(n27829,n27755,G59782);
  nand U29739(n27828,n27745,G59783);
  nand U29740(G8316,n27831,n27832,n27833);
  nand U29741(n27833,G59365,n20965);
  nand U29742(n27832,n27755,G59783);
  nand U29743(n27831,n27745,G59784);
  nand U29744(G8315,n27834,n27835,n27836);
  nand U29745(n27836,G59364,n20965);
  nand U29746(n27835,n27755,G59784);
  nand U29747(n27834,n27745,G59785);
  nand U29748(G8314,n27837,n27838,n27839);
  nand U29749(n27839,G59363,n20965);
  nand U29750(n27838,n27755,G59785);
  nand U29751(n27837,n27745,G59786);
  nand U29752(G8313,n27840,n27841,n27842);
  nand U29753(n27842,G59362,n20965);
  nand U29754(n27841,n27755,G59786);
  nand U29755(n27840,n27745,G59787);
  nand U29756(G8312,n27843,n27844,n27845);
  nand U29757(n27845,G59361,n20965);
  nand U29758(n27844,n27755,G59787);
  nand U29759(n27843,n27745,G59788);
  nand U29760(G8311,n27846,n27847,n27848);
  nand U29761(n27848,G59360,n20965);
  nand U29762(n27847,n27755,G59788);
  not U29763(n27748,G59390);
  nand U29764(n27846,n27745,G59789);
  nor U29765(n20966,n21097,G59392);
  not U29766(n21097,G59391);
  nand U29767(G3276,n27849,n27850);
  nand U29768(n27850,G58907,n27851);
  nand U29769(n27849,G59341,n27852);
  nand U29770(G3275,n27853,n27854);
  nand U29771(n27854,G58908,n27851);
  nand U29772(n27853,G59342,n27852);
  nand U29773(G3274,n27855,n27856);
  nand U29774(n27856,G58909,n27851);
  nand U29775(n27855,G59343,n27852);
  nand U29776(G3273,n27857,n27858);
  nand U29777(n27858,G58910,n27851);
  nand U29778(n27857,G59344,n27852);
  nand U29779(G3272,n27859,n27860);
  nand U29780(n27860,n27861,n20976,n27862);
  nand U29781(n27859,G58944,n27863);
  nand U29782(G3271,n27864,n27865);
  nand U29783(n27865,G58945,n27863);
  nand U29784(n27864,n27866,n27862);
  nand U29785(n27866,n20976,n27861);
  not U29786(n27861,n27867);
  nand U29787(G3270,n27868,n27869);
  nand U29788(n27869,n27870,n27871,n27872,n27873);
  nand U29789(n27868,n27874,G59108);
  nand U29790(G3269,n27875,n27876);
  nand U29791(n27876,n27874,G59109);
  nand U29792(n27875,n27877,n27873);
  nand U29793(n27877,n27878,n27879);
  nand U29794(n27879,n27880,n27881);
  nand U29795(n27878,n27870,n27882);
  nand U29796(G3268,n27883,n27884);
  nand U29797(n27884,n27874,G59110);
  nand U29798(n27883,n27885,n27873);
  nand U29799(n27885,n27886,n27887,n27888);
  nand U29800(n27888,n27870,n27889);
  nand U29801(n27887,G58978,n27890,G59118);
  nand U29802(n27886,n27891,n27880);
  nand U29803(G3266,n27892,n27893);
  nand U29804(n27893,n27874,G59111);
  nand U29805(n27892,n27894,n27873);
  nand U29806(n27894,n27895,n27896,n27897);
  nand U29807(n27897,n27870,n27898);
  nand U29808(n27896,G58978,n27899,G59118);
  nand U29809(n27895,n27900,n27880);
  nand U29810(G3265,n27901,n27902);
  nand U29811(n27902,n27874,G59112);
  not U29812(n27874,n27873);
  nand U29813(n27901,n27903,n27873);
  nand U29814(n27873,n27904,n27905,n27906);
  nand U29815(n27906,n27907,n27908);
  nand U29816(n27903,n27909,n27910,n27911);
  nand U29817(n27911,n27870,n27912);
  nand U29818(n27910,G58978,n27913);
  nand U29819(n27913,G59118,n27914);
  nand U29820(n27909,n27880,n27915);
  nor U29821(n27880,n27916,G58977);
  nand U29822(G3264,n27917,n27918);
  or U29823(n27918,n27851,G59354);
  nand U29824(n27917,G59345,n27851);
  nand U29825(G3263,n27919,n27920);
  or U29826(n27920,n27921,n27922);
  nand U29827(n27919,n27923,n27921);
  nand U29828(n27921,n27924,n27925,n27926,n27927);
  nand U29829(n27926,n27928,n27929);
  nand U29830(n27925,G58978,n27930,n27931);
  nand U29831(n27923,n27932,n27933);
  nand U29832(n27933,G58979,n27934);
  nand U29833(n27934,n27935,n27930);
  nand U29834(n27935,n27936,n27937);
  nand U29835(n27937,G58977,n27938);
  nand U29836(n27938,n27939,n27940);
  nand U29837(n27940,n27941,n27942);
  nand U29838(n27941,n27943,n27944);
  nand U29839(n27939,G59348,n27945);
  nand U29840(n27936,n27946,n27943);
  nand U29841(G3262,n27947,n27948);
  nand U29842(n27948,G59351,n27851);
  nand U29843(n27947,G59355,n27852);
  nand U29844(G3261,n27949,n27950);
  nand U29845(n27950,n27951,G59354);
  nand U29846(n27949,n27952,n27953);
  nand U29847(n27952,n27954,n27955,G58977);
  nand U29848(G3260,n27956,n27957);
  nand U29849(n27957,n27951,G59355);
  not U29850(n27951,n27953);
  nand U29851(n27956,n27953,n27958);
  nand U29852(n27953,n27924,n27959);
  nand U29853(n27959,n27960,n27928);
  nand U29854(G2747,n27961,n27962,n27963,n27964);
  nand U29855(n27964,G58979,n27965,n27966);
  nand U29856(n27963,n27967,G59117);
  nand U29857(n27962,n27968,n27969);
  nand U29858(n27961,n27970,n27971);
  nand U29859(G2745,n27863,n27972);
  nand U29860(n27972,G59353,G58943);
  nand U29861(G2744,n27973,n27974);
  nand U29862(n27974,G58979,n27928,n27960);
  nand U29863(n27973,G59352,n27975);
  nand U29864(n27975,n27976,n27907);
  nand U29865(G2743,n27977,n27978,n27979);
  or U29866(n27978,n27851,G59352);
  nand U29867(n27977,G59350,n27851);
  nand U29868(G2742,n27980,n27981,n27979);
  nand U29869(n27979,n27867,n27982);
  nand U29870(n27981,G35,n27862);
  nand U29871(n27980,G59348,n27863);
  nand U29872(G2741,n27983,n27984);
  nand U29873(n27984,n27985,n27986);
  nand U29874(n27985,n27987,n27988);
  nand U29875(n27988,n27989,n27990);
  nand U29876(n27989,n27991,n27992);
  nand U29877(n27992,n27993,n27870);
  nand U29878(n27987,n27916,n27994);
  nand U29879(n27994,n27995,n27996);
  nand U29880(n27996,n27870,n27997);
  nand U29881(n27997,n27998,n27999);
  nand U29882(n27983,G59347,n28000);
  nand U29883(G2740,n28001,n28002);
  nand U29884(n28002,G59346,n28000);
  nand U29885(n28000,n27907,n27986);
  nand U29886(G2739,n28003,n28004,n28005);
  nand U29887(n28004,G59344,n28006);
  nand U29888(n28003,n28007,G59309);
  nand U29889(G2738,n28005,n28008,n28009);
  nand U29890(n28009,G59343,n28006);
  nand U29891(G2737,n28010,n28011,n28012);
  or U29892(n28012,n28005,n28013);
  nand U29893(n28005,n28007,G59310);
  nand U29894(n28011,G59342,n28006);
  nand U29895(n28010,n28014,n28015,n28016,n28007);
  nand U29896(n28016,G59309,G58944);
  nand U29897(G2736,n28017,n28018,n28008);
  nand U29898(n28008,n28007,n28019,n28014,n28013);
  nand U29899(n28018,G59341,n28006);
  nand U29900(n28017,n28014,n28015,n28007);
  not U29901(n28007,n28006);
  nand U29902(n28006,n28020,n28021,n28022,n28023);
  nor U29903(n28023,n28024,n28025,n28026,n28027);
  nand U29904(n28027,n28028,n28029,n28030,n28031);
  nand U29905(n28026,n28032,n28033,n28034,n28035);
  nand U29906(n28025,n28036,n28037,n28038,n28039);
  nand U29907(n28024,n28040,n28041,n28042,n28043);
  nor U29908(n28022,n28044,n28045,G58947,G58946);
  nor U29909(n28045,n28019,n28014);
  not U29910(n28019,G58944);
  nand U29911(n28044,n28046,n28047,n28048,n28049);
  nor U29912(n28021,G58959,G58958,G58957,G58956);
  nor U29913(n28020,G58955,G58954,G58953,G58952);
  not U29914(n28014,G58945);
  nand U29915(G2735,n28050,n28051,n28052,n28053);
  nor U29916(n28053,n28054,n28055,n28056);
  nor U29917(n28056,n28057,n28058);
  and U29918(n28055,n28059,n28060);
  nor U29919(n28054,n28061,n28062);
  nand U29920(n28052,n28063,n28064);
  nand U29921(n28051,n28065,n28066);
  nand U29922(n28050,n28067,G59308);
  nand U29923(G2734,n28068,n28069,n28070,n28071);
  nor U29924(n28071,n28072,n28073,n28074);
  nor U29925(n28074,n28075,n28058);
  nor U29926(n28073,n28076,n28077);
  nor U29927(n28072,n28078,n28062);
  nand U29928(n28070,n28079,n28064);
  nand U29929(n28069,n28065,n28080);
  nand U29930(n28068,n28067,G59307);
  nand U29931(G2733,n28081,n28082,n28083,n28084);
  nor U29932(n28084,n28085,n28086,n28087);
  nor U29933(n28087,n28088,n28058);
  nor U29934(n28086,n28076,n28089);
  nor U29935(n28085,n28090,n28062);
  nand U29936(n28083,n28091,n28064);
  nand U29937(n28082,n28092,n28065);
  nand U29938(n28081,n28067,G59306);
  nand U29939(G2732,n28093,n28094,n28095,n28096);
  nor U29940(n28096,n28097,n28098,n28099);
  nor U29941(n28099,n28100,n28058);
  nor U29942(n28098,n28076,n28101);
  nor U29943(n28097,n28102,n28062);
  nand U29944(n28095,n28103,n28064);
  nand U29945(n28094,n28065,n28104);
  nand U29946(n28093,n28067,G59305);
  nand U29947(G2731,n28105,n28106,n28107,n28108);
  nor U29948(n28108,n28109,n28110,n28111);
  nor U29949(n28111,n28112,n28058);
  nor U29950(n28110,n28076,n28113);
  nor U29951(n28109,n28114,n28062);
  nand U29952(n28107,n28115,n28064);
  nand U29953(n28106,n28065,n28116);
  nand U29954(n28105,n28067,G59304);
  nand U29955(G2730,n28117,n28118,n28119,n28120);
  nor U29956(n28120,n28121,n28122,n28123);
  nor U29957(n28123,n28124,n28058);
  nor U29958(n28122,n28076,n28125);
  nor U29959(n28121,n28126,n28062);
  nand U29960(n28119,n28127,n28064);
  nand U29961(n28118,n28065,n28128);
  nand U29962(n28117,n28067,G59303);
  nand U29963(G2729,n28129,n28130,n28131,n28132);
  nor U29964(n28132,n28133,n28134,n28135);
  nor U29965(n28135,n28136,n28058);
  and U29966(n28134,n28059,n28137);
  nor U29967(n28133,n28138,n28062);
  nand U29968(n28131,n28139,n28064);
  nand U29969(n28130,n28065,n28140);
  nand U29970(n28129,n28067,G59302);
  nand U29971(G2728,n28141,n28142,n28143,n28144);
  nor U29972(n28144,n28145,n28146,n28147);
  nor U29973(n28147,n28148,n28058);
  nor U29974(n28146,n28076,n28149);
  nor U29975(n28145,n28150,n28062);
  nand U29976(n28143,n28151,n28064);
  nand U29977(n28142,n28065,n28152);
  nand U29978(n28141,n28067,G59301);
  nand U29979(G2727,n28153,n28154,n28155,n28156);
  nor U29980(n28156,n28157,n28158,n28159);
  nor U29981(n28159,n28160,n28058);
  nor U29982(n28158,n28076,n28161);
  nor U29983(n28157,n28162,n28062);
  nand U29984(n28155,n28163,n28064);
  nand U29985(n28154,n28065,n28164);
  nand U29986(n28153,n28067,G59300);
  nand U29987(G2726,n28165,n28166,n28167,n28168);
  nor U29988(n28168,n28169,n28170,n28171);
  nor U29989(n28171,n28172,n28058);
  and U29990(n28170,n28059,n28173);
  nor U29991(n28169,n28174,n28062);
  nand U29992(n28167,n28175,n28064);
  nand U29993(n28166,n28065,n28176);
  nand U29994(n28165,n28067,G59299);
  nand U29995(G2725,n28177,n28178,n28179,n28180);
  nor U29996(n28180,n28181,n28182,n28183);
  nor U29997(n28183,n28184,n28058);
  nor U29998(n28182,n28076,n28185);
  nor U29999(n28181,n28186,n28062);
  nand U30000(n28179,n28187,n28064);
  nand U30001(n28178,n28065,n28188);
  nand U30002(n28177,n28067,G59298);
  nand U30003(G2724,n28189,n28190,n28191,n28192);
  nor U30004(n28192,n28193,n28194,n28195);
  nor U30005(n28195,n28196,n28058);
  nor U30006(n28194,n28076,n28197);
  nor U30007(n28193,n28198,n28062);
  nand U30008(n28191,n28199,n28064);
  nand U30009(n28190,n28065,n28200);
  nand U30010(n28189,n28067,G59297);
  nand U30011(G2723,n28201,n28202,n28203,n28204);
  nor U30012(n28204,n28205,n28206,n28207,n28208);
  nor U30013(n28208,n28209,n28210);
  and U30014(n28207,G59296,n28067);
  and U30015(n28206,n28211,n28065);
  nand U30016(n28203,n28212,G59328);
  nand U30017(n28202,n28213,n28059);
  nand U30018(n28201,n28214,G59169);
  nand U30019(G2722,n28215,n28216,n28217,n28218);
  nor U30020(n28218,n28205,n28219,n28220,n28221);
  nor U30021(n28221,n28209,n28222);
  and U30022(n28220,G59295,n28067);
  and U30023(n28219,n28223,n28065);
  nand U30024(n28217,n28212,G59327);
  nand U30025(n28216,n28224,n28059);
  nand U30026(n28215,n28214,G59168);
  nand U30027(G2721,n28225,n28226,n28227,n28228);
  nor U30028(n28228,n28205,n28229,n28230,n28231);
  nor U30029(n28231,n28209,n28232);
  and U30030(n28230,G59294,n28067);
  and U30031(n28229,n28233,n28065);
  nand U30032(n28227,n28212,G59326);
  nand U30033(n28226,n28234,n28059);
  nand U30034(n28225,n28214,G59167);
  nand U30035(G2720,n28235,n28236,n28237,n28238);
  nor U30036(n28238,n28205,n28239,n28240,n28241);
  nor U30037(n28241,n28209,n28242);
  and U30038(n28240,G59293,n28067);
  and U30039(n28239,n28243,n28065);
  nand U30040(n28237,n28212,G59325);
  nand U30041(n28236,n28244,n28059);
  nand U30042(n28235,n28214,G59166);
  nand U30043(G2719,n28245,n28246,n28247,n28248);
  nor U30044(n28248,n28205,n28249,n28250,n28251);
  nor U30045(n28251,n28209,n28252);
  and U30046(n28250,G59292,n28067);
  and U30047(n28249,n28253,n28065);
  nand U30048(n28247,n28212,G59324);
  nand U30049(n28246,n28254,n28059);
  nand U30050(n28245,n28214,G59165);
  nand U30051(G2718,n28255,n28256,n28257,n28258);
  nor U30052(n28258,n28205,n28259,n28260,n28261);
  nor U30053(n28261,n28209,n28262);
  and U30054(n28260,G59291,n28067);
  and U30055(n28259,n28263,n28065);
  nand U30056(n28257,n28212,G59323);
  nand U30057(n28256,n28264,n28059);
  nand U30058(n28255,n28214,G59164);
  nand U30059(G2717,n28265,n28266,n28267,n28268);
  nor U30060(n28268,n28205,n28269,n28270,n28271);
  nor U30061(n28271,n28209,n28272);
  and U30062(n28270,G59290,n28067);
  and U30063(n28269,n28065,n28273);
  nand U30064(n28267,n28212,G59322);
  nand U30065(n28266,n28274,n28059);
  nand U30066(n28265,n28214,G59163);
  nand U30067(G2716,n28275,n28276,n28277,n28278);
  nor U30068(n28278,n28205,n28279,n28280,n28281);
  nor U30069(n28281,n28209,n28282);
  and U30070(n28280,G59289,n28067);
  and U30071(n28279,n28283,n28065);
  nand U30072(n28277,n28212,G59321);
  nand U30073(n28276,n28284,n28059);
  nand U30074(n28275,n28214,G59162);
  nand U30075(G2715,n28285,n28286,n28287,n28288);
  nor U30076(n28288,n28205,n28289,n28290,n28291);
  nor U30077(n28291,n28209,n28292);
  and U30078(n28290,G59288,n28067);
  and U30079(n28289,n28293,n28065);
  nand U30080(n28287,n28212,G59320);
  nand U30081(n28286,n28294,n28059);
  nand U30082(n28285,n28214,G59161);
  nand U30083(G2714,n28295,n28296,n28297,n28298);
  nor U30084(n28298,n28205,n28299,n28300,n28301);
  nor U30085(n28301,n28209,n28302);
  nor U30086(n28300,n28303,n28304);
  nor U30087(n28299,n28305,n28306);
  nand U30088(n28297,n28212,G59319);
  nand U30089(n28296,n28307,n28059);
  nand U30090(n28295,n28214,G59160);
  nand U30091(G2713,n28308,n28309,n28310,n28311);
  nor U30092(n28314,n28209,n28315);
  and U30093(n28313,G59286,n28067);
  and U30094(n28312,n28316,n28065);
  nand U30095(n28310,n28212,G59318);
  nand U30096(n28309,n28317,n28059);
  nand U30097(n28308,n28214,G59159);
  nand U30098(G2712,n28318,n28319,n28320,n28321);
  nor U30099(n28324,n28209,n28325);
  and U30100(n28323,G59285,n28067);
  and U30101(n28322,n28065,n28326);
  nand U30102(n28320,n28212,G59317);
  nand U30103(n28319,n28327,n28059);
  nand U30104(n28318,n28214,G59158);
  nand U30105(G2711,n28328,n28329,n28330,n28331);
  nor U30106(n28334,n28209,n28335);
  and U30107(n28333,G59284,n28067);
  and U30108(n28332,n28065,n28336);
  not U30109(n28065,n28305);
  nand U30110(n28330,n28212,G59316);
  nand U30111(n28329,n28337,n28059);
  nand U30112(n28328,n28214,G59157);
  nand U30113(G2710,n28338,n28339,n28340,n28341);
  nor U30114(n28341,n28205,n28342,n28343,n28344);
  nor U30115(n28344,n28209,n28345);
  nor U30116(n28343,n28346,n28304);
  nor U30117(n28342,n28305,n28347);
  nand U30118(n28340,n28212,G59315);
  nand U30119(n28339,n28348,n28059);
  nand U30120(n28338,n28214,G59156);
  nand U30121(G2709,n28349,n28350,n28351,n28352);
  nor U30122(n28352,n28205,n28353,n28354,n28355);
  nor U30123(n28355,n28209,n28356);
  nor U30124(n28354,n28357,n28304);
  and U30125(n28353,n28358,n28359);
  nand U30126(n28351,n28212,G59314);
  nand U30127(n28350,n28360,n28361);
  nand U30128(n28349,n28214,G59155);
  nand U30129(G2708,n28362,n28363,n28364,n28365);
  nor U30130(n28365,n28205,n28366,n28367,n28368);
  nor U30131(n28368,n28209,n28369);
  not U30132(n28209,n28064);
  nor U30133(n28367,n28370,n28304);
  and U30134(n28366,n28358,n28371);
  nor U30135(n28205,G58978,G58979,n28212);
  nand U30136(n28364,n28212,G59313);
  nand U30137(n28363,n27871,n28361);
  nand U30138(n28362,n28214,G59154);
  nand U30139(G2707,n28372,n28373,n28374,n28375);
  nor U30140(n28375,n28376,n28377,n28378);
  nor U30141(n28378,n28379,n28058);
  nor U30142(n28377,n28380,n28381);
  nor U30143(n28376,n28382,n28062);
  nand U30144(n28374,n28383,n28064);
  nand U30145(n28373,n28384,n28358);
  nand U30146(n28372,n28067,G59280);
  nand U30147(G2706,n28385,n28386,n28387,n28388);
  nor U30148(n28388,n28389,n28390,n28391);
  nor U30149(n28391,n28392,n28058);
  nor U30150(n28390,n28380,n28393);
  nor U30151(n28389,n28394,n28062);
  nand U30152(n28387,n28395,n28064);
  nand U30153(n28386,n28396,n28358);
  nand U30154(n28385,n28067,G59279);
  nand U30155(G2705,n28397,n28398,n28399,n28400);
  nor U30156(n28400,n28401,n28402,n28403);
  nor U30157(n28403,n28404,n28058);
  nor U30158(n28402,n28380,n28405);
  nor U30159(n28401,n28015,n28062);
  nand U30160(n28399,n28406,n28064);
  nand U30161(n28398,n28407,n28358);
  nand U30162(n28397,n28067,G59278);
  nand U30163(G2704,n28408,n28409,n28410,n28411);
  nor U30164(n28411,n28412,n28413,n28414);
  nor U30165(n28414,n28415,n28058);
  not U30166(n28058,n28214);
  nor U30167(n28214,n28212,G58977,n28416);
  nor U30168(n28413,n28380,n28417);
  not U30169(n28380,n28361);
  nand U30170(n28361,n28076,n28418);
  nand U30171(n28418,n28419,n27942,n28420);
  not U30172(n28076,n28059);
  nand U30173(n28059,n28421,n28422);
  nand U30174(n28422,n28063,n28062,G58978);
  nand U30175(n28421,n28423,n28424,n28420);
  nor U30176(n28412,n28013,n28062);
  nand U30177(n28410,n27969,n28064);
  nand U30178(n28064,n28425,n28426);
  nand U30179(n28426,n28420,n28424,n28427,n28428);
  not U30180(n28427,n28429);
  nand U30181(n28425,G58978,n28062,n28430);
  nand U30182(n28409,n28431,n28358);
  nand U30183(n28358,n28432,n28305);
  nand U30184(n28305,n28420,n28423,n27945,n28433);
  nand U30185(n28432,n28062,n28419,n27946);
  nand U30186(n28408,n28067,G59277);
  not U30187(n28067,n28304);
  nand U30188(n28304,n28420,n28434);
  nand U30189(n28434,n28435,n28436);
  nand U30190(n28436,n28429,n28428,n28424);
  not U30191(n28428,n28423);
  nand U30192(n28435,n28433,n28437);
  nand U30193(n28437,n28423,n27945);
  nor U30194(n28420,n27929,n28212);
  not U30195(n28212,n28062);
  nand U30196(n28062,n27924,n28438,n28439,n28440);
  nor U30197(n27924,n28441,n28442);
  nor U30198(n28442,n27995,n27916);
  nor U30199(n27995,n28443,n28444);
  nor U30200(n28444,n28445,n27929,n28446);
  nor U30201(n28443,n28447,n28448);
  nand U30202(G2703,n28449,n28450);
  nand U30203(n28450,n28451,n28063);
  nand U30204(n28449,n28452,G59308);
  nand U30205(G2702,n28453,n28454,n28455);
  nand U30206(n28455,n28452,G59307);
  nand U30207(n28454,n28451,n28079);
  nand U30208(n28453,n28456,n28457);
  nand U30209(G2701,n28458,n28459,n28460);
  nand U30210(n28460,n28452,G59306);
  nand U30211(n28459,n28451,n28091);
  nand U30212(n28458,n28456,n28461);
  nand U30213(G2700,n28462,n28463,n28464);
  nand U30214(n28464,n28452,G59305);
  nand U30215(n28463,n28451,n28103);
  nand U30216(n28462,n28456,n28465);
  nand U30217(G2699,n28466,n28467,n28468);
  nand U30218(n28468,n28452,G59304);
  nand U30219(n28467,n28451,n28115);
  nand U30220(n28466,n28456,n28469);
  nand U30221(G2698,n28470,n28471,n28472);
  nand U30222(n28472,n28452,G59303);
  nand U30223(n28471,n28451,n28127);
  nand U30224(n28470,n28456,n28473);
  nand U30225(G2697,n28474,n28475,n28476);
  nand U30226(n28476,n28452,G59302);
  nand U30227(n28475,n28451,n28139);
  nand U30228(n28474,n28456,n28137);
  nand U30229(G2696,n28477,n28478,n28479);
  nand U30230(n28479,n28452,G59301);
  nand U30231(n28478,n28451,n28151);
  nand U30232(n28477,n28456,n28480);
  nand U30233(G2695,n28481,n28482,n28483);
  nand U30234(n28483,n28452,G59300);
  nand U30235(n28482,n28451,n28163);
  nand U30236(n28481,n28456,n28484);
  nand U30237(G2694,n28485,n28486,n28487);
  nand U30238(n28487,n28452,G59299);
  nand U30239(n28486,n28451,n28175);
  nand U30240(n28485,n28456,n28173);
  nand U30241(G2693,n28488,n28489,n28490);
  nand U30242(n28490,n28452,G59298);
  nand U30243(n28489,n28451,n28187);
  nand U30244(n28488,n28456,n28491);
  nand U30245(G2692,n28492,n28493,n28494);
  nand U30246(n28494,n28452,G59297);
  nand U30247(n28493,n28451,n28199);
  nand U30248(n28492,n28456,n28495);
  nand U30249(G2691,n28496,n28497,n28498);
  nand U30250(n28498,n28452,G59296);
  nand U30251(n28497,n28451,n28499);
  nand U30252(n28496,n28456,n28213);
  nand U30253(G2690,n28500,n28501,n28502);
  nand U30254(n28502,n28452,G59295);
  nand U30255(n28501,n28451,n28503);
  nand U30256(n28500,n28456,n28224);
  nand U30257(G2689,n28504,n28505,n28506);
  nand U30258(n28506,n28452,G59294);
  nand U30259(n28505,n28451,n28507);
  nand U30260(n28504,n28456,n28234);
  nand U30261(G2688,n28508,n28509,n28510);
  nand U30262(n28510,n28452,G59293);
  nand U30263(n28509,n28451,n28511);
  nand U30264(n28508,n28456,n28244);
  nand U30265(G2687,n28512,n28513,n28514);
  nand U30266(n28514,n28452,G59292);
  nand U30267(n28513,n28451,n28515);
  nand U30268(n28512,n28456,n28254);
  nand U30269(G2686,n28516,n28517,n28518);
  nand U30270(n28518,n28452,G59291);
  nand U30271(n28517,n28451,n28519);
  nand U30272(n28516,n28456,n28264);
  nand U30273(G2685,n28520,n28521,n28522);
  nand U30274(n28522,n28452,G59290);
  nand U30275(n28521,n28451,n28523);
  nand U30276(n28520,n28456,n28274);
  nand U30277(G2684,n28524,n28525,n28526);
  nand U30278(n28526,n28452,G59289);
  nand U30279(n28525,n28451,n28527);
  nand U30280(n28524,n28456,n28284);
  nand U30281(G2683,n28528,n28529,n28530);
  nand U30282(n28530,n28452,G59288);
  nand U30283(n28529,n28451,n28531);
  nand U30284(n28528,n28456,n28294);
  nand U30285(G2682,n28532,n28533,n28534);
  nand U30286(n28534,n28452,G59287);
  nand U30287(n28533,n28451,n28535);
  nand U30288(n28532,n28456,n28307);
  nand U30289(G2681,n28536,n28537,n28538);
  nand U30290(n28538,n28452,G59286);
  nand U30291(n28537,n28451,n28539);
  nand U30292(n28536,n28456,n28317);
  nand U30293(G2680,n28540,n28541,n28542);
  nand U30294(n28542,n28452,G59285);
  nand U30295(n28541,n28451,n28543);
  nand U30296(n28540,n28456,n28327);
  nand U30297(G2679,n28544,n28545,n28546);
  nand U30298(n28546,n28452,G59284);
  nand U30299(n28545,n28451,n28547);
  nand U30300(n28544,n28456,n28337);
  nand U30301(G2678,n28548,n28549,n28550);
  nand U30302(n28550,n28452,G59283);
  nand U30303(n28549,n28451,n28551);
  nand U30304(n28548,n28456,n28348);
  nand U30305(G2677,n28552,n28553,n28554);
  nand U30306(n28554,n28452,G59282);
  nand U30307(n28553,n28451,n28555);
  nand U30308(n28552,n28456,n28360);
  nand U30309(G2676,n28556,n28557,n28558);
  nand U30310(n28558,n28452,G59281);
  nand U30311(n28557,n28451,n28559);
  nand U30312(n28556,n28456,n27871);
  nand U30313(G2675,n28560,n28561,n28562);
  nand U30314(n28562,n28452,G59280);
  nand U30315(n28561,n28451,n28383);
  nand U30316(n28560,n28456,n27881);
  nand U30317(G2674,n28563,n28564,n28565);
  nand U30318(n28565,n28452,G59279);
  nand U30319(n28564,n28451,n28395);
  nand U30320(n28563,n28456,n27891);
  nand U30321(G2673,n28566,n28567,n28568);
  nand U30322(n28568,n28452,G59278);
  nand U30323(n28567,n28451,n28406);
  nand U30324(n28566,n28456,n27900);
  nand U30325(G2672,n28569,n28570,n28571);
  nand U30326(n28571,n28452,G59277);
  nand U30327(n28570,n28451,n27969);
  nand U30328(n28569,n28456,n27915);
  nand U30329(n28574,n28577,n27907);
  nand U30330(G2671,n28578,n28579,n28580);
  nand U30331(n28580,n28581,G59276);
  nand U30332(n28579,n28582,G58902);
  nand U30333(n28578,n28583,n28063);
  nand U30334(G2670,n28584,n28585,n28586);
  nor U30335(n28586,n28587,n28588,n28589);
  nor U30336(n28589,n28590,n22157);
  not U30337(n22157,G58885);
  nor U30338(n28588,n21709,n28591);
  not U30339(n21709,G58901);
  nor U30340(n28587,n28592,n28593);
  nand U30341(n28585,n28594,n28080);
  nand U30342(n28584,n28581,G59275);
  nand U30343(G2669,n28595,n28596,n28597);
  nor U30344(n28597,n28598,n28599,n28600);
  nor U30345(n28600,n28590,n22151);
  not U30346(n22151,G58884);
  nor U30347(n28599,n21722,n28591);
  not U30348(n21722,G58900);
  nor U30349(n28598,n28601,n28593);
  nand U30350(n28596,n28594,n28092);
  nand U30351(n28595,n28581,G59274);
  nand U30352(G2668,n28602,n28603,n28604);
  nor U30353(n28604,n28605,n28606,n28607);
  nor U30354(n28607,n28590,n22145);
  not U30355(n22145,G58883);
  nor U30356(n28606,n21732,n28591);
  not U30357(n21732,G58899);
  nor U30358(n28605,n28608,n28593);
  nand U30359(n28603,n28594,n28104);
  nand U30360(n28602,n28581,G59273);
  nand U30361(G2667,n28609,n28610,n28611);
  nor U30362(n28611,n28612,n28613,n28614);
  nor U30363(n28614,n28590,n22139);
  not U30364(n22139,G58882);
  nor U30365(n28613,n21742,n28591);
  not U30366(n21742,G58898);
  nor U30367(n28612,n28615,n28593);
  nand U30368(n28610,n28594,n28116);
  nand U30369(n28609,n28581,G59272);
  nand U30370(G2666,n28616,n28617,n28618);
  nor U30371(n28618,n28619,n28620,n28621);
  nor U30372(n28621,n28590,n22133);
  not U30373(n22133,G58881);
  nor U30374(n28620,n21752,n28591);
  not U30375(n21752,G58897);
  nor U30376(n28619,n28622,n28593);
  nand U30377(n28617,n28594,n28128);
  nand U30378(n28616,n28581,G59271);
  nand U30379(G2665,n28623,n28624,n28625);
  nor U30380(n28625,n28626,n28627,n28628);
  nor U30381(n28628,n28590,n22127);
  not U30382(n22127,G58880);
  nor U30383(n28627,n21762,n28591);
  not U30384(n21762,G58896);
  nor U30385(n28626,n28629,n28593);
  nand U30386(n28624,n28594,n28140);
  nand U30387(n28623,n28581,G59270);
  nand U30388(G2664,n28630,n28631,n28632);
  nor U30389(n28632,n28633,n28634,n28635);
  nor U30390(n28635,n28590,n22121);
  not U30391(n22121,G58879);
  nor U30392(n28634,n21772,n28591);
  not U30393(n21772,G58895);
  nor U30394(n28633,n28636,n28593);
  nand U30395(n28631,n28594,n28152);
  nand U30396(n28630,n28581,G59269);
  nand U30397(G2663,n28637,n28638,n28639);
  nor U30398(n28639,n28640,n28641,n28642);
  nor U30399(n28642,n28590,n26913);
  nor U30400(n28641,n28591,n26905);
  nor U30401(n28640,n28643,n28593);
  nand U30402(n28638,n28594,n28164);
  nand U30403(n28637,n28581,G59268);
  nand U30404(G2662,n28644,n28645,n28646);
  nor U30405(n28646,n28647,n28648,n28649);
  nor U30406(n28649,n28590,n26883);
  nor U30407(n28648,n28591,n26878);
  nor U30408(n28647,n28650,n28593);
  nand U30409(n28645,n28594,n28176);
  nand U30410(n28644,n28581,G59267);
  nand U30411(G2661,n28651,n28652,n28653);
  nor U30412(n28653,n28654,n28655,n28656);
  nor U30413(n28656,n28590,n26866);
  nor U30414(n28655,n28591,n26860);
  nor U30415(n28654,n28657,n28593);
  nand U30416(n28652,n28594,n28188);
  nand U30417(n28651,n28581,G59266);
  nand U30418(G2660,n28658,n28659,n28660);
  nor U30419(n28660,n28661,n28662,n28663);
  nor U30420(n28663,n28590,n26848);
  nor U30421(n28662,n28591,n26843);
  nor U30422(n28661,n28664,n28593);
  nand U30423(n28659,n28594,n28200);
  nand U30424(n28658,n28581,G59265);
  nand U30425(G2659,n28665,n28666,n28667);
  nor U30426(n28667,n28668,n28669,n28670);
  nor U30427(n28670,n28590,n26831);
  nor U30428(n28669,n28591,n26826);
  nor U30429(n28668,n28210,n28593);
  nand U30430(n28666,n28594,n28211);
  nand U30431(n28665,n28581,G59264);
  nand U30432(G2658,n28671,n28672,n28673);
  nor U30433(n28673,n28674,n28675,n28676);
  nor U30434(n28676,n28590,n26814);
  nor U30435(n28675,n28591,n26809);
  nor U30436(n28674,n28222,n28593);
  nand U30437(n28672,n28594,n28223);
  nand U30438(n28671,n28581,G59263);
  nand U30439(G2657,n28677,n28678,n28679);
  nor U30440(n28679,n28680,n28681,n28682);
  nor U30441(n28682,n28590,n26797);
  nor U30442(n28681,n28591,n26792);
  nor U30443(n28680,n28232,n28593);
  nand U30444(n28678,n28594,n28233);
  nand U30445(n28677,n28581,G59262);
  nand U30446(G2656,n28683,n28684,n28685);
  nor U30447(n28685,n28686,n28687,n28688);
  nor U30448(n28688,n28590,n26779);
  nand U30449(n28590,n28689,n28690);
  nor U30450(n28687,n28591,n26769);
  not U30451(n28591,n28582);
  nor U30452(n28582,n28691,n28581);
  nor U30453(n28686,n28242,n28593);
  not U30454(n28593,n28583);
  nand U30455(n28684,n28594,n28243);
  nand U30456(n28683,n28581,G59261);
  nand U30457(G2655,n28692,n28693,n28694,n28695);
  nand U30458(n28695,n28696,G58886);
  nand U30459(n28694,n28583,n28515);
  nand U30460(n28693,n28594,n28253);
  nand U30461(n28692,n28581,G59260);
  nand U30462(G2654,n28697,n28698,n28699,n28700);
  nand U30463(n28700,n28696,G58885);
  nand U30464(n28699,n28583,n28519);
  nand U30465(n28698,n28594,n28263);
  nand U30466(n28697,n28581,G59259);
  nand U30467(G2653,n28701,n28702,n28703,n28704);
  nand U30468(n28704,n28696,G58884);
  nand U30469(n28703,n28583,n28523);
  nand U30470(n28702,n28594,n28273);
  nand U30471(n28701,n28581,G59258);
  nand U30472(G2652,n28705,n28706,n28707,n28708);
  nand U30473(n28708,n28696,G58883);
  nand U30474(n28707,n28583,n28527);
  nand U30475(n28706,n28594,n28283);
  nand U30476(n28705,n28581,G59257);
  nand U30477(G2651,n28709,n28710,n28711,n28712);
  nand U30478(n28712,n28696,G58882);
  nand U30479(n28711,n28583,n28531);
  nand U30480(n28710,n28594,n28293);
  nand U30481(n28709,n28581,G59256);
  nand U30482(G2650,n28713,n28714,n28715,n28716);
  nand U30483(n28716,n28696,G58881);
  nand U30484(n28715,n28583,n28535);
  nand U30485(n28714,n28594,n28717);
  nand U30486(n28713,n28581,G59255);
  nand U30487(G2649,n28718,n28719,n28720,n28721);
  nand U30488(n28721,n28696,G58880);
  nand U30489(n28720,n28583,n28539);
  nand U30490(n28719,n28594,n28316);
  nand U30491(n28718,n28581,G59254);
  nand U30492(G2648,n28722,n28723,n28724,n28725);
  nand U30493(n28725,n28696,G58879);
  nand U30494(n28724,n28583,n28543);
  nand U30495(n28723,n28594,n28326);
  nand U30496(n28722,n28581,G59253);
  nand U30497(G2647,n28726,n28727,n28728,n28729);
  nand U30498(n28729,n28696,G58878);
  nand U30499(n28728,n28583,n28547);
  nand U30500(n28727,n28594,n28336);
  nand U30501(n28726,n28581,G59252);
  nand U30502(G2646,n28730,n28731,n28732,n28733);
  nand U30503(n28733,n28696,G58877);
  nand U30504(n28732,n28583,n28551);
  nand U30505(n28731,n28594,n28734);
  nand U30506(n28730,n28581,G59251);
  nand U30507(G2645,n28735,n28736,n28737,n28738);
  nand U30508(n28738,n28696,G58876);
  nand U30509(n28737,n28583,n28555);
  nand U30510(n28736,n28594,n28359);
  nand U30511(n28735,n28581,G59250);
  nand U30512(G2644,n28739,n28740,n28741,n28742);
  nand U30513(n28742,n28696,G58875);
  nand U30514(n28741,n28583,n28559);
  nand U30515(n28740,n28594,n28371);
  nand U30516(n28739,n28581,G59249);
  nand U30517(G2643,n28743,n28744,n28745,n28746);
  nand U30518(n28746,n28696,G58874);
  nand U30519(n28745,n28583,n28383);
  nand U30520(n28744,n28594,n28384);
  nand U30521(n28743,n28581,G59248);
  nand U30522(G2642,n28747,n28748,n28749,n28750);
  nand U30523(n28750,n28696,G58873);
  nand U30524(n28749,n28583,n28395);
  nand U30525(n28748,n28594,n28396);
  nand U30526(n28747,n28581,G59247);
  nand U30527(G2641,n28751,n28752,n28753,n28754);
  nand U30528(n28754,n28696,G58872);
  nand U30529(n28753,n28583,n28406);
  nand U30530(n28752,n28594,n28407);
  nand U30531(n28751,n28581,G59246);
  nand U30532(G2640,n28755,n28756,n28757,n28758);
  nand U30533(n28758,n28696,G58871);
  nor U30534(n28696,n28581,n28759);
  nand U30535(n28757,n28583,n27969);
  nor U30536(n28583,n28760,n28581);
  nand U30537(n28756,n28594,n28431);
  nand U30538(n28755,n28581,G59245);
  nand U30539(n28763,n27870,n28764);
  nand U30540(n28764,n28765,n28766);
  nand U30541(n28766,n28767,n27965);
  nand U30542(n28767,n27998,n28768);
  or U30543(n28768,n28769,n28770);
  nor U30544(G2639,n28771,n28772);
  nand U30545(G2638,n28773,n28774,n28775);
  nand U30546(n28775,G59243,n28776);
  nand U30547(n28774,n28777,G59275);
  nand U30548(n28773,G59198,n28778);
  nand U30549(G2637,n28779,n28780,n28781);
  nand U30550(n28781,G59242,n28776);
  nand U30551(n28780,n28777,G59274);
  nand U30552(n28779,G59199,n28778);
  nand U30553(G2636,n28782,n28783,n28784);
  nand U30554(n28784,G59241,n28776);
  nand U30555(n28783,n28777,G59273);
  nand U30556(n28782,G59200,n28778);
  nand U30557(G2635,n28785,n28786,n28787);
  nand U30558(n28787,G59240,n28776);
  nand U30559(n28786,n28777,G59272);
  nand U30560(n28785,G59201,n28778);
  nand U30561(G2634,n28788,n28789,n28790);
  nand U30562(n28790,G59239,n28776);
  nand U30563(n28789,n28777,G59271);
  nand U30564(n28788,G59202,n28778);
  nand U30565(G2633,n28791,n28792,n28793);
  nand U30566(n28793,G59238,n28776);
  nand U30567(n28792,n28777,G59270);
  nand U30568(n28791,G59203,n28778);
  nand U30569(G2632,n28794,n28795,n28796);
  nand U30570(n28796,G59237,n28776);
  nand U30571(n28795,n28777,G59269);
  nand U30572(n28794,G59204,n28778);
  nand U30573(G2631,n28797,n28798,n28799);
  nand U30574(n28799,G59236,n28776);
  nand U30575(n28798,n28777,G59268);
  nand U30576(n28797,G59205,n28778);
  nand U30577(G2630,n28800,n28801,n28802);
  nand U30578(n28802,G59235,n28776);
  nand U30579(n28801,n28777,G59267);
  nand U30580(n28800,G59206,n28778);
  nand U30581(G2629,n28803,n28804,n28805);
  nand U30582(n28805,G59234,n28776);
  nand U30583(n28804,n28777,G59266);
  nand U30584(n28803,G59207,n28778);
  nand U30585(G2628,n28806,n28807,n28808);
  nand U30586(n28808,G59233,n28776);
  nand U30587(n28807,n28777,G59265);
  nand U30588(n28806,G59208,n28778);
  nand U30589(G2627,n28809,n28810,n28811);
  nand U30590(n28811,G59232,n28776);
  nand U30591(n28810,n28777,G59264);
  nand U30592(n28809,G59209,n28778);
  nand U30593(G2626,n28812,n28813,n28814);
  nand U30594(n28814,G59231,n28776);
  nand U30595(n28813,n28777,G59263);
  nand U30596(n28812,G59210,n28778);
  nand U30597(G2625,n28815,n28816,n28817);
  nand U30598(n28817,G59230,n28776);
  nand U30599(n28816,n28777,G59262);
  nand U30600(n28815,G59211,n28778);
  nand U30601(G2624,n28818,n28819,n28820);
  nand U30602(n28820,G59229,n28776);
  nand U30603(n28819,n28777,G59261);
  and U30604(n28777,n28821,n28689);
  nand U30605(n28818,G59212,n28778);
  nand U30606(G2623,n28822,n28823,n28824);
  nand U30607(n28824,G59228,n28776);
  nand U30608(n28823,G59182,n28778);
  nand U30609(n28822,n28821,G59260);
  nand U30610(G2622,n28825,n28826,n28827);
  nand U30611(n28827,G59227,n28776);
  nand U30612(n28826,G59183,n28778);
  nand U30613(n28825,n28821,G59259);
  nand U30614(G2621,n28828,n28829,n28830);
  nand U30615(n28830,G59226,n28776);
  nand U30616(n28829,G59184,n28778);
  nand U30617(n28828,n28821,G59258);
  nand U30618(G2620,n28831,n28832,n28833);
  nand U30619(n28833,G59225,n28776);
  nand U30620(n28832,G59185,n28778);
  nand U30621(n28831,n28821,G59257);
  nand U30622(G2619,n28834,n28835,n28836);
  nand U30623(n28836,G59224,n28776);
  nand U30624(n28835,G59186,n28778);
  nand U30625(n28834,n28821,G59256);
  nand U30626(G2618,n28837,n28838,n28839);
  nand U30627(n28839,G59223,n28776);
  nand U30628(n28838,G59187,n28778);
  nand U30629(n28837,n28821,G59255);
  nand U30630(G2617,n28840,n28841,n28842);
  nand U30631(n28842,G59222,n28776);
  nand U30632(n28841,G59188,n28778);
  nand U30633(n28840,n28821,G59254);
  nand U30634(G2616,n28843,n28844,n28845);
  nand U30635(n28845,G59221,n28776);
  nand U30636(n28844,G59189,n28778);
  nand U30637(n28843,n28821,G59253);
  nand U30638(G2615,n28846,n28847,n28848);
  nand U30639(n28848,G59220,n28776);
  nand U30640(n28847,G59190,n28778);
  nand U30641(n28846,n28821,G59252);
  nand U30642(G2614,n28849,n28850,n28851);
  nand U30643(n28851,G59219,n28776);
  nand U30644(n28850,G59191,n28778);
  nand U30645(n28849,n28821,G59251);
  nand U30646(G2613,n28852,n28853,n28854);
  nand U30647(n28854,G59218,n28776);
  nand U30648(n28853,G59192,n28778);
  nand U30649(n28852,n28821,G59250);
  nand U30650(G2612,n28855,n28856,n28857);
  nand U30651(n28857,G59217,n28776);
  nand U30652(n28856,G59193,n28778);
  nand U30653(n28855,n28821,G59249);
  nand U30654(G2611,n28858,n28859,n28860);
  nand U30655(n28860,G59216,n28776);
  nand U30656(n28859,G59194,n28778);
  nand U30657(n28858,n28821,G59248);
  nand U30658(G2610,n28861,n28862,n28863);
  nand U30659(n28863,G59215,n28776);
  nand U30660(n28862,G59195,n28778);
  nand U30661(n28861,n28821,G59247);
  nand U30662(G2609,n28864,n28865,n28866);
  nand U30663(n28866,G59214,n28776);
  nand U30664(n28865,G59196,n28778);
  nand U30665(n28864,n28821,G59246);
  nand U30666(G2608,n28867,n28868,n28869);
  nand U30667(n28869,G59213,n28776);
  nand U30668(n28868,G59197,n28778);
  nand U30669(n28867,n28821,G59245);
  nor U30670(n28821,n28416,n28776);
  nand U30671(n28771,n28870,n28871);
  nand U30672(n28871,n28872,n27965);
  nand U30673(n28872,n28873,n28874);
  nand U30674(n28874,n27907,n27945,n28875);
  nand U30675(n28873,n27870,n28876,n28877);
  nand U30676(n28870,n27931,G58978);
  nand U30677(G2607,n28878,n28879,n28880);
  nand U30678(n28880,n28881,G59212);
  nand U30679(n28878,n28882,G59261);
  nand U30680(G2606,n28883,n28884,n28885);
  nand U30681(n28885,n28881,G59211);
  nand U30682(n28883,n28882,G59262);
  nand U30683(G2605,n28886,n28887,n28888);
  nand U30684(n28888,n28881,G59210);
  nand U30685(n28886,n28882,G59263);
  nand U30686(G2604,n28889,n28890,n28891);
  nand U30687(n28891,n28881,G59209);
  nand U30688(n28889,n28882,G59264);
  nand U30689(G2603,n28892,n28893,n28894);
  nand U30690(n28894,n28881,G59208);
  nand U30691(n28892,n28882,G59265);
  nand U30692(G2602,n28895,n28896,n28897);
  nand U30693(n28897,n28881,G59207);
  nand U30694(n28895,n28882,G59266);
  nand U30695(G2601,n28898,n28899,n28900);
  nand U30696(n28900,n28881,G59206);
  nand U30697(n28898,n28882,G59267);
  nand U30698(G2600,n28901,n28902,n28903);
  nand U30699(n28903,n28881,G59205);
  nand U30700(n28901,n28882,G59268);
  nand U30701(G2599,n28904,n28905,n28906);
  nand U30702(n28906,n28881,G59204);
  nand U30703(n28904,n28882,G59269);
  nand U30704(G2598,n28907,n28908,n28909);
  nand U30705(n28909,n28881,G59203);
  nand U30706(n28907,n28882,G59270);
  nand U30707(G2597,n28910,n28911,n28912);
  nand U30708(n28912,n28881,G59202);
  nand U30709(n28910,n28882,G59271);
  nand U30710(G2596,n28913,n28914,n28915);
  nand U30711(n28915,n28881,G59201);
  nand U30712(n28913,n28882,G59272);
  nand U30713(G2595,n28916,n28917,n28918);
  nand U30714(n28918,n28881,G59200);
  nand U30715(n28916,n28882,G59273);
  nand U30716(G2594,n28919,n28920,n28921);
  nand U30717(n28921,n28881,G59199);
  nand U30718(n28919,n28882,G59274);
  nand U30719(G2593,n28922,n28923,n28924);
  nand U30720(n28924,n28881,G59198);
  nand U30721(n28922,n28882,G59275);
  nand U30722(G2592,n28925,n28879,n28926);
  nand U30723(n28926,n28881,G59197);
  nand U30724(n28879,n28927,G58871);
  nand U30725(n28925,n28882,G59245);
  nand U30726(G2591,n28928,n28884,n28929);
  nand U30727(n28929,n28881,G59196);
  nand U30728(n28884,n28927,G58872);
  nand U30729(n28928,n28882,G59246);
  nand U30730(G2590,n28930,n28887,n28931);
  nand U30731(n28931,n28881,G59195);
  nand U30732(n28887,n28927,G58873);
  nand U30733(n28930,n28882,G59247);
  nand U30734(G2589,n28932,n28890,n28933);
  nand U30735(n28933,n28881,G59194);
  nand U30736(n28890,n28927,G58874);
  nand U30737(n28932,n28882,G59248);
  nand U30738(G2588,n28934,n28893,n28935);
  nand U30739(n28935,n28881,G59193);
  nand U30740(n28893,n28927,G58875);
  nand U30741(n28934,n28882,G59249);
  nand U30742(G2587,n28936,n28896,n28937);
  nand U30743(n28937,n28881,G59192);
  nand U30744(n28896,n28927,G58876);
  nand U30745(n28936,n28882,G59250);
  nand U30746(G2586,n28938,n28899,n28939);
  nand U30747(n28939,n28881,G59191);
  nand U30748(n28899,n28927,G58877);
  nand U30749(n28938,n28882,G59251);
  nand U30750(G2585,n28940,n28902,n28941);
  nand U30751(n28941,n28881,G59190);
  nand U30752(n28902,n28927,G58878);
  nand U30753(n28940,n28882,G59252);
  nand U30754(G2584,n28942,n28905,n28943);
  nand U30755(n28943,n28881,G59189);
  nand U30756(n28905,n28927,G58879);
  nand U30757(n28942,n28882,G59253);
  nand U30758(G2583,n28944,n28908,n28945);
  nand U30759(n28945,n28881,G59188);
  nand U30760(n28908,n28927,G58880);
  nand U30761(n28944,n28882,G59254);
  nand U30762(G2582,n28946,n28911,n28947);
  nand U30763(n28947,n28881,G59187);
  nand U30764(n28911,n28927,G58881);
  nand U30765(n28946,n28882,G59255);
  nand U30766(G2581,n28948,n28914,n28949);
  nand U30767(n28949,n28881,G59186);
  nand U30768(n28914,n28927,G58882);
  nand U30769(n28948,n28882,G59256);
  nand U30770(G2580,n28950,n28917,n28951);
  nand U30771(n28951,n28881,G59185);
  nand U30772(n28917,n28927,G58883);
  nand U30773(n28950,n28882,G59257);
  nand U30774(G2579,n28952,n28920,n28953);
  nand U30775(n28953,n28881,G59184);
  nand U30776(n28920,n28927,G58884);
  nand U30777(n28952,n28882,G59258);
  nand U30778(G2578,n28954,n28923,n28955);
  nand U30779(n28955,n28881,G59183);
  nand U30780(n28923,n28927,G58885);
  nand U30781(n28954,n28882,G59259);
  nand U30782(G2577,n28956,n28957,n28958);
  nand U30783(n28958,n28881,G59182);
  nand U30784(n28957,n28927,G58886);
  nor U30785(n28927,n28959,n28881);
  nand U30786(n28956,n28882,G59260);
  nand U30787(n28960,n27907,n27965,n28961);
  nand U30788(n28762,n28441,n27930);
  nor U30789(n28441,n28962,n27990,n28963);
  nand U30790(G2576,n28964,n28965,n28966,n28967);
  nor U30791(n28967,n28968,n28969);
  nor U30792(n28969,n28057,n28970);
  nor U30793(n28968,n28430,n28971);
  nand U30794(n28966,n28972,n28066);
  nand U30795(n28965,n28973,G59340);
  nand U30796(n28964,n28974,n28060);
  nand U30797(G2575,n28975,n28976,n28977,n28978);
  nor U30798(n28978,n28979,n28980);
  nor U30799(n28980,n28075,n28970);
  nor U30800(n28979,n28592,n28971);
  nand U30801(n28977,n28972,n28080);
  nand U30802(n28976,n28973,G59339);
  nand U30803(n28975,n28974,n28457);
  nand U30804(G2574,n28981,n28982,n28983,n28984);
  nor U30805(n28984,n28985,n28986);
  nor U30806(n28986,n28088,n28970);
  nor U30807(n28985,n28601,n28971);
  nand U30808(n28983,n28972,n28092);
  nand U30809(n28982,n28973,G59338);
  nand U30810(n28981,n28974,n28461);
  nand U30811(G2573,n28987,n28988,n28989,n28990);
  nor U30812(n28990,n28991,n28992);
  nor U30813(n28992,n28100,n28970);
  nor U30814(n28991,n28608,n28971);
  nand U30815(n28989,n28972,n28104);
  nand U30816(n28988,n28973,G59337);
  nand U30817(n28987,n28974,n28465);
  nand U30818(G2572,n28993,n28994,n28995,n28996);
  nor U30819(n28996,n28997,n28998);
  nor U30820(n28998,n28112,n28970);
  nor U30821(n28997,n28615,n28971);
  not U30822(n28615,n28115);
  nand U30823(n28995,n28972,n28116);
  nand U30824(n28994,n28973,G59336);
  nand U30825(n28993,n28974,n28469);
  nand U30826(G2571,n28999,n29000,n29001,n29002);
  nor U30827(n29002,n29003,n29004);
  nor U30828(n29004,n28124,n28970);
  nor U30829(n29003,n28622,n28971);
  nand U30830(n29001,n28972,n28128);
  nand U30831(n29000,n28973,G59335);
  nand U30832(n28999,n28974,n28473);
  nand U30833(G2570,n29005,n29006,n29007,n29008);
  nor U30834(n29008,n29009,n29010);
  nor U30835(n29010,n28136,n28970);
  nor U30836(n29009,n28629,n28971);
  nand U30837(n29007,n28972,n28140);
  nand U30838(n29006,n28973,G59334);
  nand U30839(n29005,n28974,n28137);
  nand U30840(G2569,n29011,n29012,n29013,n29014);
  nor U30841(n29014,n29015,n29016);
  nor U30842(n29016,n28148,n28970);
  nor U30843(n29015,n28636,n28971);
  nand U30844(n29013,n28972,n28152);
  nand U30845(n29012,n28973,G59333);
  nand U30846(n29011,n28974,n28480);
  nand U30847(G2568,n29017,n29018,n29019,n29020);
  nor U30848(n29020,n29021,n29022);
  nor U30849(n29022,n28160,n28970);
  nor U30850(n29021,n28643,n28971);
  nand U30851(n29019,n28972,n28164);
  nand U30852(n29018,n28973,G59332);
  nand U30853(n29017,n28974,n28484);
  nand U30854(G2567,n29023,n29024,n29025,n29026);
  nor U30855(n29026,n29027,n29028);
  nor U30856(n29028,n28172,n28970);
  not U30857(n28172,G59172);
  nor U30858(n29027,n28650,n28971);
  nand U30859(n29025,n28972,n28176);
  nand U30860(n29024,n28973,G59331);
  nand U30861(n29023,n28974,n28173);
  nand U30862(G2566,n29029,n29030,n29031,n29032);
  nor U30863(n29032,n29033,n29034);
  nor U30864(n29034,n28184,n28970);
  not U30865(n28184,G59171);
  nor U30866(n29033,n28657,n28971);
  nand U30867(n29031,n28972,n28188);
  nand U30868(n29030,n28973,G59330);
  nand U30869(n29029,n28974,n28491);
  nand U30870(G2565,n29035,n29036,n29037,n29038);
  nor U30871(n29038,n29039,n29040);
  nor U30872(n29040,n28196,n28970);
  not U30873(n28196,G59170);
  nor U30874(n29039,n28664,n28971);
  nand U30875(n29037,n28972,n28200);
  nand U30876(n29036,n28973,G59329);
  nand U30877(n29035,n28974,n28495);
  nand U30878(G2564,n29041,n29042,n29043,n29044);
  nor U30879(n29044,n29045,n29046);
  and U30880(n29046,G59169,n29047);
  nor U30881(n29045,n28210,n28971);
  nand U30882(n29043,n28972,n28211);
  nand U30883(n29042,n28973,G59328);
  nand U30884(n29041,n28974,n28213);
  nand U30885(G2563,n29048,n29049,n29050,n29051);
  nor U30886(n29051,n29052,n29053);
  and U30887(n29053,G59168,n29047);
  nor U30888(n29052,n28222,n28971);
  nand U30889(n29050,n28972,n28223);
  nand U30890(n29049,n28973,G59327);
  nand U30891(n29048,n28974,n28224);
  nand U30892(G2562,n29054,n29055,n29056,n29057);
  nor U30893(n29057,n29058,n29059);
  and U30894(n29059,G59167,n29047);
  nor U30895(n29058,n28232,n28971);
  nand U30896(n29056,n28972,n28233);
  nand U30897(n29055,n28973,G59326);
  nand U30898(n29054,n28974,n28234);
  nand U30899(G2561,n29060,n29061,n29062,n29063);
  nor U30900(n29063,n29064,n29065);
  and U30901(n29065,G59166,n29047);
  nor U30902(n29064,n28242,n28971);
  nand U30903(n29062,n28972,n28243);
  nand U30904(n29061,n28973,G59325);
  nand U30905(n29060,n28974,n28244);
  nand U30906(G2560,n29066,n29067,n29068,n29069);
  nor U30907(n29069,n29070,n29071);
  and U30908(n29071,G59165,n29047);
  nor U30909(n29070,n28252,n28971);
  nand U30910(n29068,n28972,n28253);
  nand U30911(n29067,n28973,G59324);
  nand U30912(n29066,n28974,n28254);
  nand U30913(G2559,n29072,n29073,n29074,n29075);
  nor U30914(n29075,n29076,n29077);
  and U30915(n29077,G59164,n29047);
  nor U30916(n29076,n28262,n28971);
  nand U30917(n29074,n28972,n28263);
  nand U30918(n29073,n28973,G59323);
  nand U30919(n29072,n28974,n28264);
  nand U30920(G2558,n29078,n29079,n29080,n29081);
  nor U30921(n29081,n29082,n29083);
  and U30922(n29083,G59163,n29047);
  nor U30923(n29082,n28272,n28971);
  nand U30924(n29080,n28972,n28273);
  nand U30925(n29079,n28973,G59322);
  nand U30926(n29078,n28974,n28274);
  nand U30927(G2557,n29084,n29085,n29086,n29087);
  nor U30928(n29087,n29088,n29089);
  and U30929(n29089,G59162,n29047);
  nor U30930(n29088,n28282,n28971);
  nand U30931(n29086,n28972,n28283);
  nand U30932(n29085,n28973,G59321);
  nand U30933(n29084,n28974,n28284);
  nand U30934(G2556,n29090,n29091,n29092,n29093);
  nor U30935(n29093,n29094,n29095);
  and U30936(n29095,G59161,n29047);
  nor U30937(n29094,n28292,n28971);
  nand U30938(n29092,n28972,n28293);
  nand U30939(n29091,n28973,G59320);
  nand U30940(n29090,n28974,n28294);
  nand U30941(G2555,n29096,n29097,n29098);
  nor U30942(n29098,n29099,n29100,n29101);
  nor U30943(n29101,n29102,n29103);
  nor U30944(n29100,n29104,n29105);
  and U30945(n29099,n28717,n28972);
  nand U30946(n29097,n29106,n28535);
  nand U30947(n29096,n29047,G59160);
  nand U30948(G2554,n29107,n29108,n29109,n29110);
  nor U30949(n29110,n29111,n29112);
  and U30950(n29112,G59159,n29047);
  nor U30951(n29111,n28315,n28971);
  nand U30952(n29109,n28972,n28316);
  nand U30953(n29108,n28973,G59318);
  nand U30954(n29107,n28974,n28317);
  nand U30955(G2553,n29113,n29114,n29115,n29116);
  nor U30956(n29116,n29117,n29118);
  and U30957(n29118,G59158,n29047);
  nor U30958(n29117,n28325,n28971);
  not U30959(n28325,n28543);
  nand U30960(n29115,n28972,n28326);
  nand U30961(n29114,n28973,G59317);
  nand U30962(n29113,n28974,n28327);
  nand U30963(G2552,n29119,n29120,n29121,n29122);
  nor U30964(n29122,n29123,n29124);
  and U30965(n29124,G59157,n29047);
  nor U30966(n29123,n28335,n28971);
  nand U30967(n29121,n28972,n28336);
  nand U30968(n29120,n28973,G59316);
  nand U30969(n29119,n28974,n28337);
  nand U30970(G2551,n29125,n29126,n29127,n29128);
  nor U30971(n29128,n29129,n29130);
  nor U30972(n29130,n29131,n28970);
  nor U30973(n29129,n28345,n28971);
  nand U30974(n29127,n28972,n28734);
  nand U30975(n29126,n28973,G59315);
  nand U30976(n29125,n28974,n28348);
  nand U30977(G2550,n29132,n29133,n29134,n29135);
  nor U30978(n29135,n29136,n29137);
  nor U30979(n29137,n29138,n28970);
  nor U30980(n29136,n28356,n28971);
  nand U30981(n29134,n28972,n28359);
  nand U30982(n29133,n28973,G59314);
  nand U30983(n29132,n28974,n28360);
  nand U30984(G2549,n29139,n29140,n29141,n29142);
  nor U30985(n29142,n29143,n29144);
  nor U30986(n29144,n29145,n28970);
  nor U30987(n29143,n28369,n28971);
  nand U30988(n29141,n28972,n28371);
  nand U30989(n29140,n28973,G59313);
  nand U30990(n29139,n28974,n27871);
  nand U30991(G2548,n29146,n29147,n29148,n29149);
  nor U30992(n29149,n29150,n29151);
  nor U30993(n29151,n28379,n28970);
  nor U30994(n29150,n29152,n28971);
  nand U30995(n29148,n28972,n28384);
  nand U30996(n29147,n28973,G59312);
  nand U30997(n29146,n28974,n27881);
  nand U30998(G2547,n29153,n29154,n29155,n29156);
  nor U30999(n29156,n29157,n29158);
  nor U31000(n29158,n28392,n28970);
  nor U31001(n29157,n29159,n28971);
  nand U31002(n29155,n28972,n28396);
  nand U31003(n29154,n28973,G59311);
  nand U31004(n29153,n28974,n27891);
  nand U31005(G2546,n29160,n29161,n29162,n29163);
  nor U31006(n29163,n29164,n29165);
  nor U31007(n29165,n28404,n28970);
  nor U31008(n29164,n29166,n28971);
  not U31009(n28971,n29106);
  nand U31010(n29162,n28972,n28407);
  nand U31011(n29161,n28973,G59310);
  nand U31012(n29160,n28974,n27900);
  nand U31013(G2545,n29167,n29168,n29169,n29170);
  nand U31014(n29170,n28972,n28431);
  nor U31015(n29169,n29171,n29172);
  nor U31016(n29172,n28417,n29103);
  not U31017(n29103,n28974);
  nor U31018(n29171,n28013,n29105);
  not U31019(n29105,n28973);
  nand U31020(n29168,n29106,n27969);
  nor U31021(n29106,n29174,n29047);
  nand U31022(n29167,n29047,G59150);
  not U31023(n29047,n28970);
  nand U31024(n28970,n28001,n27927);
  nand U31025(n27927,n27928,n28416,n29175);
  or U31026(n28001,n27991,n27990);
  nand U31027(n27991,n29176,G58977,n29177);
  nand U31028(G2544,n29178,n29179,n29180,n29181);
  nor U31029(n29181,n29182,n29183,n29184);
  nor U31030(n29184,G59149,n29185,n29186);
  nor U31031(n29183,n29187,n29188);
  nor U31032(n29187,n29189,n29190);
  nor U31033(n29189,n29191,n29185);
  nor U31034(n29182,n28061,n29192);
  nand U31035(n29180,n29193,n28063);
  nand U31036(n29179,n29194,n28066);
  nand U31037(n28066,n29195,n29196);
  nand U31038(n29196,n29197,n29198);
  nand U31039(n29198,n29199,n29200);
  nand U31040(n29199,n29201,n29202,n29203);
  nand U31041(n29195,n29204,n29200,n29205);
  nand U31042(n29200,n29206,n29207,n29208);
  nand U31043(n29206,n29209,n29205);
  nand U31044(n29204,n29203,n29209);
  not U31045(n29203,n29207);
  nand U31046(n29207,n29210,n29211,n29212,n29213);
  nand U31047(n29213,n28060,n29214);
  nand U31048(n29212,n29197,n28063);
  not U31049(n28063,n28430);
  xor U31050(n28430,n29215,n29216);
  nand U31051(n29215,n29217,n29218);
  nand U31052(n29218,n29219,n27993);
  nand U31053(n29217,n29220,n28963);
  nand U31054(n29220,n29221,n29222,n29219);
  and U31055(n29219,n29223,n29224);
  nand U31056(n29224,G59308,n29225);
  nand U31057(n29223,G59181,n29226);
  nand U31058(n29222,G59149,n29227);
  nand U31059(n29221,G59276,n29228);
  nand U31060(n29211,G59149,n29229);
  nand U31061(n29210,n29230,G59340);
  nand U31062(n29178,n29231,n28060);
  xor U31063(n28060,n29232,n29233);
  nor U31064(n29233,n29234,n29235,n29236);
  nor U31065(n29236,n29173,n28057);
  not U31066(n28057,G59181);
  nor U31067(n29235,n29237,n29188);
  nor U31068(n29234,n28963,n28061);
  not U31069(n28061,G59340);
  nand U31070(G2543,n29238,n29239,n29240,n29241);
  nor U31071(n29241,n29242,n29243,n29244);
  nor U31072(n29244,n28078,n29192);
  nor U31073(n29243,n29245,n29185);
  nor U31074(n29242,n29246,n29247);
  nand U31075(n29240,n29193,n28079);
  nand U31076(n29239,n29194,n28080);
  nand U31077(n28080,n29248,n29249);
  nand U31078(n29249,n29197,n29250);
  nand U31079(n29250,n29209,n29208);
  nand U31080(n29208,n29201,n29202);
  not U31081(n29201,n29251);
  nand U31082(n29209,n29251,n29252);
  nand U31083(n29248,n29253,n29205);
  xnor U31084(n29253,n29251,n29202);
  not U31085(n29202,n29252);
  nand U31086(n29252,n29254,n29255,n29256,n29257);
  nor U31087(n29257,n29258,n29259);
  nor U31088(n29259,n28078,n29260);
  nor U31089(n29258,n29261,n29246);
  nand U31090(n29256,n29197,n28079);
  nand U31091(n29255,n29262,n29263,n29264);
  nand U31092(n29263,n28457,n29265);
  nand U31093(n29262,n29266,n28077);
  nand U31094(n29266,n29267,n29265);
  nor U31095(n29265,n28089,n28101);
  nand U31096(n29254,n28457,n29268);
  nand U31097(n29251,n29269,n29270);
  nand U31098(n29270,n29197,n29271);
  nand U31099(n29271,n29272,n29273);
  or U31100(n29269,n29273,n29272);
  nand U31101(n29238,n29231,n28457);
  not U31102(n28457,n28077);
  nand U31103(n28077,n29274,n29232);
  nand U31104(n29232,n29275,n29276,n29277);
  xnor U31105(n29277,n29278,n29174);
  nand U31106(n29274,n29279,n29280);
  nand U31107(n29280,n29276,n29275);
  xnor U31108(n29279,n29226,n29278);
  nand U31109(n29278,n29281,n29282,n29283,n29284);
  nor U31110(n29284,n29285,n29286);
  nor U31111(n29286,n29173,n28075);
  not U31112(n28075,G59180);
  nor U31113(n29285,n28963,n28078);
  not U31114(n28078,G59339);
  nand U31115(n29283,G59148,n29287);
  nand U31116(n29282,n28079,n29288);
  not U31117(n28079,n28592);
  nand U31118(n28592,n29216,n29289);
  nand U31119(n29289,n29290,n29291);
  or U31120(n29216,n29291,n29290);
  xor U31121(n29290,n29292,n28963);
  nand U31122(n29292,n29293,n29294,n29295,n29296);
  nor U31123(n29296,n29297,n29298);
  and U31124(n29298,n29225,G59307);
  and U31125(n29297,n29228,G59275);
  nand U31126(n29295,G59180,n29226);
  or U31127(n29294,n29245,n27999);
  nand U31128(n29245,n29186,n29299);
  nand U31129(n29299,n29300,n29301);
  not U31130(n29186,n29191);
  nor U31131(n29191,n29301,n29300);
  nand U31132(n29300,n29302,n29303);
  nand U31133(n29303,n27943,n29246);
  not U31134(n29246,G59148);
  nand U31135(n29302,n29304,n29305,n29306,n28689);
  nor U31136(n29306,n29307,n29308);
  nand U31137(n29308,n29309,n29310,n29311,n29312);
  nand U31138(n29312,n29313,G59100);
  nand U31139(n29311,n29314,G59092);
  nand U31140(n29310,n29315,G59084);
  nand U31141(n29309,n29316,G59076);
  nand U31142(n29307,n29317,n29318,n29319,n29320);
  nand U31143(n29320,n29321,G59068);
  nand U31144(n29319,n29322,G59060);
  nand U31145(n29318,n29323,G59052);
  nand U31146(n29317,n29324,G59044);
  nor U31147(n29305,n29325,n29326,n29327,n29328);
  nor U31148(n29328,n29329,n29330);
  nor U31149(n29327,n29331,n29332);
  nor U31150(n29326,n29333,n29334);
  nor U31151(n29325,n29335,n29336);
  nor U31152(n29304,n29337,n29338,n29339,n29340);
  nor U31153(n29340,n29341,n29342);
  nor U31154(n29339,n29343,n29344);
  nor U31155(n29338,n29345,n29346);
  nor U31156(n29337,n29347,n29348);
  nand U31157(n29293,G59148,n29227);
  nand U31158(n29281,n29349,n29350);
  nand U31159(G2542,n29351,n29352,n29353,n29354);
  nor U31160(n29354,n29355,n29356,n29357);
  nor U31161(n29357,n28090,n29192);
  nor U31162(n29356,n29358,n29185);
  nor U31163(n29355,n29359,n29247);
  nand U31164(n29353,n29193,n28091);
  nand U31165(n29352,n29194,n28092);
  xnor U31166(n28092,n29272,n29360);
  xnor U31167(n29360,n29197,n29273);
  nand U31168(n29273,n29361,n29362);
  nand U31169(n29362,n29363,n29205);
  nand U31170(n29363,n29364,n29365);
  or U31171(n29361,n29364,n29365);
  and U31172(n29272,n29366,n29367,n29368,n29369);
  nor U31173(n29369,n29370,n29371);
  nor U31174(n29371,n28090,n29260);
  nor U31175(n29370,n29261,n29359);
  not U31176(n29359,G59147);
  nand U31177(n29368,n29197,n28091);
  nand U31178(n29367,n29372,n29373,n29264);
  nand U31179(n29373,n28101,n28089);
  nand U31180(n29372,n28465,n29374);
  nand U31181(n29374,n29267,n28089);
  nand U31182(n29366,n28461,n29268);
  nand U31183(n29351,n29231,n28461);
  not U31184(n28461,n28089);
  xnor U31185(n28089,n29275,n29276);
  nor U31186(n29276,n29375,n29376);
  xnor U31187(n29275,n29377,n29174);
  nand U31188(n29377,n29378,n29379,n29380,n29381);
  nor U31189(n29381,n29382,n29383);
  nor U31190(n29383,n29173,n28088);
  nor U31191(n29382,n28963,n28090);
  not U31192(n28090,G59338);
  nand U31193(n29380,G59147,n29287);
  nand U31194(n29379,n28091,n29288);
  not U31195(n28091,n28601);
  nand U31196(n28601,n29291,n29384);
  nand U31197(n29384,n29385,n29386);
  or U31198(n29291,n29386,n29385);
  xor U31199(n29385,n27993,n29387);
  nor U31200(n29387,n29388,n29389,n29390,n29391);
  and U31201(n29391,n29225,G59306);
  nor U31202(n29390,n27999,n29358);
  nand U31203(n29358,n29392,n29301);
  nand U31204(n29301,n29393,n29394);
  or U31205(n29392,n29394,n29393);
  nand U31206(n29394,n29395,n29396);
  nand U31207(n29396,G59147,n27943);
  nand U31208(n29395,n29397,n28689);
  nand U31209(n29397,n29398,n29399,n29400,n29401);
  nor U31210(n29401,n29402,n29403,n29404,n29405);
  nor U31211(n29405,n29406,n29330);
  nor U31212(n29404,n29407,n29332);
  nor U31213(n29403,n29408,n29334);
  nor U31214(n29402,n29409,n29336);
  nor U31215(n29400,n29410,n29411,n29412,n29413);
  nor U31216(n29413,n29414,n29342);
  nor U31217(n29412,n29415,n29344);
  nor U31218(n29411,n29416,n29346);
  nor U31219(n29410,n29417,n29348);
  nor U31220(n29399,n29418,n29419,n29420,n29421);
  nor U31221(n29421,n29422,n29423);
  nor U31222(n29420,n29424,n29425);
  nor U31223(n29419,n29426,n29427);
  nor U31224(n29418,n29428,n29429);
  nor U31225(n29398,n29430,n29431,n29432,n29433);
  nor U31226(n29433,n29434,n29435);
  nor U31227(n29432,n29436,n29437);
  nor U31228(n29431,n29438,n29439);
  nor U31229(n29430,n29440,n29441);
  nor U31230(n29389,n29174,n28088);
  not U31231(n28088,G59179);
  nand U31232(n29388,n29442,n29443);
  nand U31233(n29443,G59147,n29227);
  nand U31234(n29442,G59274,n29228);
  nand U31235(n29378,n29349,n29444);
  nand U31236(G2541,n29445,n29446,n29447,n29448);
  nor U31237(n29448,n29449,n29450,n29451);
  nor U31238(n29451,n28102,n29192);
  nor U31239(n29450,n29452,n29185);
  nor U31240(n29449,n29453,n29247);
  nand U31241(n29447,n29193,n28103);
  nand U31242(n29446,n29194,n28104);
  xor U31243(n28104,n29454,n29365);
  nand U31244(n29365,n29455,n29456,n29457,n29458);
  nor U31245(n29458,n29459,n29460);
  nor U31246(n29460,n29261,n29453);
  nor U31247(n29459,n28608,n29205);
  nand U31248(n29457,n29230,G59337);
  nand U31249(n29456,n28465,n29268);
  nand U31250(n29455,n29267,n29264,n28101);
  xnor U31251(n29454,n29205,n29364);
  nand U31252(n29364,n29461,n29462);
  nand U31253(n29462,n29197,n29463);
  or U31254(n29463,n29464,n29465);
  nand U31255(n29461,n29465,n29464);
  nand U31256(n29445,n29231,n28465);
  not U31257(n28465,n28101);
  xnor U31258(n28101,n29375,n29376);
  xor U31259(n29376,n29466,n29174);
  nand U31260(n29466,n29467,n29468,n29469,n29470);
  nor U31261(n29470,n29471,n29472);
  nor U31262(n29472,n29173,n28100);
  not U31263(n28100,G59178);
  nor U31264(n29471,n28963,n28102);
  not U31265(n28102,G59337);
  nand U31266(n29469,G59146,n29287);
  nand U31267(n29468,n28103,n29288);
  not U31268(n28103,n28608);
  nand U31269(n28608,n29386,n29473);
  nand U31270(n29473,n29474,n29475);
  nand U31271(n29475,n29476,n29477);
  nand U31272(n29386,n29477,n29476,n29478);
  not U31273(n29478,n29474);
  xor U31274(n29474,n29479,n28963);
  nand U31275(n29479,n29480,n29481,n29482,n29483);
  nor U31276(n29483,n29484,n29485);
  and U31277(n29485,n29228,G59273);
  nor U31278(n29484,n29486,n29453);
  nand U31279(n29482,G59178,n29226);
  or U31280(n29481,n29452,n27999);
  nand U31281(n29452,n29487,n29488);
  nand U31282(n29488,n29489,n29490);
  not U31283(n29487,n29393);
  nor U31284(n29393,n29490,n29489);
  nand U31285(n29489,n29491,n29492);
  nand U31286(n29492,n27943,n29453);
  not U31287(n29453,G59146);
  nand U31288(n29491,n29493,n29494,n29495,n28689);
  nor U31289(n29495,n29496,n29497);
  nand U31290(n29497,n29498,n29499,n29500,n29501);
  nand U31291(n29501,n29313,G59102);
  nand U31292(n29500,n29314,G59094);
  nand U31293(n29499,n29315,G59086);
  nand U31294(n29498,n29316,G59078);
  nand U31295(n29496,n29502,n29503,n29504,n29505);
  nand U31296(n29505,n29321,G59070);
  nand U31297(n29504,n29322,G59062);
  nand U31298(n29503,n29323,G59054);
  nand U31299(n29502,n29324,G59046);
  nor U31300(n29494,n29506,n29507,n29508,n29509);
  nor U31301(n29509,n29510,n29330);
  nor U31302(n29508,n29511,n29332);
  nor U31303(n29507,n29512,n29334);
  nor U31304(n29506,n29513,n29336);
  nor U31305(n29493,n29514,n29515,n29516,n29517);
  nor U31306(n29517,n29518,n29342);
  nor U31307(n29516,n29519,n29344);
  nor U31308(n29515,n29520,n29346);
  nor U31309(n29514,n29521,n29348);
  nand U31310(n29480,G59305,n29225);
  nand U31311(n29467,n29349,n29522);
  nand U31312(G2540,n29523,n29524,n29525,n29526);
  nor U31313(n29526,n29527,n29528,n29529);
  nor U31314(n29529,n28114,n29192);
  nor U31315(n29528,n29530,n29185);
  nor U31316(n29527,n29531,n29247);
  nand U31317(n29525,n29193,n28115);
  nand U31318(n29524,n29194,n28116);
  xor U31319(n28116,n29532,n29465);
  nand U31320(n29465,n29533,n29534,n29535,n29536);
  nor U31321(n29536,n29537,n29538);
  nor U31322(n29538,n28114,n29260);
  nor U31323(n29537,n29261,n29531);
  nand U31324(n29535,n29197,n28115);
  nand U31325(n29534,n28473,n29539,n29264,n29540);
  nand U31326(n29533,n28469,n29268);
  nand U31327(n29268,n29541,n29542);
  nand U31328(n29542,n29264,n29540);
  not U31329(n29540,n29267);
  nor U31330(n29267,n28125,n29543,n28113);
  xnor U31331(n29532,n29205,n29464);
  nand U31332(n29464,n29544,n29545);
  nand U31333(n29545,n29197,n29546);
  or U31334(n29546,n29547,n29548);
  nand U31335(n29544,n29548,n29547);
  nand U31336(n29523,n29231,n28469);
  not U31337(n28469,n28113);
  nand U31338(n28113,n29549,n29375);
  or U31339(n29375,n29550,n29551);
  nand U31340(n29549,n29551,n29550);
  or U31341(n29550,n29552,n29553,n29554);
  xor U31342(n29551,n29555,n29174);
  nand U31343(n29555,n29556,n29557,n29558,n29559);
  nor U31344(n29559,n29560,n29561);
  nor U31345(n29561,n29173,n28112);
  nor U31346(n29560,n28963,n28114);
  not U31347(n28114,G59336);
  nand U31348(n29558,G59145,n29287);
  nand U31349(n29557,n28115,n29288);
  xor U31350(n28115,n29476,n29477);
  xnor U31351(n29477,n27993,n29562);
  nor U31352(n29562,n29563,n29564,n29565,n29566);
  and U31353(n29566,n29225,G59304);
  nor U31354(n29565,n27999,n29530);
  nand U31355(n29530,n29490,n29567);
  nand U31356(n29567,n29568,n29569);
  or U31357(n29490,n29569,n29568);
  nand U31358(n29568,n29570,n29571);
  nand U31359(n29571,n27943,n29531);
  not U31360(n29531,G59145);
  nand U31361(n29570,n29572,n29573,n29574,n28689);
  nor U31362(n29574,n29575,n29576);
  nand U31363(n29576,n29577,n29578,n29579,n29580);
  nand U31364(n29580,n29313,G59103);
  nand U31365(n29579,n29314,G59095);
  nand U31366(n29578,n29315,G59087);
  nand U31367(n29577,n29316,G59079);
  nand U31368(n29575,n29581,n29582,n29583,n29584);
  nand U31369(n29584,n29321,G59071);
  nand U31370(n29583,n29322,G59063);
  nand U31371(n29582,n29323,G59055);
  nand U31372(n29581,n29324,G59047);
  nor U31373(n29573,n29585,n29586,n29587,n29588);
  nor U31374(n29588,n29589,n29330);
  nor U31375(n29587,n29590,n29332);
  nor U31376(n29586,n29591,n29334);
  nor U31377(n29585,n29592,n29336);
  nor U31378(n29572,n29593,n29594,n29595,n29596);
  nor U31379(n29596,n29597,n29342);
  nor U31380(n29595,n29598,n29344);
  nor U31381(n29594,n29599,n29346);
  nor U31382(n29593,n29600,n29348);
  nor U31383(n29564,n29174,n28112);
  not U31384(n28112,G59177);
  nand U31385(n29563,n29601,n29602);
  nand U31386(n29602,G59145,n29227);
  nand U31387(n29601,G59272,n29228);
  and U31388(n29476,n29603,n29604);
  nand U31389(n29556,n29349,n29605);
  nand U31390(G2539,n29606,n29607,n29608,n29609);
  nor U31391(n29609,n29610,n29611,n29612);
  nor U31392(n29612,n28126,n29192);
  nor U31393(n29611,n29613,n29185);
  nor U31394(n29610,n29614,n29247);
  nand U31395(n29608,n29193,n28127);
  nand U31396(n29607,n29194,n28128);
  xor U31397(n28128,n29615,n29548);
  nand U31398(n29548,n29616,n29617,n29618,n29619);
  nor U31399(n29619,n29620,n29621);
  nor U31400(n29621,n29261,n29614);
  nor U31401(n29620,n28622,n29205);
  nand U31402(n29618,n29230,G59335);
  nand U31403(n29617,n28473,n29622);
  nand U31404(n29616,n29539,n29264,n28125);
  not U31405(n29539,n29543);
  xnor U31406(n29615,n29205,n29547);
  nand U31407(n29547,n29623,n29624);
  nand U31408(n29624,n29197,n29625);
  or U31409(n29625,n29626,n29627);
  nand U31410(n29623,n29627,n29626);
  nand U31411(n29606,n29231,n28473);
  not U31412(n28473,n28125);
  xor U31413(n28125,n29553,n29628);
  nor U31414(n29628,n29552,n29554);
  xnor U31415(n29553,n29629,n29226);
  nand U31416(n29629,n29630,n29631,n29632,n29633);
  nor U31417(n29633,n29634,n29635);
  nor U31418(n29635,n29173,n28124);
  not U31419(n28124,G59176);
  nor U31420(n29634,n28963,n28126);
  not U31421(n28126,G59335);
  nand U31422(n29632,G59144,n29287);
  nand U31423(n29631,n28127,n29288);
  not U31424(n28127,n28622);
  xnor U31425(n28622,n29604,n29603);
  xnor U31426(n29604,n29636,n28963);
  nand U31427(n29636,n29637,n29638,n29639,n29640);
  nor U31428(n29640,n29641,n29642);
  and U31429(n29642,n29228,G59271);
  nor U31430(n29641,n29486,n29614);
  nand U31431(n29639,G59176,n29226);
  or U31432(n29638,n29613,n27999);
  nand U31433(n29613,n29569,n29643);
  nand U31434(n29643,n29644,n29645);
  or U31435(n29569,n29645,n29644);
  nand U31436(n29644,n29646,n29647);
  nand U31437(n29647,n27943,n29614);
  not U31438(n29614,G59144);
  nand U31439(n29646,n29648,n29649,n29650,n28689);
  nor U31440(n29650,n29651,n29652);
  nand U31441(n29652,n29653,n29654,n29655,n29656);
  nand U31442(n29656,n29313,G59104);
  not U31443(n29313,n29441);
  nand U31444(n29655,n29314,G59096);
  not U31445(n29314,n29439);
  nand U31446(n29654,n29315,G59088);
  not U31447(n29315,n29437);
  nand U31448(n29653,n29316,G59080);
  not U31449(n29316,n29435);
  nand U31450(n29651,n29657,n29658,n29659,n29660);
  nand U31451(n29660,n29321,G59072);
  not U31452(n29321,n29429);
  nand U31453(n29659,n29322,G59064);
  not U31454(n29322,n29427);
  nand U31455(n29658,n29323,G59056);
  not U31456(n29323,n29425);
  nand U31457(n29657,n29324,G59048);
  not U31458(n29324,n29423);
  nor U31459(n29649,n29661,n29662,n29663,n29664);
  nor U31460(n29664,n29665,n29330);
  nor U31461(n29663,n29666,n29332);
  nor U31462(n29662,n29667,n29334);
  nor U31463(n29661,n29668,n29336);
  nor U31464(n29648,n29669,n29670,n29671,n29672);
  nor U31465(n29672,n29673,n29342);
  nor U31466(n29671,n29674,n29344);
  nor U31467(n29670,n29675,n29346);
  nor U31468(n29669,n29676,n29348);
  nand U31469(n29637,G59303,n29225);
  nand U31470(n29630,n29349,n29677);
  nand U31471(G2538,n29678,n29679,n29680,n29681);
  nor U31472(n29681,n29682,n29683,n29684);
  nor U31473(n29684,n28138,n29192);
  nor U31474(n29683,n28629,n29685);
  not U31475(n28629,n28139);
  nor U31476(n29682,n29686,n29247);
  nand U31477(n29680,n29231,n28137);
  nand U31478(n29679,n29687,n29645,n29688);
  nand U31479(n29678,n29194,n28140);
  xor U31480(n28140,n29689,n29627);
  nand U31481(n29627,n29690,n29691,n29692,n29693);
  nor U31482(n29693,n29694,n29695);
  nor U31483(n29695,n28138,n29260);
  nor U31484(n29694,n29261,n29686);
  nand U31485(n29692,n29197,n28139);
  nand U31486(n29691,n28480,n29543,n29696);
  nand U31487(n29690,n28137,n29622);
  nand U31488(n29622,n29541,n29697);
  nand U31489(n29697,n29264,n29543);
  nand U31490(n29543,n29698,n28480,n28137,n28484);
  xor U31491(n28137,n29554,n29552);
  xor U31492(n29552,n29699,n29174);
  nand U31493(n29699,n29700,n29701,n29702,n29703);
  nor U31494(n29703,n29704,n29705);
  nor U31495(n29705,n29173,n28136);
  not U31496(n28136,G59175);
  nor U31497(n29704,n28963,n28138);
  not U31498(n28138,G59334);
  nand U31499(n29702,G59143,n29287);
  nand U31500(n29701,n28139,n29288);
  nor U31501(n28139,n29706,n29603);
  nor U31502(n29603,n29707,n29708);
  and U31503(n29706,n29708,n29707);
  nand U31504(n29707,n29709,n29710,n29711);
  xor U31505(n29708,n29712,n28963);
  nand U31506(n29712,n29713,n29714,n29715,n29716);
  nor U31507(n29716,n29717,n29718);
  and U31508(n29718,n29228,G59270);
  nor U31509(n29717,n29486,n29686);
  nand U31510(n29715,G59175,n29226);
  nand U31511(n29714,n29687,n29645,n28576);
  nand U31512(n29645,n29719,n29720,n29721);
  nand U31513(n29720,n27943,n29686);
  not U31514(n29686,G59143);
  or U31515(n29719,n29722,n27943);
  nand U31516(n29687,n29723,n29724,n29725);
  nand U31517(n29724,G59143,n27943);
  nand U31518(n29723,n29722,n28689);
  nand U31519(n29722,n29726,n29727,n29728,n29729);
  nor U31520(n29729,n29730,n29731,n29732,n29733);
  nor U31521(n29733,n29734,n29330);
  nor U31522(n29732,n29735,n29332);
  nor U31523(n29731,n29736,n29334);
  nor U31524(n29730,n29737,n29336);
  nor U31525(n29728,n29738,n29739,n29740,n29741);
  nor U31526(n29741,n29742,n29342);
  nor U31527(n29740,n29743,n29344);
  nor U31528(n29739,n29744,n29346);
  nor U31529(n29738,n29745,n29348);
  nor U31530(n29727,n29746,n29747,n29748,n29749);
  nor U31531(n29749,n29750,n29423);
  nor U31532(n29748,n29751,n29425);
  nor U31533(n29747,n29752,n29427);
  nor U31534(n29746,n29753,n29429);
  nor U31535(n29726,n29754,n29755,n29756,n29757);
  nor U31536(n29757,n29758,n29435);
  nor U31537(n29756,n29759,n29437);
  nor U31538(n29755,n29760,n29439);
  nor U31539(n29754,n29761,n29441);
  nand U31540(n29713,G59302,n29225);
  nand U31541(n29700,n29349,n29762);
  xnor U31542(n29689,n29205,n29626);
  nand U31543(n29626,n29763,n29764);
  nand U31544(n29764,n29197,n29765);
  or U31545(n29765,n29766,n29767);
  nand U31546(n29763,n29767,n29766);
  nand U31547(G2537,n29768,n29769,n29770,n29771);
  nor U31548(n29771,n29772,n29773,n29774);
  nor U31549(n29774,n28150,n29192);
  nor U31550(n29773,n29775,n29185);
  nor U31551(n29772,n29776,n29247);
  nand U31552(n29770,n29193,n28151);
  nand U31553(n29769,n29194,n28152);
  xor U31554(n28152,n29777,n29767);
  nand U31555(n29767,n29778,n29779,n29780,n29781);
  nor U31556(n29781,n29782,n29783);
  nor U31557(n29783,n29261,n29776);
  nor U31558(n29782,n28636,n29205);
  not U31559(n28636,n28151);
  nand U31560(n29780,n29230,G59333);
  nand U31561(n29779,n29696,n28149);
  nor U31562(n29696,n28161,n28761,n29784);
  nand U31563(n29778,n28480,n29785);
  nand U31564(n29785,n29786,n29787);
  nand U31565(n29787,n29264,n28161);
  not U31566(n29786,n29788);
  xnor U31567(n29777,n29205,n29766);
  nand U31568(n29766,n29789,n29790);
  nand U31569(n29790,n29197,n29791);
  or U31570(n29791,n29792,n29793);
  nand U31571(n29789,n29793,n29792);
  nand U31572(n29768,n29231,n28480);
  not U31573(n28480,n28149);
  nand U31574(n28149,n29554,n29794);
  nand U31575(n29794,n29795,n29796);
  or U31576(n29554,n29796,n29795);
  and U31577(n29795,n29797,n29798);
  nand U31578(n29797,n29799,n29800);
  xor U31579(n29796,n29801,n29174);
  nand U31580(n29801,n29802,n29803,n29804,n29805);
  nor U31581(n29805,n29806,n29807);
  nor U31582(n29807,n29173,n28148);
  not U31583(n28148,G59174);
  nor U31584(n29806,n28963,n28150);
  not U31585(n28150,G59333);
  nand U31586(n29804,G59142,n29287);
  nand U31587(n29803,n28151,n29288);
  xnor U31588(n28151,n29808,n29711);
  xor U31589(n29711,n29809,n27993);
  nand U31590(n29809,n29810,n29811,n29812,n29813);
  nor U31591(n29813,n29814,n29815);
  and U31592(n29815,n29228,G59269);
  nor U31593(n29814,n29486,n29776);
  not U31594(n29776,G59142);
  nand U31595(n29812,G59174,n29226);
  or U31596(n29811,n29775,n27999);
  nand U31597(n29775,n29725,n29816);
  nand U31598(n29816,n29817,n29818);
  not U31599(n29725,n29721);
  nor U31600(n29721,n29818,n29817);
  and U31601(n29817,n29819,n29820);
  nand U31602(n29820,G59142,n27943);
  nand U31603(n29819,n29821,n28689);
  nand U31604(n29821,n29822,n29823,n29824,n29825);
  nor U31605(n29825,n29826,n29827,n29828,n29829);
  nor U31606(n29829,n29830,n29330);
  nor U31607(n29828,n29831,n29332);
  nor U31608(n29827,n29832,n29334);
  nor U31609(n29826,n29833,n29336);
  nor U31610(n29824,n29834,n29835,n29836,n29837);
  nor U31611(n29837,n29838,n29342);
  nor U31612(n29836,n29839,n29344);
  nor U31613(n29835,n29840,n29346);
  nor U31614(n29834,n29841,n29348);
  nor U31615(n29823,n29842,n29843,n29844,n29845);
  nor U31616(n29845,n29846,n29423);
  nor U31617(n29844,n29847,n29425);
  nor U31618(n29843,n29848,n29427);
  nor U31619(n29842,n29849,n29429);
  nor U31620(n29822,n29850,n29851,n29852,n29853);
  nor U31621(n29853,n29854,n29435);
  nor U31622(n29852,n29855,n29437);
  nor U31623(n29851,n29856,n29439);
  nor U31624(n29850,n29857,n29441);
  nand U31625(n29818,n29858,n29859);
  nand U31626(n29810,G59301,n29225);
  nand U31627(n29808,n29710,n29709);
  nand U31628(n29802,n29349,n29860);
  nand U31629(G2536,n29861,n29862,n29863,n29864);
  nor U31630(n29864,n29865,n29866,n29867);
  nor U31631(n29867,n28162,n29192);
  nor U31632(n29866,n28643,n29685);
  nor U31633(n29865,n29868,n29247);
  nand U31634(n29863,n29231,n28484);
  nand U31635(n29862,n29688,n29869);
  nand U31636(n29861,n29194,n28164);
  xor U31637(n28164,n29870,n29793);
  nand U31638(n29793,n29871,n29872,n29873,n29874);
  nor U31639(n29874,n29875,n29876);
  nor U31640(n29876,n29261,n29868);
  nor U31641(n29875,n28643,n29205);
  not U31642(n28643,n28163);
  nand U31643(n29873,n29230,G59332);
  nand U31644(n29872,n28484,n29788);
  not U31645(n28484,n28161);
  nand U31646(n29871,n29698,n29264,n28161);
  xnor U31647(n28161,n29799,n29877);
  and U31648(n29877,n29798,n29800);
  nand U31649(n29800,n29878,n29879,n29880);
  nand U31650(n29880,n29349,n29881);
  nand U31651(n29798,n29882,n29881,n29349);
  nand U31652(n29882,n29878,n29879);
  or U31653(n29879,n29883,n29174);
  nand U31654(n29878,n29174,n29883);
  nand U31655(n29883,n29884,n29885,n29886,n29887);
  nor U31656(n29887,n29888,n29889);
  nor U31657(n29889,n29173,n28160);
  not U31658(n28160,G59173);
  nor U31659(n29888,n28963,n28162);
  not U31660(n28162,G59332);
  nand U31661(n29886,G59141,n29287);
  nand U31662(n29885,n28163,n29288);
  xor U31663(n28163,n29709,n29710);
  xnor U31664(n29709,n29890,n28963);
  nand U31665(n29890,n29891,n29892,n29893,n29894);
  nor U31666(n29894,n29895,n29896);
  and U31667(n29896,n29228,G59268);
  nor U31668(n29895,n29486,n29868);
  not U31669(n29868,G59141);
  nand U31670(n29893,G59173,n29226);
  nand U31671(n29892,n28576,n29869);
  xor U31672(n29869,n29858,n29859);
  nand U31673(n29859,n29897,n29898);
  nand U31674(n29898,G59141,n27943);
  nand U31675(n29897,n29899,n28689);
  nand U31676(n29899,n29900,n29901,n29902,n29903);
  nor U31677(n29903,n29904,n29905,n29906,n29907);
  nor U31678(n29907,n29908,n29330);
  nand U31679(n29330,n29909,n29910);
  nor U31680(n29906,n29911,n29332);
  nand U31681(n29332,n29912,n29910);
  nor U31682(n29905,n29913,n29334);
  nand U31683(n29334,n29914,n29910);
  nor U31684(n29904,n29915,n29336);
  nand U31685(n29336,n29916,n29910);
  and U31686(n29910,n29917,n29918);
  nor U31687(n29902,n29919,n29920,n29921,n29922);
  nor U31688(n29922,n29923,n29342);
  nand U31689(n29342,n29924,n29909);
  nor U31690(n29921,n29925,n29344);
  nand U31691(n29344,n29924,n29912);
  nor U31692(n29920,n29926,n29346);
  nand U31693(n29346,n29924,n29914);
  nor U31694(n29919,n29927,n29348);
  nand U31695(n29348,n29924,n29916);
  and U31696(n29924,n29928,n29918);
  nor U31697(n29901,n29929,n29930,n29931,n29932);
  nor U31698(n29932,n29933,n29423);
  nand U31699(n29423,n29934,n29909);
  nor U31700(n29931,n29935,n29425);
  nand U31701(n29425,n29934,n29912);
  nor U31702(n29930,n29936,n29427);
  nand U31703(n29427,n29934,n29914);
  nor U31704(n29929,n29937,n29429);
  nand U31705(n29429,n29934,n29916);
  nor U31706(n29934,n29918,n29928);
  not U31707(n29928,n29917);
  nor U31708(n29900,n29938,n29939,n29940,n29941);
  nor U31709(n29941,n29942,n29435);
  nand U31710(n29435,n29943,n29909);
  nor U31711(n29909,n29944,n29945);
  nor U31712(n29940,n29946,n29437);
  nand U31713(n29437,n29943,n29912);
  nor U31714(n29912,G59112,n29945);
  nor U31715(n29939,n29947,n29439);
  nand U31716(n29439,n29943,n29914);
  nor U31717(n29914,n29948,n29944);
  nor U31718(n29938,n29949,n29441);
  nand U31719(n29441,n29943,n29916);
  nor U31720(n29916,n29948,G59112);
  nor U31721(n29943,n29918,n29917);
  nand U31722(n29858,n29950,n29951);
  nand U31723(n29951,n29952,G59140);
  nand U31724(n29950,n29350,n28689);
  nand U31725(n29350,n29953,n29954,n29955,n29956);
  nor U31726(n29956,n29957,n29958,n29959,n29960);
  nor U31727(n29960,n29961,n29962);
  nor U31728(n29959,n29963,n29964);
  nor U31729(n29958,n29965,n29966);
  nor U31730(n29957,n29967,n29968);
  nor U31731(n29955,n29969,n29970,n29971,n29972);
  nor U31732(n29972,n29973,n29974);
  nor U31733(n29971,n29975,n29976);
  nor U31734(n29970,n29977,n29978);
  nor U31735(n29969,n29979,n29980);
  nor U31736(n29954,n29981,n29982,n29983,n29984);
  nor U31737(n29984,n29341,n29985);
  nor U31738(n29983,n29343,n29986);
  nor U31739(n29982,n29345,n29987);
  nor U31740(n29981,n29347,n29988);
  nor U31741(n29953,n29989,n29990,n29991,n29992);
  nor U31742(n29992,n29329,n29993);
  nor U31743(n29991,n29331,n29994);
  nor U31744(n29990,n29333,n29995);
  nor U31745(n29989,n29335,n29996);
  nand U31746(n29891,G59300,n29225);
  nand U31747(n29884,n29349,n29997);
  nand U31748(n29799,n29998,n29999);
  nand U31749(n29999,n30000,n30001);
  not U31750(n29698,n29784);
  xnor U31751(n29870,n29205,n29792);
  nand U31752(n29792,n30002,n30003);
  nand U31753(n30003,n29197,n30004);
  or U31754(n30004,n30005,n30006);
  nand U31755(n30002,n30006,n30005);
  nand U31756(G2535,n30007,n30008,n30009,n30010);
  nor U31757(n30010,n30011,n30012,n30013);
  nor U31758(n30013,n28174,n29192);
  and U31759(n30012,n30014,n29688);
  nor U31760(n30011,n30015,n29247);
  nand U31761(n30009,n29193,n28175);
  nand U31762(n30008,n29194,n28176);
  xor U31763(n28176,n30016,n30006);
  nand U31764(n30006,n30017,n30018,n30019,n30020);
  nor U31765(n30020,n30021,n30022);
  nor U31766(n30022,n28174,n29260);
  not U31767(n28174,G59331);
  nor U31768(n30021,n29261,n30015);
  nand U31769(n30019,n29197,n28175);
  nand U31770(n30018,n28491,n29784,n30023);
  nand U31771(n30017,n28173,n29788);
  nand U31772(n29788,n29541,n30024);
  nand U31773(n30024,n29264,n29784);
  nand U31774(n29784,n28173,n30025,n28491,n28495);
  xnor U31775(n30016,n29205,n30005);
  nand U31776(n30005,n30026,n30027);
  nand U31777(n30027,n29197,n30028);
  or U31778(n30028,n30029,n30030);
  nand U31779(n30026,n30030,n30029);
  nand U31780(n30007,n29231,n28173);
  xor U31781(n28173,n30001,n30031);
  and U31782(n30031,n29998,n30000);
  nand U31783(n30000,n30032,n30033,n30034);
  nand U31784(n30034,n29349,n30035);
  nand U31785(n29998,n30036,n30035,n29349);
  nand U31786(n30036,n30032,n30033);
  nand U31787(n30033,n29226,n28650,n30037);
  not U31788(n28650,n28175);
  nand U31789(n30032,n30038,n29174);
  nand U31790(n30038,n30037,n30039);
  nand U31791(n30039,n28175,n29288);
  nor U31792(n28175,n30040,n29710);
  nor U31793(n29710,n30041,n30042,n30043);
  and U31794(n30040,n30041,n30044);
  or U31795(n30044,n30043,n30042);
  xor U31796(n30041,n30045,n28963);
  nand U31797(n30045,n30046,n30047,n30048,n30049);
  nor U31798(n30049,n30050,n30051);
  and U31799(n30051,n29228,G59267);
  nor U31800(n30050,n29486,n30015);
  nand U31801(n30048,G59172,n29226);
  nand U31802(n30047,n28576,n30014);
  nand U31803(n30014,n30052,n30053,n30054);
  nand U31804(n30054,n29952,n30015);
  not U31805(n30015,G59140);
  not U31806(n29952,n30055);
  nand U31807(n30053,G59140,n30055,n27943);
  nand U31808(n30055,G59139,n30056);
  nand U31809(n30052,n29444,n28689);
  nand U31810(n29444,n30057,n30058,n30059,n30060);
  nor U31811(n30060,n30061,n30062,n30063,n30064);
  nor U31812(n30064,n29434,n29962);
  nor U31813(n30063,n29436,n29964);
  nor U31814(n30062,n29438,n29966);
  nor U31815(n30061,n29440,n29968);
  nor U31816(n30059,n30065,n30066,n30067,n30068);
  nor U31817(n30068,n29422,n29974);
  nor U31818(n30067,n29424,n29976);
  nor U31819(n30066,n29426,n29978);
  nor U31820(n30065,n29428,n29980);
  nor U31821(n30058,n30069,n30070,n30071,n30072);
  nor U31822(n30072,n29414,n29985);
  nor U31823(n30071,n29415,n29986);
  nor U31824(n30070,n29416,n29987);
  nor U31825(n30069,n29417,n29988);
  nor U31826(n30057,n30073,n30074,n30075,n30076);
  nor U31827(n30076,n29406,n29993);
  nor U31828(n30075,n29407,n29994);
  nor U31829(n30074,n29408,n29995);
  nor U31830(n30073,n29409,n29996);
  nand U31831(n30046,G59299,n29225);
  and U31832(n30037,n30077,n30078,n30079);
  nand U31833(n30079,G59172,n30080);
  nand U31834(n30078,G59140,n29287);
  nand U31835(n30077,G59331,n27993);
  nand U31836(n30001,n30081,n30082);
  nand U31837(n30082,n30083,n30084);
  nand U31838(G2534,n30085,n30086,n30087,n30088);
  nor U31839(n30088,n30089,n30090,n30091);
  nor U31840(n30091,n28186,n29192);
  not U31841(n28186,G59330);
  and U31842(n30090,n30092,n29688);
  nor U31843(n30089,n30093,n29247);
  nand U31844(n30087,n29193,n28187);
  nand U31845(n30086,n29194,n28188);
  xor U31846(n28188,n30094,n30030);
  nand U31847(n30030,n30095,n30096,n30097,n30098);
  nor U31848(n30098,n30099,n30100);
  nor U31849(n30100,n29261,n30093);
  nor U31850(n30099,n28657,n29205);
  nand U31851(n30097,n29230,G59330);
  nand U31852(n30096,n28185,n30023);
  nor U31853(n30023,n28197,n28761,n30101);
  nand U31854(n30095,n28491,n30102);
  nand U31855(n30102,n30103,n30104);
  nand U31856(n30104,n29264,n28197);
  not U31857(n30103,n30105);
  xnor U31858(n30094,n29205,n30029);
  nand U31859(n30029,n30106,n30107);
  nand U31860(n30107,n29197,n30108);
  or U31861(n30108,n30109,n30110);
  nand U31862(n30106,n30110,n30109);
  nand U31863(n30085,n29231,n28491);
  not U31864(n28491,n28185);
  xnor U31865(n28185,n30084,n30111);
  and U31866(n30111,n30081,n30083);
  nand U31867(n30083,n30112,n30113,n30114);
  nand U31868(n30114,n29349,n30115);
  nand U31869(n30081,n30116,n30115,n29349);
  nand U31870(n30116,n30112,n30113);
  nand U31871(n30113,n29226,n28657,n30117);
  nand U31872(n30112,n30118,n29174);
  nand U31873(n30118,n30117,n30119);
  nand U31874(n30119,n28187,n29288);
  not U31875(n28187,n28657);
  xnor U31876(n28657,n30043,n30042);
  xor U31877(n30042,n27993,n30120);
  nor U31878(n30120,n30121,n30122,n30123);
  and U31879(n30123,n29228,G59266);
  nor U31880(n30122,n29486,n30093);
  nand U31881(n30121,n30124,n30125,n30126);
  nand U31882(n30126,G59171,n29226);
  nand U31883(n30125,n28576,n30092);
  nand U31884(n30092,n30127,n30128);
  nand U31885(n30128,n29522,n28689);
  nand U31886(n29522,n30129,n30130,n30131,n30132);
  nor U31887(n30132,n30133,n30134,n30135,n30136);
  nor U31888(n30136,n30137,n29962);
  nor U31889(n30135,n30138,n29964);
  nor U31890(n30134,n30139,n29966);
  nor U31891(n30133,n30140,n29968);
  nor U31892(n30131,n30141,n30142,n30143,n30144);
  nor U31893(n30144,n30145,n29974);
  nor U31894(n30143,n30146,n29976);
  nor U31895(n30142,n30147,n29978);
  nor U31896(n30141,n30148,n29980);
  nor U31897(n30130,n30149,n30150,n30151,n30152);
  nor U31898(n30152,n29518,n29985);
  nor U31899(n30151,n29519,n29986);
  nor U31900(n30150,n29520,n29987);
  nor U31901(n30149,n29521,n29988);
  nor U31902(n30129,n30153,n30154,n30155,n30156);
  nor U31903(n30156,n29510,n29993);
  nor U31904(n30155,n29511,n29994);
  nor U31905(n30154,n29512,n29995);
  nor U31906(n30153,n29513,n29996);
  nand U31907(n30127,n30157,n27943);
  xnor U31908(n30157,n30093,n30056);
  nor U31909(n30056,n30158,n30159);
  not U31910(n30093,G59139);
  nand U31911(n30124,G59298,n29225);
  and U31912(n30117,n30160,n30161,n30162);
  nand U31913(n30162,G59171,n30080);
  nand U31914(n30161,G59139,n29287);
  nand U31915(n30160,G59330,n27993);
  nand U31916(n30084,n30163,n30164);
  nand U31917(n30164,n30165,n30166);
  nand U31918(G2533,n30167,n30168,n30169,n30170);
  nor U31919(n30170,n30171,n30172,n30173);
  nor U31920(n30173,n28198,n29192);
  not U31921(n28198,G59329);
  and U31922(n30172,n30174,n29688);
  nor U31923(n30171,n30159,n29247);
  nand U31924(n30169,n29193,n28199);
  nand U31925(n30168,n29194,n28200);
  xor U31926(n28200,n30175,n30110);
  nand U31927(n30110,n30176,n30177,n30178,n30179);
  nor U31928(n30179,n30180,n30181);
  nor U31929(n30181,n29261,n30159);
  nor U31930(n30180,n28664,n29205);
  nand U31931(n30178,n29230,G59329);
  nand U31932(n30177,n28495,n30105);
  nand U31933(n30176,n30025,n29264,n28197);
  not U31934(n30025,n30101);
  xnor U31935(n30175,n29205,n30109);
  nand U31936(n30109,n30182,n30183);
  nand U31937(n30183,n29197,n30184);
  or U31938(n30184,n30185,n30186);
  nand U31939(n30182,n30186,n30185);
  nand U31940(n30167,n29231,n28495);
  not U31941(n28495,n28197);
  xnor U31942(n28197,n30166,n30187);
  and U31943(n30187,n30163,n30165);
  nand U31944(n30165,n30188,n30189,n30190);
  nand U31945(n30163,n30192,n30191,n29349);
  nand U31946(n30192,n30188,n30189);
  nand U31947(n30189,n29226,n28664,n30193);
  nand U31948(n30188,n30194,n29174);
  nand U31949(n30194,n30193,n30195);
  nand U31950(n30195,n28199,n29288);
  not U31951(n28199,n28664);
  nand U31952(n28664,n30043,n30196);
  nand U31953(n30196,n30197,n30198);
  or U31954(n30043,n30198,n30197);
  xor U31955(n30197,n30199,n28963);
  nand U31956(n30199,n30200,n30201,n30202,n30203);
  nor U31957(n30203,n30204,n30205);
  and U31958(n30205,n29228,G59265);
  nor U31959(n30204,n29486,n30159);
  not U31960(n30159,G59138);
  nand U31961(n30202,G59170,n29226);
  nand U31962(n30201,n28576,n30174);
  nand U31963(n30174,n30206,n30207,n30208);
  or U31964(n30208,n30158,G59138);
  nand U31965(n30207,G59138,n30158,n27943);
  nand U31966(n30158,n30209,G59137);
  nand U31967(n30206,n29605,n28689);
  nand U31968(n29605,n30210,n30211,n30212,n30213);
  nor U31969(n30213,n30214,n30215,n30216,n30217);
  nor U31970(n30217,n30218,n29962);
  nor U31971(n30216,n30219,n29964);
  nor U31972(n30215,n30220,n29966);
  nor U31973(n30214,n30221,n29968);
  nor U31974(n30212,n30222,n30223,n30224,n30225);
  nor U31975(n30225,n30226,n29974);
  nor U31976(n30224,n30227,n29976);
  nor U31977(n30223,n30228,n29978);
  nor U31978(n30222,n30229,n29980);
  nor U31979(n30211,n30230,n30231,n30232,n30233);
  nor U31980(n30233,n29597,n29985);
  nor U31981(n30232,n29598,n29986);
  nor U31982(n30231,n29599,n29987);
  nor U31983(n30230,n29600,n29988);
  nor U31984(n30210,n30234,n30235,n30236,n30237);
  nor U31985(n30237,n29589,n29993);
  nor U31986(n30236,n29590,n29994);
  nor U31987(n30235,n29591,n29995);
  nor U31988(n30234,n29592,n29996);
  nand U31989(n30200,G59297,n29225);
  and U31990(n30193,n30238,n30239,n30240);
  nand U31991(n30240,G59170,n30080);
  nand U31992(n30239,G59138,n29287);
  nand U31993(n30238,G59329,n27993);
  nand U31994(n30166,n30241,n30242);
  nand U31995(n30242,n30243,n30244);
  nand U31996(G2532,n30245,n30246,n30247,n30248);
  nor U31997(n30248,n30249,n30250,n30251);
  nor U31998(n30251,n30252,n29192);
  and U31999(n30250,n30253,n29688);
  nor U32000(n30249,n30254,n29247);
  nand U32001(n30247,n29193,n28499);
  nand U32002(n30246,n29194,n28211);
  xor U32003(n28211,n30255,n30186);
  nand U32004(n30186,n30256,n30257,n30258,n30259);
  nor U32005(n30259,n30260,n30261);
  nor U32006(n30261,n30252,n29260);
  not U32007(n30252,G59328);
  nor U32008(n30260,n29261,n30254);
  nand U32009(n30258,n29197,n28499);
  nand U32010(n30257,n28234,n30262,n28224,n30101);
  nand U32011(n30256,n28213,n30105);
  nand U32012(n30105,n29541,n30263);
  nand U32013(n30263,n29264,n30101);
  nand U32014(n30101,n28244,n30264,n28224,n30265);
  and U32015(n30265,n28213,n28234);
  xnor U32016(n30255,n29205,n30185);
  nand U32017(n30185,n30266,n30267);
  nand U32018(n30267,n29197,n30268);
  or U32019(n30268,n30269,n30270);
  nand U32020(n30266,n30270,n30269);
  nand U32021(n30245,n29231,n28213);
  xor U32022(n28213,n30244,n30271);
  and U32023(n30271,n30241,n30243);
  nand U32024(n30243,n30272,n30273,n30274);
  nand U32025(n30241,n30276,n30275,n29349);
  nand U32026(n30276,n30272,n30273);
  nand U32027(n30273,n29226,n28210,n30277);
  nand U32028(n30272,n30278,n29174);
  nand U32029(n30278,n30277,n30279);
  nand U32030(n30279,n28499,n29288);
  not U32031(n28499,n28210);
  nand U32032(n28210,n30280,n30198);
  or U32033(n30198,n30281,n30282,n30283);
  nand U32034(n30280,n30281,n30284);
  or U32035(n30284,n30283,n30282);
  xor U32036(n30281,n27993,n30285);
  nor U32037(n30285,n30286,n30287,n30288);
  and U32038(n30288,n29228,G59264);
  nor U32039(n30287,n29486,n30254);
  nand U32040(n30286,n30289,n30290,n30291);
  nand U32041(n30291,G59169,n29226);
  nand U32042(n30290,n28576,n30253);
  nand U32043(n30253,n30292,n30293);
  nand U32044(n30293,n29677,n28689);
  nand U32045(n29677,n30294,n30295,n30296,n30297);
  nor U32046(n30297,n30298,n30299,n30300,n30301);
  nor U32047(n30301,n30302,n29962);
  nor U32048(n30300,n30303,n29964);
  nor U32049(n30299,n30304,n29966);
  nor U32050(n30298,n30305,n29968);
  nor U32051(n30296,n30306,n30307,n30308,n30309);
  nor U32052(n30309,n30310,n29974);
  nor U32053(n30308,n30311,n29976);
  nor U32054(n30307,n30312,n29978);
  nor U32055(n30306,n30313,n29980);
  nor U32056(n30295,n30314,n30315,n30316,n30317);
  nor U32057(n30317,n29673,n29985);
  nor U32058(n30316,n29674,n29986);
  nor U32059(n30315,n29675,n29987);
  nor U32060(n30314,n29676,n29988);
  nor U32061(n30294,n30318,n30319,n30320,n30321);
  nor U32062(n30321,n29665,n29993);
  nor U32063(n30320,n29666,n29994);
  nor U32064(n30319,n29667,n29995);
  nor U32065(n30318,n29668,n29996);
  nand U32066(n30292,n30322,n27943);
  xnor U32067(n30322,n30254,n30209);
  nor U32068(n30209,n30323,n30324);
  not U32069(n30254,G59137);
  nand U32070(n30289,G59296,n29225);
  and U32071(n30277,n30325,n30326,n30327);
  nand U32072(n30327,G59169,n30080);
  nand U32073(n30326,G59137,n29287);
  nand U32074(n30325,G59328,n27993);
  nand U32075(n30244,n30328,n30329);
  nand U32076(n30329,n30330,n30331);
  nand U32077(G2531,n30332,n30333,n30334,n30335);
  nor U32078(n30335,n30336,n30337,n30338);
  nor U32079(n30338,n30339,n29192);
  not U32080(n30339,G59327);
  and U32081(n30337,n30340,n29688);
  nor U32082(n30336,n30323,n29247);
  nand U32083(n30334,n29193,n28503);
  nand U32084(n30333,n29194,n28223);
  xor U32085(n28223,n30341,n30270);
  nand U32086(n30270,n30342,n30343,n30344,n30345);
  nor U32087(n30345,n30346,n30347);
  nor U32088(n30347,n29261,n30323);
  nor U32089(n30346,n28222,n29205);
  nand U32090(n30344,n29230,G59327);
  nand U32091(n30343,n28224,n30348);
  nand U32092(n30348,n30349,n30350);
  nand U32093(n30350,n29264,n30351);
  nand U32094(n30342,n30262,n28234,n30352);
  xnor U32095(n30341,n29205,n30269);
  nand U32096(n30269,n30353,n30354);
  nand U32097(n30354,n29197,n30355);
  or U32098(n30355,n30356,n30357);
  nand U32099(n30353,n30357,n30356);
  nand U32100(n30332,n29231,n28224);
  not U32101(n28224,n30352);
  xnor U32102(n30352,n30330,n30358);
  and U32103(n30358,n30331,n30328);
  nand U32104(n30328,n30359,n30360,n29349);
  nand U32105(n30359,n30361,n30362);
  nand U32106(n30331,n30361,n30362,n30363);
  nand U32107(n30362,n29226,n28222,n30364);
  nand U32108(n30361,n30365,n29174);
  nand U32109(n30365,n30364,n30366);
  nand U32110(n30366,n28503,n29288);
  not U32111(n28503,n28222);
  xnor U32112(n28222,n30283,n30282);
  xor U32113(n30282,n30367,n28963);
  nand U32114(n30367,n30368,n30369,n30370,n30371);
  nor U32115(n30371,n30372,n30373);
  and U32116(n30373,n29228,G59263);
  nor U32117(n30372,n29486,n30323);
  not U32118(n30323,G59136);
  nand U32119(n30370,G59168,n29226);
  nand U32120(n30369,n28576,n30340);
  nand U32121(n30340,n30374,n30375,n30376);
  or U32122(n30376,n30324,G59136);
  nand U32123(n30375,G59136,n30324,n27943);
  nand U32124(n30324,n30377,n30378);
  nand U32125(n30374,n29762,n28689);
  nand U32126(n29762,n30379,n30380,n30381,n30382);
  nor U32127(n30382,n30383,n30384,n30385,n30386);
  nor U32128(n30386,n29758,n29962);
  nor U32129(n30385,n29759,n29964);
  nor U32130(n30384,n29760,n29966);
  nor U32131(n30383,n29761,n29968);
  nor U32132(n30381,n30387,n30388,n30389,n30390);
  nor U32133(n30390,n29750,n29974);
  nor U32134(n30389,n29751,n29976);
  nor U32135(n30388,n29752,n29978);
  nor U32136(n30387,n29753,n29980);
  nor U32137(n30380,n30391,n30392,n30393,n30394);
  nor U32138(n30394,n29742,n29985);
  nor U32139(n30393,n29743,n29986);
  nor U32140(n30392,n29744,n29987);
  nor U32141(n30391,n29745,n29988);
  nor U32142(n30379,n30395,n30396,n30397,n30398);
  nor U32143(n30398,n29734,n29993);
  nor U32144(n30397,n29735,n29994);
  nor U32145(n30396,n29736,n29995);
  nor U32146(n30395,n29737,n29996);
  nand U32147(n30368,G59295,n29225);
  and U32148(n30364,n30399,n30400,n30401);
  nand U32149(n30401,G59168,n30080);
  nand U32150(n30400,G59136,n29287);
  nand U32151(n30399,G59327,n27993);
  nand U32152(n30330,n30402,n30403);
  nand U32153(n30403,n30404,n30405);
  nand U32154(G2530,n30406,n30407,n30408,n30409);
  nor U32155(n30409,n30410,n30411,n30412);
  nor U32156(n30412,n30413,n29192);
  not U32157(n30413,G59326);
  and U32158(n30411,n30414,n29688);
  nor U32159(n30410,n30415,n29247);
  nand U32160(n30408,n29193,n28507);
  nand U32161(n30407,n29194,n28233);
  xor U32162(n28233,n30416,n30357);
  nand U32163(n30357,n30417,n30418,n30419,n30420);
  nor U32164(n30420,n30421,n30422);
  nor U32165(n30422,n29261,n30415);
  nor U32166(n30421,n28232,n29205);
  nand U32167(n30419,n29230,G59326);
  nand U32168(n30418,n30262,n30351);
  nor U32169(n30262,n30423,n30424,n28761);
  or U32170(n30417,n30351,n30349);
  nor U32171(n30349,n30425,n30426);
  nor U32172(n30426,n28244,n28761);
  xnor U32173(n30416,n29205,n30356);
  nand U32174(n30356,n30427,n30428);
  nand U32175(n30428,n29197,n30429);
  or U32176(n30429,n30430,n30431);
  nand U32177(n30427,n30431,n30430);
  nand U32178(n30406,n29231,n28234);
  not U32179(n28234,n30351);
  xnor U32180(n30351,n30404,n30432);
  and U32181(n30432,n30405,n30402);
  nand U32182(n30402,n30433,n30434,n29349);
  nand U32183(n30433,n30435,n30436);
  nand U32184(n30405,n30435,n30436,n30437);
  nand U32185(n30436,n29226,n28232,n30438);
  nand U32186(n30435,n30439,n29174);
  nand U32187(n30439,n30438,n30440);
  nand U32188(n30440,n28507,n29288);
  not U32189(n28507,n28232);
  nand U32190(n28232,n30283,n30441);
  nand U32191(n30441,n30442,n30443);
  or U32192(n30283,n30443,n30442);
  xor U32193(n30442,n27993,n30444);
  nor U32194(n30444,n30445,n30446,n30447);
  and U32195(n30447,n29228,G59262);
  nor U32196(n30446,n29486,n30415);
  nand U32197(n30445,n30448,n30449,n30450);
  nand U32198(n30450,G59167,n29226);
  nand U32199(n30449,n28576,n30414);
  nand U32200(n30414,n30451,n30452);
  nand U32201(n30452,n29860,n28689);
  nand U32202(n29860,n30453,n30454,n30455,n30456);
  nor U32203(n30456,n30457,n30458,n30459,n30460);
  nor U32204(n30460,n29854,n29962);
  nor U32205(n30459,n29855,n29964);
  nor U32206(n30458,n29856,n29966);
  nor U32207(n30457,n29857,n29968);
  nor U32208(n30455,n30461,n30462,n30463,n30464);
  nor U32209(n30464,n29846,n29974);
  nor U32210(n30463,n29847,n29976);
  nor U32211(n30462,n29848,n29978);
  nor U32212(n30461,n29849,n29980);
  nor U32213(n30454,n30465,n30466,n30467,n30468);
  nor U32214(n30468,n29838,n29985);
  nor U32215(n30467,n29839,n29986);
  nor U32216(n30466,n29840,n29987);
  nor U32217(n30465,n29841,n29988);
  nor U32218(n30453,n30469,n30470,n30471,n30472);
  nor U32219(n30472,n29830,n29993);
  nor U32220(n30471,n29831,n29994);
  nor U32221(n30470,n29832,n29995);
  nor U32222(n30469,n29833,n29996);
  xnor U32223(n30451,n30378,n30377);
  nor U32224(n30377,n30473,n30474);
  nor U32225(n30378,n30415,n28689);
  not U32226(n30415,G59135);
  nand U32227(n30448,G59294,n29225);
  and U32228(n30438,n30475,n30476,n30477);
  nand U32229(n30477,G59167,n30080);
  nand U32230(n30476,G59135,n29287);
  nand U32231(n30475,G59326,n27993);
  nand U32232(n30404,n30478,n30479);
  nand U32233(n30479,n30480,n30481);
  not U32234(n30480,n30482);
  nand U32235(G2529,n30483,n30484,n30485,n30486);
  nor U32236(n30486,n30487,n30488,n30489);
  nor U32237(n30489,n30490,n29192);
  not U32238(n30490,G59325);
  and U32239(n30488,n30491,n29688);
  nor U32240(n30487,n30474,n29247);
  nand U32241(n30485,n29193,n28511);
  nand U32242(n30484,n29194,n28243);
  xor U32243(n28243,n30492,n30431);
  nand U32244(n30431,n30493,n30494);
  nand U32245(n30494,n29197,n30495);
  or U32246(n30495,n30496,n30497);
  nand U32247(n30493,n30497,n30496);
  xnor U32248(n30492,n30430,n29205);
  nand U32249(n30430,n30498,n30499,n30500,n30501);
  nor U32250(n30501,n30502,n30503);
  nor U32251(n30503,n29261,n30474);
  nor U32252(n30502,n28242,n29205);
  nand U32253(n30500,n29230,G59325);
  nand U32254(n30499,n28244,n30425);
  nand U32255(n30425,n29541,n30504);
  nand U32256(n30504,n30424,n29264);
  not U32257(n30424,n30264);
  nand U32258(n30498,n29264,n30264,n30423);
  not U32259(n30423,n28244);
  nand U32260(n30264,n30505,n30506);
  nand U32261(n30506,n30507,n30508);
  or U32262(n30507,n30509,n28254);
  nand U32263(n30505,n28254,n30509);
  nand U32264(n30483,n29231,n28244);
  xor U32265(n28244,n30510,n30482);
  nand U32266(n30510,n30478,n30481);
  nand U32267(n30481,n30511,n30512,n30513);
  nand U32268(n30478,n30515,n30514,n29349);
  nand U32269(n30515,n30511,n30512);
  nand U32270(n30512,n29226,n28242,n30516);
  nand U32271(n30511,n30517,n29174);
  nand U32272(n30517,n30516,n30518);
  nand U32273(n30518,n28511,n29288);
  not U32274(n28511,n28242);
  nand U32275(n28242,n30443,n30519);
  nand U32276(n30519,n30520,n30521);
  or U32277(n30443,n30521,n30520);
  and U32278(n30520,n30522,n30523);
  nand U32279(n30523,n30524,n30525);
  xor U32280(n30521,n30526,n28963);
  nand U32281(n30526,n30527,n30528,n30529,n30530);
  nor U32282(n30530,n30531,n30532);
  and U32283(n30532,n29228,G59261);
  nor U32284(n30531,n29486,n30474);
  nand U32285(n30529,G59166,n29226);
  nand U32286(n30528,n28576,n30491);
  nand U32287(n30491,n30533,n30534,n30535);
  nand U32288(n30535,n30536,n30474);
  not U32289(n30474,G59134);
  nand U32290(n30534,G59134,n30473,n27943);
  not U32291(n30473,n30536);
  nor U32292(n30536,n30537,n30538,n30539);
  nand U32293(n30533,n29997,n28689);
  nand U32294(n29997,n30540,n30541,n30542,n30543);
  nor U32295(n30543,n30544,n30545,n30546,n30547);
  nor U32296(n30547,n29942,n29962);
  nor U32297(n30546,n29946,n29964);
  nor U32298(n30545,n29947,n29966);
  nor U32299(n30544,n29949,n29968);
  nor U32300(n30542,n30548,n30549,n30550,n30551);
  nor U32301(n30551,n29933,n29974);
  nor U32302(n30550,n29935,n29976);
  nor U32303(n30549,n29936,n29978);
  nor U32304(n30548,n29937,n29980);
  nor U32305(n30541,n30552,n30553,n30554,n30555);
  nor U32306(n30555,n29923,n29985);
  nor U32307(n30554,n29925,n29986);
  nor U32308(n30553,n29926,n29987);
  nor U32309(n30552,n29927,n29988);
  nor U32310(n30540,n30556,n30557,n30558,n30559);
  nor U32311(n30559,n29908,n29993);
  nor U32312(n30558,n29911,n29994);
  nor U32313(n30557,n29913,n29995);
  nor U32314(n30556,n29915,n29996);
  nand U32315(n30527,G59293,n29225);
  and U32316(n30516,n30560,n30561,n30562);
  nand U32317(n30562,G59166,n30080);
  nand U32318(n30561,G59134,n29287);
  nand U32319(n30560,G59325,n27993);
  nand U32320(G2528,n30563,n30564,n30565,n30566);
  nor U32321(n30566,n30567,n30568,n30569);
  nor U32322(n30569,G59133,n29185,n30570,n30539);
  nor U32323(n30568,n30571,n30538);
  nor U32324(n30571,n30572,n29190);
  nor U32325(n30572,n30573,n29185);
  nor U32326(n30573,n30570,n30539);
  nor U32327(n30567,n30574,n29192);
  nand U32328(n30565,n29193,n28515);
  nand U32329(n30564,n29194,n28253);
  xor U32330(n28253,n30575,n30497);
  nand U32331(n30497,n30576,n30577,n30578,n30579);
  nor U32332(n30579,n30580,n30581);
  nor U32333(n30581,n30574,n29260);
  not U32334(n30574,G59324);
  nor U32335(n30580,n29261,n30538);
  not U32336(n30538,G59133);
  nand U32337(n30578,n29197,n28515);
  nand U32338(n30577,n29264,n30582);
  xor U32339(n30582,n30509,n30583);
  xor U32340(n30583,n28254,n30508);
  nand U32341(n30509,n30584,n30585);
  nand U32342(n30585,n30586,n30587);
  nand U32343(n30586,n30588,n30589);
  or U32344(n30584,n30588,n30589);
  nand U32345(n30576,n28254,n29214);
  xnor U32346(n30575,n29205,n30496);
  nand U32347(n30496,n30590,n30591);
  nand U32348(n30591,n29197,n30592);
  or U32349(n30592,n30593,n30594);
  nand U32350(n30590,n30594,n30593);
  nand U32351(n30563,n29231,n28254);
  and U32352(n28254,n30482,n30595);
  nand U32353(n30595,n30596,n30597);
  xnor U32354(n30596,n29226,n30598);
  nand U32355(n30482,n30599,n30600);
  xnor U32356(n30599,n30598,n29174);
  nand U32357(n30598,n30601,n30602,n30603,n30604);
  nand U32358(n30604,n28515,n29288);
  not U32359(n28515,n28252);
  xor U32360(n28252,n30605,n30524);
  nand U32361(n30524,n30606,n30607);
  nand U32362(n30607,n30608,n30609);
  nand U32363(n30605,n30525,n30522);
  nand U32364(n30522,n30610,n30508,n28576);
  nand U32365(n30525,n30611,n30612,n30613);
  nand U32366(n30613,n28576,n30508);
  nand U32367(n30508,n30614,n30615,n30616,n30617);
  nor U32368(n30617,n30618,n30619,n30620,n30621);
  nor U32369(n30621,n29965,n30622);
  nor U32370(n30620,n29963,n30623);
  nor U32371(n30619,n29961,n30624);
  nor U32372(n30618,n29977,n30625);
  nor U32373(n30616,n30626,n30627,n30628,n30629);
  nor U32374(n30629,n29975,n30630);
  nor U32375(n30628,n29973,n30631);
  nor U32376(n30627,n29345,n30632);
  nor U32377(n30626,n29343,n30633);
  nor U32378(n30615,n30634,n30635,n30636,n30637);
  nor U32379(n30637,n29341,n30638);
  nor U32380(n30636,n29333,n30639);
  nor U32381(n30635,n29331,n30640);
  nor U32382(n30634,n29329,n30641);
  nor U32383(n30614,n30642,n30643,n30644,n30645);
  nor U32384(n30645,n29967,n30646);
  nor U32385(n30644,n29979,n30647);
  nor U32386(n30643,n29347,n30648);
  nor U32387(n30642,n29335,n30649);
  nand U32388(n30612,n30650,n27993);
  nand U32389(n30611,n30610,n28963);
  nand U32390(n30610,n30651,n30652,n30650);
  and U32391(n30650,n30653,n30654);
  nand U32392(n30654,G59292,n29225);
  nand U32393(n30653,G59165,n29226);
  nand U32394(n30652,G59133,n29227);
  nand U32395(n30651,G59260,n29228);
  nand U32396(n30603,G59133,n29287);
  nand U32397(n30602,G59324,n27993);
  nand U32398(n30601,G59165,n30080);
  nand U32399(G2527,n30655,n30656,n30657,n30658);
  nor U32400(n30658,n30659,n30660,n30661);
  nor U32401(n30661,n28262,n29685);
  nor U32402(n30660,n30588,n30662);
  nor U32403(n30659,n30663,n29192);
  nand U32404(n30657,n29194,n28263);
  xor U32405(n28263,n30664,n30594);
  nand U32406(n30594,n30665,n30666,n30667,n30668);
  nor U32407(n30668,n30669,n30670);
  nor U32408(n30670,n30663,n29260);
  not U32409(n30663,G59323);
  nor U32410(n30669,n29261,n30570);
  not U32411(n30570,G59132);
  nand U32412(n30667,n29197,n28519);
  nand U32413(n30666,n30671,n29264);
  xor U32414(n30671,n30589,n30672);
  xnor U32415(n30672,n30587,n28264);
  nand U32416(n30589,n30673,n30674);
  nand U32417(n30674,n30675,n30676);
  or U32418(n30676,n30677,n30678);
  nand U32419(n30673,n30678,n30677);
  nand U32420(n30665,n28264,n29214);
  not U32421(n28264,n30588);
  nand U32422(n30588,n30597,n30679);
  nand U32423(n30679,n30680,n30681);
  not U32424(n30597,n30600);
  nor U32425(n30600,n30681,n30680);
  xor U32426(n30680,n30682,n29174);
  nand U32427(n30682,n30683,n30684,n30685,n30686);
  nand U32428(n30686,n28519,n29288);
  not U32429(n28519,n28262);
  xor U32430(n28262,n30687,n30609);
  nand U32431(n30609,n30688,n30689);
  nand U32432(n30689,n30690,n30691);
  nand U32433(n30687,n30606,n30608);
  nand U32434(n30608,n30692,n30693);
  nand U32435(n30693,n28576,n30587);
  xnor U32436(n30692,n27993,n30694);
  nand U32437(n30606,n30694,n30587,n28576);
  nand U32438(n30587,n30695,n30696,n30697,n30698);
  nor U32439(n30698,n30699,n30700,n30701,n30702);
  nor U32440(n30702,n29438,n30622);
  nor U32441(n30701,n29436,n30623);
  nor U32442(n30700,n29434,n30624);
  nor U32443(n30699,n29426,n30625);
  nor U32444(n30697,n30703,n30704,n30705,n30706);
  nor U32445(n30706,n29424,n30630);
  nor U32446(n30705,n29422,n30631);
  nor U32447(n30704,n29416,n30632);
  nor U32448(n30703,n29415,n30633);
  nor U32449(n30696,n30707,n30708,n30709,n30710);
  nor U32450(n30710,n29414,n30638);
  nor U32451(n30709,n29408,n30639);
  nor U32452(n30708,n29407,n30640);
  nor U32453(n30707,n29406,n30641);
  nor U32454(n30695,n30711,n30712,n30713,n30714);
  nor U32455(n30714,n29440,n30646);
  nor U32456(n30713,n29428,n30647);
  nor U32457(n30712,n29417,n30648);
  nor U32458(n30711,n29409,n30649);
  nand U32459(n30694,n30715,n30716,n30717,n30718);
  nand U32460(n30718,G59291,n29225);
  nand U32461(n30717,G59164,n29226);
  nand U32462(n30716,G59132,n29227);
  nand U32463(n30715,G59259,n29228);
  nand U32464(n30685,G59132,n29287);
  nand U32465(n30684,G59323,n27993);
  nand U32466(n30683,G59164,n30080);
  xnor U32467(n30664,n29205,n30593);
  nand U32468(n30593,n30719,n30720);
  nand U32469(n30720,n29197,n30721);
  nand U32470(n30721,n30722,n30723);
  or U32471(n30719,n30723,n30722);
  nand U32472(n30656,n30724,n30537,n29688);
  nand U32473(n30537,G59132,n27943);
  nand U32474(n30655,G59132,n30725);
  nand U32475(n30725,n29247,n30726);
  nand U32476(n30726,n29688,n30539);
  not U32477(n30539,n30724);
  nor U32478(n30724,n30727,n30728,n30729);
  nand U32479(G2526,n30730,n30731,n30732,n30733);
  nor U32480(n30733,n30734,n30735,n30736);
  nor U32481(n30736,G59131,n29185,n30737,n30729);
  nor U32482(n30735,n30738,n30728);
  nor U32483(n30738,n30739,n30740);
  nor U32484(n30739,G59130,n29185);
  nor U32485(n30734,n30741,n29192);
  nand U32486(n30732,n29193,n28523);
  nand U32487(n30731,n29194,n28273);
  xnor U32488(n28273,n30722,n30742);
  xnor U32489(n30742,n29197,n30723);
  nand U32490(n30723,n30743,n30744);
  nand U32491(n30744,n30745,n29205);
  nand U32492(n30745,n30746,n30747);
  or U32493(n30743,n30746,n30747);
  and U32494(n30722,n30748,n30749,n30750,n30751);
  nor U32495(n30751,n30752,n30753);
  nor U32496(n30753,n30741,n29260);
  not U32497(n30741,G59322);
  nor U32498(n30752,n29261,n30728);
  not U32499(n30728,G59131);
  nand U32500(n30750,n29197,n28523);
  nand U32501(n30749,n30754,n29264);
  xor U32502(n30754,n30678,n30755);
  xnor U32503(n30755,n30675,n30677);
  not U32504(n30675,n30756);
  nand U32505(n30678,n30757,n30758);
  nand U32506(n30758,n30759,n30760);
  or U32507(n30760,n30761,n30762);
  not U32508(n30759,n30763);
  nand U32509(n30757,n30762,n30761);
  nand U32510(n30748,n28274,n29214);
  nand U32511(n30730,n29231,n28274);
  not U32512(n28274,n30677);
  nand U32513(n30677,n30681,n30764);
  nand U32514(n30764,n30765,n30766);
  or U32515(n30681,n30766,n30765);
  xor U32516(n30765,n30767,n29174);
  nand U32517(n30767,n30768,n30769,n30770,n30771);
  nand U32518(n30771,n28523,n29288);
  not U32519(n28523,n28272);
  xor U32520(n28272,n30772,n30690);
  or U32521(n30690,n30773,n30774);
  nor U32522(n30774,n30775,n30776);
  nand U32523(n30772,n30691,n30688);
  nand U32524(n30688,n30777,n30756,n28576);
  nand U32525(n30691,n30778,n30779,n30780);
  nand U32526(n30780,n28576,n30756);
  nand U32527(n30756,n30781,n30782,n30783,n30784);
  nor U32528(n30784,n30785,n30786,n30787,n30788);
  nor U32529(n30788,n30139,n30622);
  nor U32530(n30787,n30138,n30623);
  nor U32531(n30786,n30137,n30624);
  nor U32532(n30785,n30147,n30625);
  nor U32533(n30783,n30789,n30790,n30791,n30792);
  nor U32534(n30792,n30146,n30630);
  nor U32535(n30791,n30145,n30631);
  nor U32536(n30790,n29520,n30632);
  nor U32537(n30789,n29519,n30633);
  nor U32538(n30782,n30793,n30794,n30795,n30796);
  nor U32539(n30796,n29518,n30638);
  nor U32540(n30795,n29512,n30639);
  nor U32541(n30794,n29511,n30640);
  nor U32542(n30793,n29510,n30641);
  nor U32543(n30781,n30797,n30798,n30799,n30800);
  nor U32544(n30800,n30140,n30646);
  nor U32545(n30799,n30148,n30647);
  nor U32546(n30798,n29521,n30648);
  nor U32547(n30797,n29513,n30649);
  nand U32548(n30779,n30801,n27993);
  nand U32549(n30778,n30777,n28963);
  nand U32550(n30777,n30802,n30803,n30801);
  and U32551(n30801,n30804,n30805);
  nand U32552(n30805,G59290,n29225);
  nand U32553(n30804,G59163,n29226);
  nand U32554(n30803,G59131,n29227);
  nand U32555(n30802,G59258,n29228);
  nand U32556(n30770,G59131,n29287);
  nand U32557(n30769,G59322,n27993);
  nand U32558(n30768,G59163,n30080);
  nand U32559(n30766,n30806,n30807);
  nand U32560(G2525,n30808,n30809,n30810,n30811);
  nor U32561(n30811,n30812,n30813,n30814);
  nor U32562(n30814,n28282,n29685);
  not U32563(n28282,n28527);
  nor U32564(n30813,n30762,n30662);
  nor U32565(n30812,n30815,n29192);
  nand U32566(n30810,n29194,n28283);
  xnor U32567(n28283,n30747,n30816);
  xnor U32568(n30816,n29197,n30746);
  nand U32569(n30746,n30817,n30818,n30819,n30820);
  nor U32570(n30820,n30821,n30822);
  nor U32571(n30822,n30815,n29260);
  not U32572(n30815,G59321);
  nor U32573(n30821,n29261,n30737);
  not U32574(n30737,G59130);
  nand U32575(n30819,n29197,n28527);
  nand U32576(n30818,n29264,n30823);
  xnor U32577(n30823,n30762,n30824);
  xnor U32578(n30824,n30761,n30763);
  nand U32579(n30761,n30825,n30826);
  nand U32580(n30826,n30827,n30828);
  or U32581(n30828,n30829,n30830);
  not U32582(n30827,n30831);
  nand U32583(n30825,n30830,n30829);
  nand U32584(n30817,n28284,n29214);
  not U32585(n28284,n30762);
  xnor U32586(n30762,n30807,n30806);
  xnor U32587(n30807,n30832,n29174);
  nand U32588(n30832,n30833,n30834,n30835,n30836);
  nand U32589(n30836,n28527,n29288);
  xnor U32590(n28527,n30775,n30837);
  nor U32591(n30837,n30773,n30776);
  and U32592(n30776,n30838,n30839,n30840);
  nand U32593(n30840,n30841,n27993);
  nor U32594(n30773,n30839,n30838);
  nand U32595(n30838,n28576,n30763);
  nand U32596(n30763,n30842,n30843,n30844,n30845);
  nor U32597(n30845,n30846,n30847,n30848,n30849);
  nor U32598(n30849,n29590,n30640);
  nor U32599(n30848,n29591,n30639);
  nor U32600(n30847,n29599,n30632);
  nor U32601(n30846,n30228,n30625);
  nor U32602(n30844,n30850,n30851,n30852,n30853);
  nor U32603(n30853,n29598,n30633);
  nor U32604(n30852,n29600,n30648);
  nor U32605(n30851,n30221,n30646);
  nor U32606(n30850,n29589,n30641);
  nor U32607(n30843,n30854,n30855,n30856,n30857);
  nor U32608(n30857,n30227,n30630);
  nor U32609(n30856,n30229,n30647);
  nor U32610(n30855,n30218,n30624);
  nor U32611(n30854,n29597,n30638);
  nor U32612(n30842,n30858,n30859,n30860,n30861);
  nor U32613(n30861,n30219,n30623);
  nor U32614(n30860,n30226,n30631);
  nor U32615(n30859,n29592,n30649);
  nor U32616(n30858,n30220,n30622);
  nand U32617(n30839,n30862,n28963);
  nand U32618(n30862,n30863,n30864,n30841);
  and U32619(n30841,n30865,n30866);
  nand U32620(n30866,G59289,n29225);
  nand U32621(n30865,G59162,n29226);
  nand U32622(n30864,G59130,n29227);
  nand U32623(n30863,G59257,n29228);
  nand U32624(n30775,n30867,n30868);
  nand U32625(n30868,n30869,n30870,n30871);
  nand U32626(n30835,G59130,n29287);
  nand U32627(n30834,G59321,n27993);
  nand U32628(n30833,G59162,n30080);
  nand U32629(n30747,n30872,n30873,n30874);
  or U32630(n30874,n29205,n30875);
  nor U32631(n30875,n30876,n30877,n30878);
  nand U32632(n30872,n30878,n30879,n30877);
  nand U32633(n30809,n30880,n30727,n29688);
  nand U32634(n30727,G59130,n27943);
  nand U32635(n30808,G59130,n30740);
  nand U32636(n30740,n29247,n30881);
  nand U32637(n30881,n29688,n30729);
  not U32638(n30729,n30880);
  nor U32639(n30880,n30882,n30883,n30884,n30885);
  nand U32640(G2524,n30886,n30887,n30888,n30889);
  nor U32641(n30889,n30890,n30891,n30892);
  nor U32642(n30892,G59129,n30885,n30893);
  nor U32643(n30891,n30894,n30883);
  nor U32644(n30894,n30895,n30896);
  nor U32645(n30895,G59128,n29185);
  nor U32646(n30890,n30897,n29192);
  nand U32647(n30888,n29193,n28531);
  nand U32648(n30887,n29194,n28293);
  xnor U32649(n28293,n30898,n30899);
  nor U32650(n30899,n30876,n30900);
  not U32651(n30876,n30901);
  xnor U32652(n30898,n30878,n29205);
  nand U32653(n30878,n30902,n30903,n30904,n30905);
  nor U32654(n30905,n30906,n30907);
  nor U32655(n30907,n30897,n29260);
  not U32656(n30897,G59320);
  nor U32657(n30906,n29261,n30883);
  not U32658(n30883,G59129);
  nand U32659(n30904,n29197,n28531);
  nand U32660(n30903,n30908,n29264);
  xnor U32661(n30908,n30909,n30830);
  not U32662(n30830,n28294);
  xnor U32663(n30909,n30829,n30831);
  nand U32664(n30829,n30910,n30911);
  nand U32665(n30911,n30912,n30913);
  nand U32666(n30913,n28307,n30914);
  nand U32667(n30910,n30915,n29102);
  nand U32668(n30902,n28294,n29214);
  nand U32669(n30886,n29231,n28294);
  nor U32670(n28294,n30806,n30916);
  and U32671(n30916,n30917,n30918);
  nor U32672(n30806,n30918,n30917);
  xor U32673(n30917,n30919,n29174);
  nand U32674(n30919,n30920,n30921,n30922,n30923);
  nand U32675(n30923,n28531,n29288);
  not U32676(n28531,n28292);
  xnor U32677(n28292,n30924,n30925);
  and U32678(n30925,n30871,n30867);
  nand U32679(n30867,n30926,n30927,n30928);
  nand U32680(n30928,n28576,n30831);
  nand U32681(n30927,n30929,n28963);
  nand U32682(n30926,n30930,n27993);
  nand U32683(n30871,n30929,n30831,n28576);
  nand U32684(n30831,n30931,n30932,n30933,n30934);
  nor U32685(n30934,n30935,n30936,n30937,n30938);
  nor U32686(n30938,n29666,n30640);
  nor U32687(n30937,n29667,n30639);
  nor U32688(n30936,n29675,n30632);
  nor U32689(n30935,n30312,n30625);
  nor U32690(n30933,n30939,n30940,n30941,n30942);
  nor U32691(n30942,n29674,n30633);
  nor U32692(n30941,n29676,n30648);
  nor U32693(n30940,n30305,n30646);
  nor U32694(n30939,n29665,n30641);
  nor U32695(n30932,n30943,n30944,n30945,n30946);
  nor U32696(n30946,n30311,n30630);
  nor U32697(n30945,n30313,n30647);
  nor U32698(n30944,n30302,n30624);
  nor U32699(n30943,n29673,n30638);
  nor U32700(n30931,n30947,n30948,n30949,n30950);
  nor U32701(n30950,n30303,n30623);
  nor U32702(n30949,n30310,n30631);
  nor U32703(n30948,n29668,n30649);
  nor U32704(n30947,n30304,n30622);
  nand U32705(n30929,n30951,n30952,n30930);
  and U32706(n30930,n30953,n30954);
  nand U32707(n30954,G59288,n29225);
  nand U32708(n30953,G59161,n29226);
  nand U32709(n30952,G59129,n29227);
  nand U32710(n30951,G59256,n29228);
  nand U32711(n30924,n30870,n30869);
  nand U32712(n30922,G59129,n29287);
  nand U32713(n30921,G59320,n27993);
  nand U32714(n30920,G59161,n30080);
  nand U32715(G2523,n30955,n30956,n30957,n30958);
  nor U32716(n30958,n30959,n30960,n30961);
  and U32717(n30961,n30896,G59128);
  nand U32718(n30896,n30962,n30963);
  nand U32719(n30963,n29688,n30884);
  nor U32720(n30960,G59128,n30893);
  nand U32721(n30893,n30964,G59127,n29688);
  nor U32722(n30959,n29104,n29192);
  nand U32723(n30957,n29193,n28535);
  nand U32724(n30956,n29194,n28717);
  not U32725(n28717,n28306);
  nand U32726(n28306,n30965,n30966);
  nand U32727(n30966,n30967,n30873,n30968);
  nand U32728(n30968,n30969,n30901);
  nand U32729(n30965,n30901,n30900);
  nand U32730(n30900,n30873,n30970);
  nand U32731(n30970,n30877,n30969);
  or U32732(n30969,n30879,n29197);
  not U32733(n30877,n30967);
  nand U32734(n30967,n30971,n30972);
  nand U32735(n30972,n30973,n29205);
  nand U32736(n30901,n29197,n30879);
  nand U32737(n30879,n30974,n30975,n30976,n30977);
  nor U32738(n30977,n30978,n30979);
  nor U32739(n30979,n29104,n29260);
  not U32740(n29104,G59319);
  nor U32741(n30978,n29261,n30885);
  nand U32742(n30976,n29197,n28535);
  nand U32743(n30975,n29264,n30980);
  xnor U32744(n30980,n28307,n30981);
  xnor U32745(n30981,n30912,n30915);
  and U32746(n30912,n30982,n30983);
  nand U32747(n30983,n30984,n30985,n28327);
  nand U32748(n30974,n28307,n29214);
  nand U32749(n30955,n29231,n28307);
  not U32750(n28307,n29102);
  nand U32751(n29102,n30986,n30918);
  nand U32752(n30918,n30987,n30988,n30989);
  xnor U32753(n30989,n30990,n29174);
  nand U32754(n30986,n30991,n30992);
  nand U32755(n30992,n30988,n30987);
  xnor U32756(n30991,n29226,n30990);
  nand U32757(n30990,n30993,n30994,n30995,n30996);
  nand U32758(n30996,n28535,n29288);
  not U32759(n28535,n28302);
  nand U32760(n28302,n30997,n30998);
  or U32761(n30998,n30869,n30999);
  nand U32762(n30869,n31000,n31001);
  nand U32763(n31001,n31002,n31003);
  nand U32764(n30997,n31004,n31003,n31002);
  nand U32765(n31002,n31005,n31006);
  nand U32766(n31004,n31000,n30870);
  not U32767(n30870,n30999);
  nor U32768(n30999,n27999,n30915,n31007);
  not U32769(n30915,n30914);
  nand U32770(n31000,n31007,n31008);
  nand U32771(n31008,n28576,n30914);
  nand U32772(n30914,n31009,n31010,n31011,n31012);
  nor U32773(n31012,n31013,n31014,n31015,n31016);
  nor U32774(n31016,n29760,n30622);
  nor U32775(n31015,n29759,n30623);
  nor U32776(n31014,n29758,n30624);
  nor U32777(n31013,n29752,n30625);
  nor U32778(n31011,n31017,n31018,n31019,n31020);
  nor U32779(n31020,n29751,n30630);
  nor U32780(n31019,n29750,n30631);
  nor U32781(n31018,n29744,n30632);
  nor U32782(n31017,n29743,n30633);
  nor U32783(n31010,n31021,n31022,n31023,n31024);
  nor U32784(n31024,n29742,n30638);
  nor U32785(n31023,n29736,n30639);
  nor U32786(n31022,n29735,n30640);
  nor U32787(n31021,n29734,n30641);
  nor U32788(n31009,n31025,n31026,n31027,n31028);
  nor U32789(n31028,n29761,n30646);
  nor U32790(n31027,n29753,n30647);
  nor U32791(n31026,n29745,n30648);
  nor U32792(n31025,n29737,n30649);
  xor U32793(n31007,n27993,n31029);
  nor U32794(n31029,n31030,n31031,n31032,n31033);
  and U32795(n31033,n29228,G59255);
  nor U32796(n31032,n29486,n30885);
  not U32797(n30885,G59128);
  and U32798(n31031,n29226,G59160);
  nor U32799(n31030,n31034,n28303);
  not U32800(n28303,G59287);
  nand U32801(n30995,G59128,n29287);
  nand U32802(n30994,G59319,n27993);
  nand U32803(n30993,G59160,n30080);
  nand U32804(G2522,n31035,n31036,n31037,n31038);
  nor U32805(n31038,n31039,n31040,n31041);
  nor U32806(n31041,G59127,n30882,n29185);
  nor U32807(n31040,n30962,n30884);
  and U32808(n30962,n29247,n31042);
  nand U32809(n31042,n29688,n30882);
  not U32810(n30882,n30964);
  nor U32811(n30964,n31043,n31044,n31045);
  nor U32812(n31039,n31046,n29192);
  nand U32813(n31037,n29193,n28539);
  nand U32814(n31036,n29194,n28316);
  nand U32815(n28316,n31047,n31048,n31049);
  or U32816(n31049,n30873,n31050);
  nand U32817(n30873,n29197,n31051);
  nand U32818(n31048,n31050,n30973,n29197);
  not U32819(n30973,n31051);
  nand U32820(n31047,n31052,n29205);
  xnor U32821(n31052,n31051,n31050);
  not U32822(n31050,n30971);
  nand U32823(n30971,n31053,n31054);
  nand U32824(n31054,n29197,n31055);
  or U32825(n31055,n31056,n31057);
  nand U32826(n31053,n31057,n31056);
  nand U32827(n31051,n31058,n31059,n31060,n31061);
  nor U32828(n31061,n31062,n31063);
  nor U32829(n31063,n31046,n29260);
  not U32830(n31046,G59318);
  nor U32831(n31062,n29261,n30884);
  not U32832(n30884,G59127);
  nand U32833(n31060,n29197,n28539);
  nand U32834(n31059,n29264,n31064);
  xor U32835(n31064,n31065,n31066);
  nand U32836(n31066,n28327,n30985);
  nand U32837(n31065,n30984,n30982);
  nand U32838(n30982,n28317,n31067);
  or U32839(n30984,n31067,n28317);
  nand U32840(n31058,n28317,n29214);
  nand U32841(n31035,n29231,n28317);
  xor U32842(n28317,n30988,n30987);
  xor U32843(n30987,n31068,n29226);
  nand U32844(n31068,n31069,n31070,n31071,n31072);
  nand U32845(n31072,n28539,n29288);
  not U32846(n28539,n28315);
  xnor U32847(n28315,n31006,n31073);
  and U32848(n31073,n31005,n31003);
  nand U32849(n31003,n31074,n31067,n28576);
  nand U32850(n31005,n31075,n31076,n31077);
  nand U32851(n31077,n28576,n31067);
  nand U32852(n31067,n31078,n31079,n31080,n31081);
  nor U32853(n31081,n31082,n31083,n31084,n31085);
  nor U32854(n31085,n29856,n30622);
  nor U32855(n31084,n29855,n30623);
  nor U32856(n31083,n29854,n30624);
  nor U32857(n31082,n29848,n30625);
  nor U32858(n31080,n31086,n31087,n31088,n31089);
  nor U32859(n31089,n29847,n30630);
  nor U32860(n31088,n29846,n30631);
  nor U32861(n31087,n29840,n30632);
  nor U32862(n31086,n29839,n30633);
  nor U32863(n31079,n31090,n31091,n31092,n31093);
  nor U32864(n31093,n29838,n30638);
  nor U32865(n31092,n29832,n30639);
  nor U32866(n31091,n29831,n30640);
  nor U32867(n31090,n29830,n30641);
  nor U32868(n31078,n31094,n31095,n31096,n31097);
  nor U32869(n31097,n29857,n30646);
  nor U32870(n31096,n29849,n30647);
  nor U32871(n31095,n29841,n30648);
  nor U32872(n31094,n29833,n30649);
  nand U32873(n31076,n31074,n28963);
  nand U32874(n31074,n31098,n31099,n31100);
  nand U32875(n31099,G59127,n29227);
  nand U32876(n31098,G59254,n29228);
  nand U32877(n31075,n31100,n27993);
  and U32878(n31100,n31101,n31102);
  nand U32879(n31102,G59286,n29225);
  nand U32880(n31101,G59159,n29226);
  nand U32881(n31006,n31103,n31104);
  nand U32882(n31104,n31105,n31106);
  not U32883(n31105,n31107);
  nand U32884(n31071,G59127,n29287);
  nand U32885(n31070,G59318,n27993);
  nand U32886(n31069,G59159,n30080);
  nand U32887(G2521,n31108,n31109,n31110,n31111);
  nor U32888(n31111,n31112,n31113,n31114);
  nor U32889(n31114,G59126,n29185,n31044,n31045);
  not U32890(n31044,G59125);
  nor U32891(n31113,n31115,n31043);
  nor U32892(n31115,n31116,n31117);
  nor U32893(n31116,G59125,n29185);
  nor U32894(n31112,n31118,n29192);
  nand U32895(n31110,n29193,n28543);
  nand U32896(n31109,n29194,n28326);
  xnor U32897(n28326,n31119,n31056);
  nand U32898(n31056,n31120,n31121,n31122,n31123);
  nor U32899(n31123,n31124,n31125);
  nor U32900(n31125,n31118,n29260);
  not U32901(n31118,G59317);
  nor U32902(n31124,n29261,n31043);
  not U32903(n31043,G59126);
  nand U32904(n31122,n29197,n28543);
  nand U32905(n31121,n31126,n29264);
  xor U32906(n31126,n28327,n30985);
  nand U32907(n31120,n28327,n29214);
  xnor U32908(n31119,n29197,n31057);
  nor U32909(n31057,n31127,n31128);
  nor U32910(n31127,n31129,n31130);
  nand U32911(n31108,n29231,n28327);
  nor U32912(n28327,n30988,n31131);
  and U32913(n31131,n31132,n31133);
  nor U32914(n30988,n31133,n31132);
  xor U32915(n31132,n31134,n29174);
  nand U32916(n31134,n31135,n31136,n31137,n31138);
  nand U32917(n31138,n28543,n29288);
  xor U32918(n28543,n31139,n31107);
  nand U32919(n31139,n31103,n31106);
  nand U32920(n31106,n31140,n31141,n31142);
  nand U32921(n31142,n28576,n30985);
  nand U32922(n31141,n31143,n27993);
  nand U32923(n31140,n31144,n28963);
  nand U32924(n31103,n31144,n30985,n28576);
  nand U32925(n30985,n31145,n31146,n31147,n31148);
  nor U32926(n31148,n31149,n31150,n31151,n31152);
  nor U32927(n31152,n29913,n30639);
  nand U32928(n30639,n31153,n31154);
  nor U32929(n31151,n29915,n30649);
  nand U32930(n30649,n31153,n31155);
  nor U32931(n31150,n29927,n30648);
  nand U32932(n30648,n31156,n31155);
  nor U32933(n31149,n29937,n30647);
  nand U32934(n30647,n31157,n31155);
  nor U32935(n31147,n31158,n31159,n31160,n31161);
  nor U32936(n31161,n29926,n30632);
  nand U32937(n30632,n31156,n31154);
  nor U32938(n31160,n29933,n30631);
  nand U32939(n30631,n31157,n31162);
  nor U32940(n31159,n29908,n30641);
  nand U32941(n30641,n31153,n31162);
  nor U32942(n31158,n29911,n30640);
  nand U32943(n30640,n31153,n31163);
  nor U32944(n31153,n31164,n31165);
  nor U32945(n31146,n31166,n31167,n31168,n31169);
  nor U32946(n31169,n29936,n30625);
  nand U32947(n30625,n31157,n31154);
  nor U32948(n31168,n29942,n30624);
  nand U32949(n30624,n31170,n31162);
  nor U32950(n31167,n29946,n30623);
  nand U32951(n30623,n31170,n31163);
  nor U32952(n31166,n29925,n30633);
  nand U32953(n30633,n31156,n31163);
  nor U32954(n31145,n31171,n31172,n31173,n31174);
  nor U32955(n31174,n29949,n30646);
  nand U32956(n30646,n31170,n31155);
  nor U32957(n31173,n29947,n30622);
  nand U32958(n30622,n31170,n31154);
  nor U32959(n31170,n31175,n31176);
  nor U32960(n31172,n29935,n30630);
  nand U32961(n30630,n31157,n31163);
  nor U32962(n31157,n31176,n31164);
  not U32963(n31164,n31175);
  nor U32964(n31171,n29923,n30638);
  nand U32965(n30638,n31156,n31162);
  nor U32966(n31156,n31175,n31165);
  not U32967(n31165,n31176);
  nand U32968(n31176,n31177,n31178,n31179);
  not U32969(n31179,n31180);
  nand U32970(n31178,G59109,n31181);
  nand U32971(n31177,n31182,G59111);
  xnor U32972(n31175,G59110,n31181);
  nand U32973(n31144,n31183,n31184,n31143);
  and U32974(n31143,n31185,n31186);
  nand U32975(n31186,G59285,n29225);
  nand U32976(n31185,G59158,n29226);
  nand U32977(n31184,G59126,n29227);
  nand U32978(n31183,G59253,n29228);
  nand U32979(n31137,G59126,n29287);
  nand U32980(n31136,G59317,n27993);
  nand U32981(n31135,G59158,n30080);
  or U32982(n31133,n31187,n31188);
  nand U32983(G2520,n31189,n31190,n31191,n31192);
  nor U32984(n31192,n31193,n31194,n31195);
  nor U32985(n31195,G59125,n31045,n29185);
  and U32986(n31194,n31117,G59125);
  nand U32987(n31117,n29247,n31196);
  nand U32988(n31196,n29688,n31045);
  or U32989(n31045,n31197,n31198);
  nor U32990(n31193,n31199,n29192);
  not U32991(n31199,G59316);
  nand U32992(n31191,n29193,n28547);
  nand U32993(n31190,n29194,n28336);
  xor U32994(n28336,n31129,n31200);
  nor U32995(n31200,n31130,n31128);
  nor U32996(n31128,n31201,n31202);
  and U32997(n31130,n31202,n31201);
  nand U32998(n31201,n31203,n31204,n31205,n31206);
  nand U32999(n31206,n31207,n28337);
  nand U33000(n31205,n28547,n29197);
  nand U33001(n31204,G59125,n29229);
  nand U33002(n31203,n29230,G59316);
  xnor U33003(n31202,n29205,n31208);
  nand U33004(n31208,n31209,n31210,n31211,n31212);
  nand U33005(n31212,n31213,n31214,n31215,n31216);
  nor U33006(n31216,n31217,n31218,n31219,n31220);
  nor U33007(n31220,n29347,n31221);
  nor U33008(n31219,n29979,n31222);
  nor U33009(n31218,n29335,n31223);
  nand U33010(n31217,n31224,n31225);
  nand U33011(n31225,n31226,G58996);
  nand U33012(n31224,n31227,G58988);
  nor U33013(n31215,n31228,n31229,n31230,n31231);
  nor U33014(n31231,n29345,n31232);
  nor U33015(n31230,n29973,n31233);
  nor U33016(n31229,n29967,n31234);
  nor U33017(n31228,n29329,n31235);
  nor U33018(n31214,n31236,n31237,n31238,n31239);
  nor U33019(n31239,n29977,n31240);
  nor U33020(n31238,n29975,n31241);
  nor U33021(n31237,n29341,n31242);
  nor U33022(n31236,n29343,n31243);
  nor U33023(n31213,n31244,n31245,n31246,n29205);
  nor U33024(n31246,n29963,n31247);
  nor U33025(n31245,n29965,n31248);
  nor U33026(n31244,n29961,n31249);
  nand U33027(n31211,n31250,n29881);
  nand U33028(n29881,n31251,n31252,n31253,n31254);
  nor U33029(n31254,n31255,n31256,n31257,n31258);
  nor U33030(n31258,n29965,n31259);
  nor U33031(n31257,n29963,n31260);
  nor U33032(n31256,n29961,n31261);
  nor U33033(n31255,n29977,n31262);
  nor U33034(n31253,n31263,n31264,n31265,n31266);
  nor U33035(n31266,n29975,n31267);
  nor U33036(n31265,n29973,n31268);
  nor U33037(n31264,n29345,n31269);
  nor U33038(n31263,n29343,n31270);
  nor U33039(n31252,n31271,n31272,n31273,n31274);
  nor U33040(n31274,n29341,n31275);
  nor U33041(n31273,n29333,n31276);
  nor U33042(n31272,n29331,n31277);
  nor U33043(n31271,n29329,n31278);
  nor U33044(n31251,n31279,n31280,n31281,n31282);
  nor U33045(n31282,n29967,n31283);
  nor U33046(n31281,n29979,n31284);
  nor U33047(n31280,n29347,n31285);
  nor U33048(n31279,n29335,n31286);
  nand U33049(n31210,n29264,n31287);
  nand U33050(n31287,n31288,n31289,n31290,n31291);
  nor U33051(n31291,n31292,n31293,n31294,n31295);
  nor U33052(n31295,n29967,n31296);
  nor U33053(n31294,n29965,n31297);
  nor U33054(n31293,n29963,n31298);
  nor U33055(n31292,n29961,n31299);
  nor U33056(n31290,n31300,n31301,n31302,n31303);
  nor U33057(n31303,n29979,n31304);
  nor U33058(n31302,n29977,n31305);
  nor U33059(n31301,n29975,n31306);
  nor U33060(n31300,n29973,n31307);
  nor U33061(n31289,n31308,n31309,n31310,n31311);
  nor U33062(n31311,n29347,n31312);
  nor U33063(n31310,n29345,n31313);
  nor U33064(n31309,n29343,n31314);
  nor U33065(n31308,n29341,n31315);
  nor U33066(n31288,n31316,n31317,n31318,n31319);
  nor U33067(n31319,n29335,n31320);
  nor U33068(n31318,n29333,n31321);
  nor U33069(n31317,n29331,n31322);
  nor U33070(n31316,n29329,n31323);
  nand U33071(n31209,n31324,n31325);
  nand U33072(n31129,n31326,n31327);
  nand U33073(n31189,n29231,n28337);
  nand U33074(n28337,n31328,n31329);
  nand U33075(n31329,n31330,n31331);
  or U33076(n31330,n31188,n31332);
  not U33077(n31188,n31333);
  nand U33078(n31328,n31187,n31333);
  nand U33079(n31333,n31334,n31335);
  nand U33080(n31335,n28576,G59100);
  nor U33081(n31187,n31331,n31332);
  nor U33082(n31332,n29967,n31334,n27999);
  nor U33083(n31334,n31336,n31337);
  and U33084(n31337,n31338,n29174);
  nor U33085(n31336,n31338,n28547,n29174);
  not U33086(n28547,n28335);
  nand U33087(n28335,n31107,n31339);
  nand U33088(n31339,n31340,n31341);
  xnor U33089(n31340,n28963,n31342);
  nand U33090(n31107,n31343,n31344);
  xnor U33091(n31343,n27993,n31342);
  and U33092(n31342,n31345,n31346,n31347,n31348);
  nand U33093(n31348,G59284,n29225);
  nand U33094(n31347,G59157,n29226);
  nand U33095(n31346,G59125,n29227);
  nand U33096(n31345,G59252,n29228);
  nand U33097(n31338,n31349,n31350,n31351);
  nand U33098(n31351,G59157,n30080);
  nand U33099(n31350,G59125,n29287);
  nand U33100(n31349,G59316,n27993);
  or U33101(n31331,n31352,n31353);
  and U33102(n31353,n31354,n31355);
  nand U33103(G2519,n31356,n31357,n31358,n31359);
  nor U33104(n31359,n31360,n31361,n31362);
  nor U33105(n31362,n28345,n29685);
  and U33106(n31361,n28348,n29231);
  nor U33107(n31360,n31363,n29192);
  not U33108(n31363,G59315);
  nand U33109(n31358,n29194,n28734);
  not U33110(n28734,n28347);
  nand U33111(n28347,n31364,n31365);
  nand U33112(n31365,n31366,n31367,n31368);
  nand U33113(n31366,n31369,n31326);
  nand U33114(n31364,n31370,n31326);
  nand U33115(n31326,n31371,n31372);
  xnor U33116(n31371,n31373,n29205);
  not U33117(n31370,n31327);
  nand U33118(n31327,n31369,n31374);
  nand U33119(n31374,n31368,n31367);
  nand U33120(n31368,n31375,n31376);
  nand U33121(n31369,n31377,n31378);
  xnor U33122(n31378,n29197,n31373);
  nand U33123(n31373,n31379,n31380,n31381,n31382);
  nand U33124(n31382,n31383,n31384,n31385,n31386);
  nor U33125(n31386,n31387,n31388,n31389,n31390);
  nor U33126(n31390,n29417,n31221);
  nor U33127(n31389,n29428,n31222);
  nor U33128(n31388,n29409,n31223);
  nand U33129(n31387,n31391,n31392);
  nand U33130(n31392,n31226,G58997);
  nand U33131(n31391,n31227,G58989);
  nor U33132(n31385,n31393,n31394,n31395,n31396);
  nor U33133(n31396,n29416,n31232);
  nor U33134(n31395,n29422,n31233);
  nor U33135(n31394,n29440,n31234);
  nor U33136(n31393,n29406,n31235);
  nor U33137(n31384,n31397,n31398,n31399,n31400);
  nor U33138(n31400,n29426,n31240);
  nor U33139(n31399,n29424,n31241);
  nor U33140(n31398,n29414,n31242);
  nor U33141(n31397,n29415,n31243);
  nor U33142(n31383,n31401,n31402,n31403,n29205);
  nor U33143(n31403,n29436,n31247);
  nor U33144(n31402,n29438,n31248);
  nor U33145(n31401,n29434,n31249);
  nand U33146(n31381,n31250,n30035);
  nand U33147(n30035,n31404,n31405,n31406,n31407);
  nor U33148(n31407,n31408,n31409,n31410,n31411);
  nor U33149(n31411,n29438,n31259);
  nor U33150(n31410,n29436,n31260);
  nor U33151(n31409,n29434,n31261);
  nor U33152(n31408,n29426,n31262);
  nor U33153(n31406,n31412,n31413,n31414,n31415);
  nor U33154(n31415,n29424,n31267);
  nor U33155(n31414,n29422,n31268);
  nor U33156(n31413,n29416,n31269);
  nor U33157(n31412,n29415,n31270);
  nor U33158(n31405,n31416,n31417,n31418,n31419);
  nor U33159(n31419,n29414,n31275);
  nor U33160(n31418,n29408,n31276);
  nor U33161(n31417,n29407,n31277);
  nor U33162(n31416,n29406,n31278);
  nor U33163(n31404,n31420,n31421,n31422,n31423);
  nor U33164(n31423,n29440,n31283);
  nor U33165(n31422,n29428,n31284);
  nor U33166(n31421,n29417,n31285);
  nor U33167(n31420,n29409,n31286);
  nand U33168(n31380,n31324,n31424);
  nand U33169(n31424,n31425,n31426,n31427,n31428);
  nor U33170(n31428,n31429,n31430,n31431,n31432);
  nor U33171(n31432,n29436,n31433);
  nor U33172(n31431,n29434,n31434);
  nor U33173(n31430,n29428,n31435);
  nor U33174(n31429,n29424,n31436);
  nor U33175(n31427,n31437,n31438,n31439,n31440);
  nor U33176(n31440,n29422,n31441);
  nor U33177(n31439,n29417,n31442);
  nor U33178(n31438,n29415,n31443);
  nor U33179(n31437,n29414,n31444);
  nor U33180(n31426,n31445,n31446,n31447,n31448);
  nor U33181(n31448,n29409,n31449);
  nor U33182(n31447,n29407,n31450);
  nor U33183(n31446,n29406,n31451);
  nor U33184(n31445,n29440,n31452);
  nor U33185(n31425,n31453,n31454,n31455,n31456);
  nor U33186(n31456,n29438,n31457);
  nor U33187(n31455,n29426,n31458);
  nor U33188(n31454,n29416,n31459);
  nor U33189(n31453,n29408,n31460);
  nand U33190(n31379,n29264,n31461);
  nand U33191(n31461,n31462,n31463,n31464,n31465);
  nor U33192(n31465,n31466,n31467,n31468,n31469);
  nor U33193(n31469,n29440,n31296);
  nor U33194(n31468,n29438,n31297);
  nor U33195(n31467,n29436,n31298);
  nor U33196(n31466,n29434,n31299);
  nor U33197(n31464,n31470,n31471,n31472,n31473);
  nor U33198(n31473,n29428,n31304);
  nor U33199(n31472,n29426,n31305);
  nor U33200(n31471,n29424,n31306);
  nor U33201(n31470,n29422,n31307);
  nor U33202(n31463,n31474,n31475,n31476,n31477);
  nor U33203(n31477,n29417,n31312);
  nor U33204(n31476,n29416,n31313);
  nor U33205(n31475,n29415,n31314);
  nor U33206(n31474,n29414,n31315);
  nor U33207(n31462,n31478,n31479,n31480,n31481);
  nor U33208(n31481,n29409,n31320);
  nor U33209(n31480,n29408,n31321);
  nor U33210(n31479,n29407,n31322);
  nor U33211(n31478,n29406,n31323);
  not U33212(n31377,n31372);
  nand U33213(n31372,n31482,n31483,n31484,n31485);
  nand U33214(n31485,n28348,n31207);
  xor U33215(n28348,n31355,n31486);
  nor U33216(n31486,n31352,n31487);
  not U33217(n31487,n31354);
  nand U33218(n31354,n31488,n31489);
  nand U33219(n31489,n28576,G59101);
  nor U33220(n31352,n27999,n29440,n31488);
  xor U33221(n31488,n31490,n29174);
  nand U33222(n31490,n31491,n31492,n31493,n31494);
  nand U33223(n31494,n28551,n29288);
  nand U33224(n31493,G59124,n29287);
  nand U33225(n31492,G59315,n27993);
  nand U33226(n31491,G59156,n30080);
  nand U33227(n31355,n31495,n31496);
  nand U33228(n31496,n31497,n31498);
  nand U33229(n31497,n31499,n31500);
  nand U33230(n31500,n28576,G59102);
  not U33231(n31495,n31501);
  nand U33232(n31484,n29197,n28551);
  not U33233(n28551,n28345);
  nand U33234(n28345,n31341,n31502);
  nand U33235(n31502,n31503,n31504);
  not U33236(n31341,n31344);
  nor U33237(n31344,n31504,n31503);
  xor U33238(n31503,n27993,n31505);
  nor U33239(n31505,n31506,n31507,n31508,n31509);
  and U33240(n31509,n29228,G59251);
  and U33241(n31508,n29227,G59124);
  nor U33242(n31507,n29174,n29131);
  not U33243(n29131,G59156);
  nor U33244(n31506,n31034,n28346);
  not U33245(n28346,G59283);
  nand U33246(n31483,G59124,n29229);
  nand U33247(n31482,n29230,G59315);
  nand U33248(n31357,n31510,n31198,n29688);
  nand U33249(n31198,G59124,n27943);
  nand U33250(n31356,G59124,n31511);
  nand U33251(n31511,n29247,n31512);
  nand U33252(n31512,n29688,n31197);
  not U33253(n31197,n31510);
  nor U33254(n31510,n31513,n31514,n31515);
  nand U33255(G2518,n31516,n31517,n31518,n31519);
  nor U33256(n31519,n31520,n31521,n31522);
  nor U33257(n31522,G59123,n29185,n31514,n31515);
  nor U33258(n31521,n31523,n31513);
  nor U33259(n31523,n31524,n29190);
  nor U33260(n31524,n31525,n29185);
  nor U33261(n31525,n31514,n31515);
  nor U33262(n31520,n31526,n29192);
  not U33263(n31526,G59314);
  nand U33264(n31518,n29193,n28555);
  nand U33265(n31517,n29194,n28359);
  xor U33266(n28359,n31376,n31527);
  and U33267(n31527,n31375,n31367);
  nand U33268(n31367,n31528,n31529);
  or U33269(n31375,n31529,n31528);
  xnor U33270(n31528,n31530,n29205);
  nand U33271(n31530,n31531,n31532,n31533,n31534);
  nand U33272(n31534,n31535,n31536,n31537,n31538);
  nor U33273(n31538,n31539,n31540,n31541,n31542);
  nor U33274(n31542,n29521,n31221);
  nor U33275(n31541,n30148,n31222);
  nor U33276(n31540,n29513,n31223);
  nand U33277(n31539,n31543,n31544);
  nand U33278(n31544,n31226,G58998);
  nand U33279(n31543,n31227,G58990);
  nor U33280(n31537,n31545,n31546,n31547,n31548);
  nor U33281(n31548,n29520,n31232);
  nor U33282(n31547,n30145,n31233);
  nor U33283(n31546,n30140,n31234);
  nor U33284(n31545,n29510,n31235);
  nor U33285(n31536,n31549,n31550,n31551,n31552);
  nor U33286(n31552,n30147,n31240);
  nor U33287(n31551,n30146,n31241);
  nor U33288(n31550,n29518,n31242);
  nor U33289(n31549,n29519,n31243);
  nor U33290(n31535,n31553,n31554,n31555,n29205);
  nor U33291(n31555,n30138,n31247);
  nor U33292(n31554,n30139,n31248);
  nor U33293(n31553,n30137,n31249);
  nand U33294(n31533,n31250,n30115);
  nand U33295(n30115,n31556,n31557,n31558,n31559);
  nor U33296(n31559,n31560,n31561,n31562,n31563);
  nor U33297(n31563,n30139,n31259);
  nor U33298(n31562,n30138,n31260);
  nor U33299(n31561,n30137,n31261);
  nor U33300(n31560,n30147,n31262);
  nor U33301(n31558,n31564,n31565,n31566,n31567);
  nor U33302(n31567,n30146,n31267);
  nor U33303(n31566,n30145,n31268);
  nor U33304(n31565,n29520,n31269);
  nor U33305(n31564,n29519,n31270);
  nor U33306(n31557,n31568,n31569,n31570,n31571);
  nor U33307(n31571,n29518,n31275);
  nor U33308(n31570,n29512,n31276);
  nor U33309(n31569,n29511,n31277);
  nor U33310(n31568,n29510,n31278);
  nor U33311(n31556,n31572,n31573,n31574,n31575);
  nor U33312(n31575,n30140,n31283);
  nor U33313(n31574,n30148,n31284);
  nor U33314(n31573,n29521,n31285);
  nor U33315(n31572,n29513,n31286);
  nand U33316(n31532,n31324,n31576);
  nand U33317(n31576,n31577,n31578,n31579,n31580);
  nor U33318(n31580,n31581,n31582,n31583,n31584);
  nor U33319(n31584,n30138,n31433);
  nor U33320(n31583,n30137,n31434);
  nor U33321(n31582,n30148,n31435);
  nor U33322(n31581,n30146,n31436);
  nor U33323(n31579,n31585,n31586,n31587,n31588);
  nor U33324(n31588,n30145,n31441);
  nor U33325(n31587,n29521,n31442);
  nor U33326(n31586,n29519,n31443);
  nor U33327(n31585,n29518,n31444);
  nor U33328(n31578,n31589,n31590,n31591,n31592);
  nor U33329(n31592,n29513,n31449);
  nor U33330(n31591,n29511,n31450);
  nor U33331(n31590,n29510,n31451);
  nor U33332(n31589,n30140,n31452);
  nor U33333(n31577,n31593,n31594,n31595,n31596);
  nor U33334(n31596,n30139,n31457);
  nor U33335(n31595,n30147,n31458);
  nor U33336(n31594,n29520,n31459);
  nor U33337(n31593,n29512,n31460);
  nand U33338(n31531,n29264,n31597);
  nand U33339(n31597,n31598,n31599,n31600,n31601);
  nor U33340(n31601,n31602,n31603,n31604,n31605);
  nor U33341(n31605,n30140,n31296);
  nor U33342(n31604,n30139,n31297);
  nor U33343(n31603,n30138,n31298);
  nor U33344(n31602,n30137,n31299);
  nor U33345(n31600,n31606,n31607,n31608,n31609);
  nor U33346(n31609,n30148,n31304);
  nor U33347(n31608,n30147,n31305);
  nor U33348(n31607,n30146,n31306);
  nor U33349(n31606,n30145,n31307);
  nor U33350(n31599,n31610,n31611,n31612,n31613);
  nor U33351(n31613,n29521,n31312);
  nor U33352(n31612,n29520,n31313);
  nor U33353(n31611,n29519,n31314);
  nor U33354(n31610,n29518,n31315);
  nor U33355(n31598,n31614,n31615,n31616,n31617);
  nor U33356(n31617,n29513,n31320);
  nor U33357(n31616,n29512,n31321);
  nor U33358(n31615,n29511,n31322);
  nor U33359(n31614,n29510,n31323);
  nand U33360(n31529,n31618,n31619,n31620,n31621);
  nand U33361(n31621,n28360,n31207);
  nand U33362(n31620,n28555,n29197);
  nand U33363(n31619,G59123,n29229);
  nand U33364(n31618,n29230,G59314);
  nand U33365(n31376,n31622,n31623);
  nand U33366(n31623,n31624,n31625);
  nand U33367(n31624,n31626,n31627);
  or U33368(n31622,n31627,n31626);
  xor U33369(n28360,n31498,n31628);
  nor U33370(n31628,n31629,n31501);
  nor U33371(n31501,n30140,n31499,n27999);
  nor U33372(n31629,n31630,n31631);
  not U33373(n31631,n31499);
  nor U33374(n31499,n31632,n31633);
  and U33375(n31633,n31634,n29174);
  nor U33376(n31632,n31634,n28555,n29174);
  not U33377(n28555,n28356);
  nand U33378(n28356,n31504,n31635);
  nand U33379(n31635,n31636,n31637);
  or U33380(n31504,n31637,n31636);
  xor U33381(n31636,n27993,n31638);
  nor U33382(n31638,n31639,n31640,n31641,n31642);
  and U33383(n31642,n29228,G59250);
  nor U33384(n31641,n29486,n31513);
  not U33385(n31513,G59123);
  nor U33386(n31640,n29174,n29138);
  not U33387(n29138,G59155);
  nor U33388(n31639,n31034,n28357);
  not U33389(n28357,G59282);
  nand U33390(n31637,n31643,n31644);
  nand U33391(n31634,n31645,n31646,n31647);
  nand U33392(n31647,G59155,n30080);
  nand U33393(n31646,G59123,n29287);
  nand U33394(n31645,G59314,n27993);
  nor U33395(n31630,n30140,n27999);
  nand U33396(n31498,n31648,n31649);
  nand U33397(n31649,n31650,n31651);
  nand U33398(G2517,n31652,n31653,n31654,n31655);
  nor U33399(n31655,n31656,n31657,n31658);
  nor U33400(n31658,G59122,n31515,n29185);
  not U33401(n31515,n31659);
  nor U33402(n31657,n31660,n31514);
  nor U33403(n31660,n31661,n29190);
  nor U33404(n31661,n31659,n29185);
  nor U33405(n31659,n31662,n31663);
  nor U33406(n31656,n31664,n29192);
  nand U33407(n31653,n29194,n28371);
  xor U33408(n28371,n31665,n31627);
  xor U33409(n31627,n31666,n29205);
  nand U33410(n31666,n31667,n31668,n31669,n31670);
  nor U33411(n31670,n31671,n31672);
  nor U33412(n31672,n28691,n31673);
  and U33413(n31671,n30191,n31250);
  nand U33414(n30191,n31674,n31675,n31676,n31677);
  nor U33415(n31677,n31678,n31679,n31680,n31681);
  nor U33416(n31681,n30220,n31259);
  nor U33417(n31680,n30219,n31260);
  nor U33418(n31679,n30218,n31261);
  nor U33419(n31678,n30228,n31262);
  nor U33420(n31676,n31682,n31683,n31684,n31685);
  nor U33421(n31685,n30227,n31267);
  nor U33422(n31684,n30226,n31268);
  nor U33423(n31683,n29599,n31269);
  nor U33424(n31682,n29598,n31270);
  nor U33425(n31675,n31686,n31687,n31688,n31689);
  nor U33426(n31689,n29597,n31275);
  nor U33427(n31688,n29591,n31276);
  nor U33428(n31687,n29590,n31277);
  nor U33429(n31686,n29589,n31278);
  nor U33430(n31674,n31690,n31691,n31692,n31693);
  nor U33431(n31693,n30221,n31283);
  nor U33432(n31692,n30229,n31284);
  nor U33433(n31691,n29600,n31285);
  nor U33434(n31690,n29592,n31286);
  nand U33435(n31669,n29264,n31694);
  nand U33436(n31694,n31695,n31696,n31697,n31698);
  nor U33437(n31698,n31699,n31700,n31701,n31702);
  nor U33438(n31702,n30221,n31296);
  nor U33439(n31701,n30220,n31297);
  nor U33440(n31700,n30219,n31298);
  nor U33441(n31699,n30218,n31299);
  nor U33442(n31697,n31703,n31704,n31705,n31706);
  nor U33443(n31706,n30229,n31304);
  nor U33444(n31705,n30228,n31305);
  nor U33445(n31704,n30227,n31306);
  nor U33446(n31703,n30226,n31307);
  nor U33447(n31696,n31707,n31708,n31709,n31710);
  nor U33448(n31710,n29600,n31312);
  nor U33449(n31709,n29599,n31313);
  nor U33450(n31708,n29598,n31314);
  nor U33451(n31707,n29597,n31315);
  nor U33452(n31695,n31711,n31712,n31713,n31714);
  nor U33453(n31714,n29592,n31320);
  nor U33454(n31713,n29591,n31321);
  nor U33455(n31712,n29590,n31322);
  nor U33456(n31711,n29589,n31323);
  nand U33457(n31668,n31715,n31716,n31717,n31718);
  nor U33458(n31718,n31719,n31720,n31721,n31722);
  nor U33459(n31722,n29600,n31221);
  nor U33460(n31721,n30229,n31222);
  nor U33461(n31720,n29592,n31223);
  nand U33462(n31719,n31723,n31724);
  nand U33463(n31724,n31226,G58999);
  nand U33464(n31723,n31227,G58991);
  nor U33465(n31717,n31725,n31726,n31727,n31728);
  nor U33466(n31728,n29599,n31232);
  nor U33467(n31727,n30226,n31233);
  nor U33468(n31726,n30221,n31234);
  nor U33469(n31725,n29589,n31235);
  nor U33470(n31716,n31729,n31730,n31731,n31732);
  nor U33471(n31732,n30228,n31240);
  nor U33472(n31731,n30227,n31241);
  nor U33473(n31730,n29597,n31242);
  nor U33474(n31729,n29598,n31243);
  nor U33475(n31715,n31733,n31734,n31735,n29205);
  nor U33476(n31735,n30219,n31247);
  nor U33477(n31734,n30220,n31248);
  nor U33478(n31733,n30218,n31249);
  nand U33479(n31667,n31324,n31736);
  nand U33480(n31736,n31737,n31738,n31739,n31740);
  nor U33481(n31740,n31741,n31742,n31743,n31744);
  nor U33482(n31744,n30219,n31433);
  nor U33483(n31743,n30218,n31434);
  nor U33484(n31742,n30229,n31435);
  nor U33485(n31741,n30227,n31436);
  nor U33486(n31739,n31745,n31746,n31747,n31748);
  nor U33487(n31748,n30226,n31441);
  nor U33488(n31747,n29600,n31442);
  nor U33489(n31746,n29598,n31443);
  nor U33490(n31745,n29597,n31444);
  nor U33491(n31738,n31749,n31750,n31751,n31752);
  nor U33492(n31752,n29592,n31449);
  nor U33493(n31751,n29590,n31450);
  nor U33494(n31750,n29589,n31451);
  nor U33495(n31749,n30221,n31452);
  nor U33496(n31737,n31753,n31754,n31755,n31756);
  nor U33497(n31756,n30220,n31457);
  nor U33498(n31755,n30228,n31458);
  nor U33499(n31754,n29599,n31459);
  nor U33500(n31753,n29591,n31460);
  xor U33501(n31665,n31625,n31626);
  and U33502(n31626,n31757,n31758,n31759,n31760);
  nand U33503(n31760,n27871,n31207);
  nand U33504(n31759,G59122,n29229);
  nand U33505(n31758,n29197,n28559);
  nand U33506(n31757,n29230,G59313);
  nand U33507(n31625,n31761,n31762);
  nand U33508(n31762,n31763,n31764);
  nand U33509(n31652,n29193,n28559);
  nand U33510(G2516,n31765,n31766,n31767,n31768);
  nor U33511(n31768,n31769,n31770,n31771);
  nor U33512(n31771,G59121,n31662,n29185);
  nor U33513(n31770,n31772,n31663);
  nor U33514(n31772,n31773,n29190);
  and U33515(n31773,n31662,n29688);
  nand U33516(n31662,n27943,n31774);
  nand U33517(n31774,n31775,n31776);
  nor U33518(n31769,n28382,n29192);
  nand U33519(n31766,n29194,n28384);
  xor U33520(n28384,n31764,n31777);
  and U33521(n31777,n31761,n31763);
  or U33522(n31763,n31778,n31779);
  nand U33523(n31761,n31779,n31778);
  nand U33524(n31778,n31780,n31781,n31782,n31783);
  nand U33525(n31783,n27881,n31207);
  nand U33526(n31782,G59121,n29229);
  nand U33527(n31781,n29197,n28383);
  nand U33528(n31780,n29230,G59312);
  xnor U33529(n31779,n29205,n31784);
  nand U33530(n31784,n31785,n31786,n31787,n31788);
  nor U33531(n31788,n31789,n31790);
  nor U33532(n31790,n28691,n31791);
  nor U33533(n31789,n31792,n28761);
  nor U33534(n31792,n31793,n31794,n31795,n31796);
  nand U33535(n31796,n31797,n31798,n31799,n31800);
  nand U33536(n31800,n31801,G58984);
  nand U33537(n31799,n31802,G58992);
  nand U33538(n31798,n31803,G59000);
  nand U33539(n31797,n31804,G59008);
  nand U33540(n31795,n31805,n31806,n31807,n31808);
  nand U33541(n31808,n31809,G59016);
  nand U33542(n31807,n31810,G59024);
  nand U33543(n31806,n31811,G59032);
  nand U33544(n31805,n31812,G59040);
  nand U33545(n31794,n31813,n31814,n31815,n31816);
  nand U33546(n31816,n31817,G59048);
  nand U33547(n31815,n31818,G59056);
  nand U33548(n31814,n31819,G59064);
  nand U33549(n31813,n31820,G59072);
  nand U33550(n31793,n31821,n31822,n31823,n31824);
  nand U33551(n31824,n31825,G59080);
  nand U33552(n31823,n31826,G59088);
  nand U33553(n31822,n31827,G59096);
  nand U33554(n31821,n31828,G59104);
  nand U33555(n31787,n31250,n30275);
  nand U33556(n30275,n31829,n31830,n31831,n31832);
  nor U33557(n31832,n31833,n31834,n31835,n31836);
  nor U33558(n31836,n30304,n31259);
  nor U33559(n31835,n30303,n31260);
  nor U33560(n31834,n30302,n31261);
  nor U33561(n31833,n30312,n31262);
  nor U33562(n31831,n31837,n31838,n31839,n31840);
  nor U33563(n31840,n30311,n31267);
  nor U33564(n31839,n30310,n31268);
  nor U33565(n31838,n29675,n31269);
  nor U33566(n31837,n29674,n31270);
  nor U33567(n31830,n31841,n31842,n31843,n31844);
  nor U33568(n31844,n29673,n31275);
  nor U33569(n31843,n29667,n31276);
  nor U33570(n31842,n29666,n31277);
  nor U33571(n31841,n29665,n31278);
  nor U33572(n31829,n31845,n31846,n31847,n31848);
  nor U33573(n31848,n30305,n31283);
  nor U33574(n31847,n30313,n31284);
  nor U33575(n31846,n29676,n31285);
  nor U33576(n31845,n29668,n31286);
  nand U33577(n31786,n31849,n31850,n31851,n31852);
  nor U33578(n31852,n31853,n31854,n31855,n31856);
  nor U33579(n31856,n29676,n31221);
  nor U33580(n31855,n30313,n31222);
  nor U33581(n31854,n29668,n31223);
  nand U33582(n31853,n31857,n31858);
  nand U33583(n31858,n31226,G59000);
  nand U33584(n31857,n31227,G58992);
  nor U33585(n31851,n31859,n31860,n31861,n31862);
  nor U33586(n31862,n29675,n31232);
  nor U33587(n31861,n30310,n31233);
  nor U33588(n31860,n30305,n31234);
  nor U33589(n31859,n29665,n31235);
  nor U33590(n31850,n31863,n31864,n31865,n31866);
  nor U33591(n31866,n30312,n31240);
  nor U33592(n31865,n30311,n31241);
  nor U33593(n31864,n29673,n31242);
  nor U33594(n31863,n29674,n31243);
  nor U33595(n31849,n31867,n31868,n31869,n29205);
  nor U33596(n31869,n30303,n31247);
  nor U33597(n31868,n30304,n31248);
  nor U33598(n31867,n30302,n31249);
  nand U33599(n31785,n31324,n31870);
  nand U33600(n31870,n31871,n31872,n31873,n31874);
  nor U33601(n31874,n31875,n31876,n31877,n31878);
  nor U33602(n31878,n30303,n31433);
  nor U33603(n31877,n30302,n31434);
  nor U33604(n31876,n30313,n31435);
  nor U33605(n31875,n30311,n31436);
  nor U33606(n31873,n31879,n31880,n31881,n31882);
  nor U33607(n31882,n30310,n31441);
  nor U33608(n31881,n29676,n31442);
  nor U33609(n31880,n29674,n31443);
  nor U33610(n31879,n29673,n31444);
  nor U33611(n31872,n31883,n31884,n31885,n31886);
  nor U33612(n31886,n29668,n31449);
  nor U33613(n31885,n29666,n31450);
  nor U33614(n31884,n29665,n31451);
  nor U33615(n31883,n30305,n31452);
  nor U33616(n31871,n31887,n31888,n31889,n31890);
  nor U33617(n31890,n30304,n31457);
  nor U33618(n31889,n30312,n31458);
  nor U33619(n31888,n29675,n31459);
  nor U33620(n31887,n29667,n31460);
  nand U33621(n31764,n31891,n31892);
  nand U33622(n31892,n31893,n31894);
  nand U33623(n31765,n29193,n28383);
  nand U33624(G2515,n31895,n31896,n31897,n31898);
  nor U33625(n31898,n31899,n31900,n31901);
  and U33626(n31901,n31775,n31776,n29688);
  not U33627(n29688,n29185);
  nor U33628(n31900,n31902,n31775);
  nor U33629(n31902,n31903,n29190);
  nor U33630(n31903,n29185,n31776);
  nand U33631(n31776,G59118,n27943,G59119);
  nor U33632(n31899,n28394,n29192);
  not U33633(n28394,G59311);
  nand U33634(n31896,n29194,n28396);
  xor U33635(n28396,n31893,n31904);
  and U33636(n31904,n31894,n31891);
  nand U33637(n31891,n31905,n31906);
  nand U33638(n31906,n31907,n31908);
  nand U33639(n31894,n31907,n31908,n31909);
  not U33640(n31909,n31905);
  nand U33641(n31905,n31910,n31911,n31912,n31913);
  nand U33642(n31913,n27891,n31207);
  nand U33643(n31207,n29541,n28761);
  nand U33644(n31912,G59120,n29229);
  not U33645(n29229,n29261);
  nand U33646(n31911,n29197,n28395);
  nand U33647(n31910,n29230,G59311);
  not U33648(n29230,n29260);
  nand U33649(n31908,n29197,n31914,n31915);
  nand U33650(n31914,n31916,n31917,n31918,n31919);
  nor U33651(n31919,n31920,n31921,n31922,n31923);
  nor U33652(n31923,n29736,n31924);
  nor U33653(n31922,n29737,n31223);
  nor U33654(n31921,n29745,n31221);
  nor U33655(n31920,n29753,n31222);
  nor U33656(n31918,n31925,n31926,n31927,n31928);
  nor U33657(n31928,n29750,n31233);
  nor U33658(n31927,n29761,n31234);
  nor U33659(n31926,n29734,n31235);
  nor U33660(n31925,n29735,n31929);
  nor U33661(n31917,n31930,n31931,n31932,n31933);
  nor U33662(n31933,n29751,n31241);
  nor U33663(n31932,n29742,n31242);
  nor U33664(n31931,n29743,n31243);
  nor U33665(n31930,n29744,n31232);
  nor U33666(n31916,n31934,n31935,n31936,n31937);
  nor U33667(n31937,n29759,n31247);
  nor U33668(n31936,n29760,n31248);
  nor U33669(n31935,n29758,n31249);
  nor U33670(n31934,n29752,n31240);
  nand U33671(n31907,n31938,n29205);
  nand U33672(n31938,n31915,n31939,n31940,n31941);
  nand U33673(n31940,n31324,n31942);
  nand U33674(n31942,n31943,n31944,n31945,n31946);
  nor U33675(n31946,n31947,n31948,n31949,n31950);
  nor U33676(n31950,n29759,n31433);
  nor U33677(n31949,n29758,n31434);
  nor U33678(n31948,n29753,n31435);
  nor U33679(n31947,n29751,n31436);
  nor U33680(n31945,n31951,n31952,n31953,n31954);
  nor U33681(n31954,n29750,n31441);
  nor U33682(n31953,n29745,n31442);
  nor U33683(n31952,n29743,n31443);
  nor U33684(n31951,n29742,n31444);
  nor U33685(n31944,n31955,n31956,n31957,n31958);
  nor U33686(n31958,n29737,n31449);
  nor U33687(n31957,n29735,n31450);
  nor U33688(n31956,n29734,n31451);
  nor U33689(n31955,n29761,n31452);
  nor U33690(n31943,n31959,n31960,n31961,n31962);
  nor U33691(n31962,n29760,n31457);
  nor U33692(n31961,n29752,n31458);
  nor U33693(n31960,n29744,n31459);
  nor U33694(n31959,n29736,n31460);
  nand U33695(n31939,n31250,n30360);
  nand U33696(n30360,n31963,n31964,n31965,n31966);
  nor U33697(n31966,n31967,n31968,n31969,n31970);
  nor U33698(n31970,n29760,n31259);
  nor U33699(n31969,n29759,n31260);
  nor U33700(n31968,n29758,n31261);
  nor U33701(n31967,n29752,n31262);
  nor U33702(n31965,n31971,n31972,n31973,n31974);
  nor U33703(n31974,n29751,n31267);
  nor U33704(n31973,n29750,n31268);
  nor U33705(n31972,n29744,n31269);
  nor U33706(n31971,n29743,n31270);
  nor U33707(n31964,n31975,n31976,n31977,n31978);
  nor U33708(n31978,n29742,n31275);
  nor U33709(n31977,n29736,n31276);
  nor U33710(n31976,n29735,n31277);
  nor U33711(n31975,n29734,n31278);
  nor U33712(n31963,n31979,n31980,n31981,n31982);
  nor U33713(n31982,n29761,n31283);
  nor U33714(n31981,n29753,n31284);
  nor U33715(n31980,n29745,n31285);
  nor U33716(n31979,n29737,n31286);
  and U33717(n31915,n31983,n31984);
  nand U33718(n31984,n29264,n31985);
  nand U33719(n31985,n31986,n31987,n31988,n31989);
  nor U33720(n31989,n31990,n31991,n31992,n31993);
  nor U33721(n31993,n29761,n31296);
  nor U33722(n31992,n29760,n31297);
  nor U33723(n31991,n29759,n31298);
  nor U33724(n31990,n29758,n31299);
  nor U33725(n31988,n31994,n31995,n31996,n31997);
  nor U33726(n31997,n29753,n31304);
  nor U33727(n31996,n29752,n31305);
  nor U33728(n31995,n29751,n31306);
  nor U33729(n31994,n29750,n31307);
  nor U33730(n31987,n31998,n31999,n32000,n32001);
  nor U33731(n32001,n29745,n31312);
  nor U33732(n32000,n29744,n31313);
  nor U33733(n31999,n29743,n31314);
  nor U33734(n31998,n29742,n31315);
  nor U33735(n31986,n32002,n32003,n32004,n32005);
  nor U33736(n32005,n29737,n31320);
  nor U33737(n32004,n29736,n31321);
  nor U33738(n32003,n29735,n31322);
  nor U33739(n32002,n29734,n31323);
  nand U33740(n31983,G59110,n32006);
  nand U33741(n31893,n32007,n32008);
  nand U33742(n32008,n32009,n32010);
  nand U33743(n31895,n29193,n28395);
  nand U33744(G2514,n32011,n32012,n32013,n32014);
  nor U33745(n32014,n32015,n32016,n32017);
  nor U33746(n32017,G59119,n32018,n29185);
  nor U33747(n32016,n32019,n32020);
  nor U33748(n32019,n32021,n29190);
  nor U33749(n32015,n28015,n29192);
  nand U33750(n32012,n29194,n28407);
  xor U33751(n28407,n32010,n32022);
  and U33752(n32022,n32009,n32007);
  or U33753(n32007,n32023,n32024);
  nand U33754(n32009,n32024,n32023);
  xor U33755(n32023,n32025,n29205);
  nand U33756(n32025,n32026,n32027,n32028,n32029);
  nor U33757(n32029,n32030,n32031,n32032,n32033);
  nor U33758(n32033,n32034,n28761);
  nor U33759(n32034,n32035,n32036,n32037,n32038);
  nand U33760(n32038,n32039,n32040,n32041,n32042);
  nand U33761(n32042,n31801,G58986);
  nand U33762(n32041,n31802,G58994);
  nand U33763(n32040,n31803,G59002);
  nand U33764(n32039,n31804,G59010);
  nand U33765(n32037,n32043,n32044,n32045,n32046);
  nand U33766(n32046,n31809,G59018);
  nand U33767(n32045,n31810,G59026);
  nand U33768(n32044,n31811,G59034);
  nand U33769(n32043,n31812,G59042);
  nand U33770(n32036,n32047,n32048,n32049,n32050);
  nand U33771(n32050,n31817,G59050);
  nand U33772(n32049,n31818,G59058);
  nand U33773(n32048,n31819,G59066);
  nand U33774(n32047,n31820,G59074);
  nand U33775(n32035,n32051,n32052,n32053,n32054);
  nand U33776(n32054,n31825,G59082);
  nand U33777(n32053,n31826,G59090);
  nand U33778(n32052,n31827,G59098);
  nand U33779(n32051,n31828,G59106);
  nor U33780(n32032,n32055,n32056,n32057,n32058);
  nand U33781(n32058,n29197,n32059,n32060,n32061);
  nand U33782(n32061,n32062,G59074);
  nand U33783(n32060,n32063,G59042);
  nand U33784(n32059,n32064,G59010);
  nand U33785(n32057,n32065,n32066,n32067,n32068);
  nand U33786(n32068,n31226,G59002);
  nand U33787(n32067,n31227,G58994);
  nand U33788(n32066,n32069,G58986);
  nand U33789(n32065,n32070,G59106);
  nand U33790(n32056,n32071,n32072,n32073,n32074);
  nand U33791(n32074,n32075,G59050);
  nand U33792(n32073,n32076,G59034);
  nand U33793(n32072,n32077,G59026);
  nand U33794(n32071,n32078,G59018);
  nand U33795(n32055,n32079,n32080,n32081,n32082);
  nor U33796(n32082,n32083,n32084);
  nor U33797(n32084,n29855,n31247);
  nor U33798(n32083,n29856,n31248);
  nand U33799(n32081,n32085,G59082);
  nand U33800(n32080,n32086,G59058);
  nand U33801(n32079,n32087,G59066);
  nand U33802(n32028,G59111,n32006);
  nand U33803(n32027,n31324,n32088);
  nand U33804(n32088,n32089,n32090,n32091,n32092);
  nor U33805(n32092,n32093,n32094,n32095,n32096);
  nor U33806(n32096,n29855,n31433);
  nor U33807(n32095,n29854,n31434);
  nor U33808(n32094,n29849,n31435);
  nor U33809(n32093,n29847,n31436);
  nor U33810(n32091,n32097,n32098,n32099,n32100);
  nor U33811(n32100,n29846,n31441);
  nor U33812(n32099,n29841,n31442);
  nor U33813(n32098,n29839,n31443);
  nor U33814(n32097,n29838,n31444);
  nor U33815(n32090,n32101,n32102,n32103,n32104);
  nor U33816(n32104,n29833,n31449);
  nor U33817(n32103,n29831,n31450);
  nor U33818(n32102,n29830,n31451);
  nor U33819(n32101,n29857,n31452);
  nor U33820(n32089,n32105,n32106,n32107,n32108);
  nor U33821(n32108,n29856,n31457);
  nor U33822(n32107,n29848,n31458);
  nor U33823(n32106,n29840,n31459);
  nor U33824(n32105,n29832,n31460);
  nand U33825(n32026,n31250,n30434);
  nand U33826(n30434,n32109,n32110,n32111,n32112);
  nor U33827(n32112,n32113,n32114,n32115,n32116);
  nor U33828(n32116,n29856,n31259);
  nor U33829(n32115,n29855,n31260);
  nor U33830(n32114,n29854,n31261);
  nor U33831(n32113,n29848,n31262);
  nor U33832(n32111,n32117,n32118,n32119,n32120);
  nor U33833(n32120,n29847,n31267);
  nor U33834(n32119,n29846,n31268);
  nor U33835(n32118,n29840,n31269);
  nor U33836(n32117,n29839,n31270);
  nor U33837(n32110,n32121,n32122,n32123,n32124);
  nor U33838(n32124,n29838,n31275);
  nor U33839(n32123,n29832,n31276);
  nor U33840(n32122,n29831,n31277);
  nor U33841(n32121,n29830,n31278);
  nor U33842(n32109,n32125,n32126,n32127,n32128);
  nor U33843(n32128,n29857,n31283);
  nor U33844(n32127,n29849,n31284);
  nor U33845(n32126,n29841,n31285);
  nor U33846(n32125,n29833,n31286);
  and U33847(n32024,n32129,n32130,n32131,n32132);
  nand U33848(n32132,n27900,n29264);
  nor U33849(n32131,n32133,n32134);
  nor U33850(n32134,n28015,n29260);
  nor U33851(n32133,n29261,n32020);
  nand U33852(n32130,n29197,n28406);
  nand U33853(n32129,n27900,n29214);
  nand U33854(n32010,n32135,n32136);
  nand U33855(n32136,n29197,n32137);
  nand U33856(n32137,n32138,n32139);
  not U33857(n32138,n32140);
  nand U33858(n32011,n29193,n28406);
  nand U33859(G2513,n32141,n32142,n32143,n32144);
  nor U33860(n32144,n32145,n32021,n32146);
  nor U33861(n32146,n32018,n29247);
  nor U33862(n32021,G59118,n29185);
  nand U33863(n29185,n32147,n32148);
  nor U33864(n32145,n28013,n29192);
  nand U33865(n32143,n29194,n28431);
  xnor U33866(n28431,n29205,n32149);
  nor U33867(n32149,n32150,n32151);
  not U33868(n32151,n32135);
  nand U33869(n32135,n32152,n32140);
  nor U33870(n32150,n32152,n32140);
  nand U33871(n32140,n32153,n32154,n28691,n32155);
  nor U33872(n32155,n32156,n32157,n32158);
  nor U33873(n32158,n28013,n29260);
  nand U33874(n29260,n32159,n28689,n32160);
  nor U33875(n32157,n28417,n28761);
  nor U33876(n32156,n29261,n32018);
  nand U33877(n32154,n29197,n27969);
  nand U33878(n32153,n27915,n29214);
  not U33879(n29214,n29541);
  nor U33880(n29541,n31324,n31250);
  xnor U33881(n32152,n32139,n29205);
  nand U33882(n32139,n32163,n32164,n32165,n32166);
  nor U33883(n32166,n32161,n32162,n32167,n32168);
  nor U33884(n32168,n32169,n28761);
  nor U33885(n32169,n32170,n32171,n32172,n32173);
  nand U33886(n32173,n32174,n32175,n32176,n32177);
  nand U33887(n32177,n31801,G58987);
  not U33888(n31801,n31323);
  nand U33889(n31323,n32178,n32179);
  nand U33890(n32176,n31802,G58995);
  not U33891(n31802,n31322);
  nand U33892(n31322,n32178,n32180);
  nand U33893(n32175,n31803,G59003);
  not U33894(n31803,n31321);
  nand U33895(n31321,n32181,n32179);
  nand U33896(n32174,n31804,G59011);
  not U33897(n31804,n31320);
  nand U33898(n31320,n32181,n32180);
  nand U33899(n32172,n32182,n32183,n32184,n32185);
  nand U33900(n32185,n31809,G59019);
  not U33901(n31809,n31315);
  nand U33902(n31315,n32178,n32186);
  nand U33903(n32184,n31810,G59027);
  not U33904(n31810,n31314);
  nand U33905(n31314,n32178,n32187);
  nor U33906(n32178,n32188,n32189);
  nand U33907(n32183,n31811,G59035);
  not U33908(n31811,n31313);
  nand U33909(n31313,n32181,n32186);
  nand U33910(n32182,n31812,G59043);
  not U33911(n31812,n31312);
  nand U33912(n31312,n32181,n32187);
  nor U33913(n32181,n32190,n32188);
  nand U33914(n32171,n32191,n32192,n32193,n32194);
  nand U33915(n32194,n31817,G59051);
  not U33916(n31817,n31307);
  nand U33917(n31307,n32179,n32195);
  nand U33918(n32193,n31818,G59059);
  not U33919(n31818,n31306);
  nand U33920(n31306,n32180,n32195);
  nand U33921(n32192,n31819,G59067);
  not U33922(n31819,n31305);
  nand U33923(n31305,n32179,n32196);
  nor U33924(n32179,n32197,G59112);
  nand U33925(n32191,n31820,G59075);
  not U33926(n31820,n31304);
  nand U33927(n31304,n32180,n32196);
  nor U33928(n32180,n32197,n29944);
  nand U33929(n32170,n32198,n32199,n32200,n32201);
  nand U33930(n32201,n31825,G59083);
  not U33931(n31825,n31299);
  nand U33932(n31299,n32186,n32195);
  nand U33933(n32200,n31826,G59091);
  not U33934(n31826,n31298);
  nand U33935(n31298,n32187,n32195);
  and U33936(n32195,n32190,n32188);
  not U33937(n32190,n32189);
  nand U33938(n32199,n31827,G59099);
  not U33939(n31827,n31297);
  nand U33940(n31297,n32196,n32186);
  and U33941(n32186,n32197,n29944);
  nand U33942(n32198,n31828,G59107);
  not U33943(n31828,n31296);
  nand U33944(n31296,n32196,n32187);
  and U33945(n32187,G59112,n32197);
  and U33946(n32196,n32189,n32188);
  nor U33947(n32167,n32202,n32203,n32204,n32205);
  nand U33948(n32205,n29197,n32206,n32207,n32208);
  nand U33949(n32208,n32062,G59075);
  not U33950(n32062,n31222);
  nand U33951(n31222,n32209,n32210);
  nand U33952(n32207,n32063,G59043);
  not U33953(n32063,n31221);
  nand U33954(n31221,n32211,n32212);
  nand U33955(n32206,n32064,G59011);
  not U33956(n32064,n31223);
  nand U33957(n31223,n32212,n32210);
  nand U33958(n32204,n32213,n32214,n32215,n32216);
  nand U33959(n32216,n31226,G59003);
  not U33960(n31226,n31924);
  nand U33961(n31924,n32217,n32212);
  nand U33962(n32215,n31227,G58995);
  not U33963(n31227,n31929);
  nand U33964(n31929,n32218,n32210);
  nand U33965(n32214,n32069,G58987);
  not U33966(n32069,n31235);
  nand U33967(n31235,n32218,n32217);
  nand U33968(n32213,n32070,G59107);
  not U33969(n32070,n31234);
  nand U33970(n31234,n32211,n32209);
  nand U33971(n32203,n32219,n32220,n32221,n32222);
  nand U33972(n32222,n32075,G59051);
  not U33973(n32075,n31233);
  nand U33974(n31233,n32223,n32217);
  nand U33975(n32221,n32076,G59035);
  not U33976(n32076,n31232);
  nand U33977(n31232,n32224,n32212);
  nor U33978(n32212,n28381,n27900);
  nand U33979(n32220,n32077,G59027);
  not U33980(n32077,n31243);
  nand U33981(n31243,n32218,n32211);
  nand U33982(n32219,n32078,G59019);
  not U33983(n32078,n31242);
  nand U33984(n31242,n32224,n32218);
  nor U33985(n32218,n28405,n28381);
  not U33986(n28381,n27881);
  nand U33987(n32202,n32225,n32226,n32227,n32228);
  nor U33988(n32228,n32229,n32230);
  nor U33989(n32230,n29946,n31247);
  nand U33990(n31247,n32223,n32211);
  nor U33991(n32211,n27915,n27891);
  nor U33992(n32229,n29947,n31248);
  nand U33993(n31248,n32224,n32209);
  nand U33994(n32227,n32085,G59083);
  not U33995(n32085,n31249);
  nand U33996(n31249,n32224,n32223);
  nor U33997(n32224,n28417,n27891);
  nand U33998(n32226,n32086,G59059);
  not U33999(n32086,n31241);
  nand U34000(n31241,n32223,n32210);
  nor U34001(n32210,n27915,n28393);
  nor U34002(n32223,n28405,n27881);
  nand U34003(n32225,n32087,G59067);
  not U34004(n32087,n31240);
  nand U34005(n31240,n32217,n32209);
  nor U34006(n32209,n27900,n27881);
  nor U34007(n32217,n28393,n28417);
  not U34008(n28417,n27915);
  nand U34009(n32165,G59112,n32006);
  nand U34010(n32164,n31324,n32231);
  nand U34011(n32231,n32232,n32233,n32234,n32235);
  nor U34012(n32235,n32236,n32237,n32238,n32239);
  nor U34013(n32239,n29946,n31433);
  nor U34014(n32238,n29942,n31434);
  nor U34015(n32237,n29937,n31435);
  nor U34016(n32236,n29935,n31436);
  nor U34017(n32234,n32240,n32241,n32242,n32243);
  nor U34018(n32243,n29933,n31441);
  nor U34019(n32242,n29927,n31442);
  nor U34020(n32241,n29925,n31443);
  nor U34021(n32240,n29923,n31444);
  nor U34022(n32233,n32244,n32245,n32246,n32247);
  nor U34023(n32247,n29915,n31449);
  nor U34024(n32246,n29911,n31450);
  nor U34025(n32245,n29908,n31451);
  nor U34026(n32244,n29949,n31452);
  nor U34027(n32232,n32248,n32249,n32250,n32251);
  nor U34028(n32251,n29947,n31457);
  nor U34029(n32250,n29936,n31458);
  nor U34030(n32249,n29926,n31459);
  nor U34031(n32248,n29913,n31460);
  nand U34032(n32163,n31250,n30514);
  nand U34033(n30514,n32252,n32253,n32254,n32255);
  nor U34034(n32255,n32256,n32257,n32258,n32259);
  nor U34035(n32259,n29947,n31259);
  nand U34036(n31259,n32260,n32261);
  nor U34037(n32258,n29946,n31260);
  nand U34038(n31260,n32262,n32260);
  nor U34039(n32257,n29942,n31261);
  nand U34040(n31261,n32260,n32263);
  nor U34041(n32256,n29936,n31262);
  nand U34042(n31262,n32264,n32261);
  nor U34043(n32254,n32265,n32266,n32267,n32268);
  nor U34044(n32268,n29935,n31267);
  nand U34045(n31267,n32262,n32264);
  nor U34046(n32267,n29933,n31268);
  nand U34047(n31268,n32263,n32264);
  nor U34048(n32266,n29926,n31269);
  nand U34049(n31269,n32269,n32261);
  nor U34050(n32265,n29925,n31270);
  nand U34051(n31270,n32269,n32262);
  nor U34052(n32253,n32270,n32271,n32272,n32273);
  nor U34053(n32273,n29923,n31275);
  nand U34054(n31275,n32269,n32263);
  nor U34055(n32272,n29913,n31276);
  nand U34056(n31276,n32274,n32261);
  nor U34057(n32261,n32275,n28406);
  nor U34058(n32271,n29911,n31277);
  nand U34059(n31277,n32274,n32262);
  nor U34060(n32262,n27969,n29166);
  nor U34061(n32270,n29908,n31278);
  nand U34062(n31278,n32274,n32263);
  nor U34063(n32263,n29166,n32275);
  nor U34064(n32252,n32276,n32277,n32278,n32279);
  nor U34065(n32279,n29949,n31283);
  nand U34066(n31283,n32280,n32260);
  nor U34067(n32260,n28395,n28383);
  nor U34068(n32278,n29937,n31284);
  nand U34069(n31284,n32280,n32264);
  nor U34070(n32264,n29159,n28383);
  nor U34071(n32277,n29927,n31285);
  nand U34072(n31285,n32280,n32269);
  nor U34073(n32269,n29152,n28395);
  nor U34074(n32276,n29915,n31286);
  nand U34075(n31286,n32280,n32274);
  nor U34076(n32274,n29159,n29152);
  nor U34077(n32280,n27969,n28406);
  nor U34078(n31250,n27916,n28959,n32281);
  nand U34079(n32282,n32283,n32284,n32285,n32286);
  nand U34080(n32142,n29193,n27969);
  not U34081(n29193,n29685);
  nand U34082(n29685,n32147,n32287);
  nand U34083(n32287,n32288,n32289,n32290,n32291);
  nand U34084(n32141,n29231,n27915);
  not U34085(n29231,n30662);
  nand U34086(n30662,n32147,n32292);
  nand U34087(n32292,n32293,n32294,n32295,n32296);
  nor U34088(n32296,n32297,n32298);
  not U34089(n32294,n32299);
  nor U34090(n32147,n27929,n29190);
  not U34091(n29190,n29247);
  nand U34092(n29247,n28438,n32300);
  nand U34093(n32300,n27907,n32301);
  nand U34094(n32301,n32302,n32303,n32304,n32305);
  nand U34095(n32305,n28691,n28419,n32306);
  nand U34096(n32304,n32307,n27930);
  nand U34097(n32307,n32308,n32309);
  nand U34098(n32309,n32306,n32310,n32311);
  nand U34099(n32308,n32312,n27965);
  nand U34100(n32312,n32313,n32314);
  nand U34101(n32314,n32315,n32006);
  nand U34102(n32315,n27942,n27944);
  nand U34103(n32313,n32160,n27945);
  nand U34104(n32303,n27965,n32316);
  nand U34105(n28438,n27928,n28416,n27960);
  nand U34106(G2512,n32317,n32318,n32319);
  nand U34107(n32319,n27967,G59116);
  nand U34108(n32318,n27968,n28406);
  nand U34109(n32317,n27970,n27899);
  nand U34110(G2511,n32320,n32321,n32322);
  nand U34111(n32322,n27967,G59115);
  nand U34112(n32321,n27968,n28395);
  nand U34113(n32320,n27970,n27890);
  nand U34114(G2510,n32323,n32324,n32325);
  nand U34115(n32325,n27967,G59114);
  nand U34116(n32324,n27968,n28383);
  and U34117(n27968,n32326,n27966);
  nand U34118(n32326,n32327,n32328);
  nand U34119(n32328,n29174,n27929);
  nand U34120(n32323,n27970,n32329);
  nor U34121(n27970,n27967,G58977,n29174);
  not U34122(n27967,n27966);
  nor U34123(G2509,n32330,n27966);
  nand U34124(n27966,n32331,n27905,n32332);
  nand U34125(n27905,G59346,n32333);
  nand U34126(n32331,n27916,n32333);
  nand U34127(G2508,n32334,n32335,n32336,n32337);
  nor U34128(n32337,n32338,n32339,n32340);
  nor U34129(n32340,n26769,n32341);
  nor U34130(n32339,n32342,n32343);
  nor U34131(n32338,n29968,n32344);
  nand U34132(n32336,n32345,G59107);
  nand U34133(n32335,n32346,n32347);
  nand U34134(n32334,G58871,n32348);
  nand U34135(G2507,n32349,n32350,n32351,n32352);
  nor U34136(n32352,n32353,n32354,n32355);
  nor U34137(n32355,n26792,n32341);
  nor U34138(n32354,n32356,n32343);
  nor U34139(n32353,n29968,n32357);
  nand U34140(n32351,n32345,G59106);
  nand U34141(n32350,n32358,n32347);
  nand U34142(n32349,G58872,n32348);
  nand U34143(G2506,n32359,n32360,n32361,n32362);
  nor U34144(n32362,n32363,n32364,n32365);
  nor U34145(n32365,n26809,n32341);
  nor U34146(n32364,n32366,n32343);
  nor U34147(n32363,n29968,n32367);
  nand U34148(n32361,n32345,G59105);
  nand U34149(n32360,n32368,n32347);
  nand U34150(n32359,G58873,n32348);
  nand U34151(G2505,n32369,n32370,n32371,n32372);
  nor U34152(n32372,n32373,n32374,n32375);
  nor U34153(n32375,n26826,n32341);
  nor U34154(n32374,n32376,n32343);
  nor U34155(n32373,n29968,n32377);
  nand U34156(n32371,n32345,G59104);
  nand U34157(n32370,n32378,n32347);
  nand U34158(n32369,G58874,n32348);
  nand U34159(G2504,n32379,n32380,n32381,n32382);
  nor U34160(n32382,n32383,n32384,n32385);
  nor U34161(n32385,n26843,n32341);
  nor U34162(n32384,n32386,n32343);
  nor U34163(n32383,n29968,n32387);
  nand U34164(n32381,n32345,G59103);
  nand U34165(n32380,n32388,n32347);
  nand U34166(n32379,G58875,n32348);
  nand U34167(G2503,n32389,n32390,n32391,n32392);
  nor U34168(n32392,n32393,n32394,n32395);
  nor U34169(n32395,n26860,n32341);
  nor U34170(n32394,n32396,n32343);
  nor U34171(n32393,n29968,n32397);
  nand U34172(n32391,n32345,G59102);
  nand U34173(n32390,n32398,n32347);
  nand U34174(n32389,G58876,n32348);
  nand U34175(G2502,n32399,n32400,n32401,n32402);
  nor U34176(n32402,n32403,n32404,n32405);
  nor U34177(n32405,n26878,n32341);
  nor U34178(n32404,n32406,n32343);
  nor U34179(n32403,n29968,n32407);
  nand U34180(n32401,n32345,G59101);
  nand U34181(n32400,n32408,n32347);
  nand U34182(n32399,G58877,n32348);
  nand U34183(G2501,n32409,n32410,n32411,n32412);
  nor U34184(n32412,n32413,n32414,n32415);
  nor U34185(n32415,n26905,n32341);
  nand U34186(n32341,n32416,n29968,n32417);
  nor U34187(n32414,n32418,n32343);
  nor U34188(n32413,n29968,n32419);
  nand U34189(n32411,n32345,G59100);
  and U34190(n32345,n32420,n32421);
  nand U34191(n32421,n32422,n32423,n32424);
  nand U34192(n32424,G58977,n31452);
  nand U34193(n32422,n32425,n32426);
  nand U34194(n32420,n32427,n32428);
  nand U34195(n32410,n32429,n32347);
  nand U34196(n32347,n32430,n32431);
  or U34197(n32431,n32426,n29174);
  nand U34198(n32430,n32416,G58977);
  not U34199(n32416,n31452);
  nand U34200(n32409,G58878,n32348);
  nand U34201(n32348,n32432,n32433);
  nand U34202(n32433,n32427,n32425);
  nand U34203(n32425,n32434,n32435);
  not U34204(n32427,n32343);
  nand U34205(n32343,n32436,n32437);
  or U34206(n32432,n32435,n32426);
  nand U34207(n32426,n32438,n32439);
  nand U34208(n32435,n29968,n31452,n32417);
  nand U34209(n29968,n32440,n32441);
  nand U34210(G2500,n32442,n32443,n32444,n32445);
  nor U34211(n32445,n32446,n32447,n32448);
  nor U34212(n32448,n32449,n26779);
  nor U34213(n32447,n32450,n32451);
  nor U34214(n32446,n29947,n32452);
  nand U34215(n32444,n32453,G58887);
  nand U34216(n32443,n32454,n32455);
  nand U34217(n32442,n32456,n32457);
  nand U34218(G2499,n32458,n32459,n32460,n32461);
  nor U34219(n32461,n32462,n32463,n32464);
  nor U34220(n32464,n32449,n26797);
  nor U34221(n32463,n32450,n32465);
  nor U34222(n32462,n29856,n32452);
  nand U34223(n32460,n32453,G58888);
  nand U34224(n32459,n32466,n32455);
  nand U34225(n32458,n32456,n32467);
  nand U34226(G2498,n32468,n32469,n32470,n32471);
  nor U34227(n32471,n32472,n32473,n32474);
  nor U34228(n32474,n32449,n26814);
  nor U34229(n32473,n32450,n32475);
  nor U34230(n32472,n29760,n32452);
  nand U34231(n32470,n32453,G58889);
  nand U34232(n32469,n32476,n32455);
  nand U34233(n32468,n32456,n32477);
  nand U34234(G2497,n32478,n32479,n32480,n32481);
  nor U34235(n32481,n32482,n32483,n32484);
  nor U34236(n32484,n32449,n26831);
  nor U34237(n32483,n32450,n32485);
  nor U34238(n32482,n30304,n32452);
  nand U34239(n32480,n32453,G58890);
  nand U34240(n32479,n32486,n32455);
  nand U34241(n32478,n32456,n32487);
  nand U34242(G2496,n32488,n32489,n32490,n32491);
  nor U34243(n32491,n32492,n32493,n32494);
  nor U34244(n32494,n32449,n26848);
  nor U34245(n32493,n32450,n32495);
  nor U34246(n32492,n30220,n32452);
  nand U34247(n32490,n32453,G58891);
  nand U34248(n32489,n32496,n32455);
  nand U34249(n32488,n32456,n32497);
  nand U34250(G2495,n32498,n32499,n32500,n32501);
  nor U34251(n32501,n32502,n32503,n32504);
  nor U34252(n32504,n32449,n26866);
  nor U34253(n32503,n32450,n32505);
  nor U34254(n32502,n30139,n32452);
  nand U34255(n32500,n32453,G58892);
  nand U34256(n32499,n32506,n32455);
  nand U34257(n32498,n32456,n32507);
  nand U34258(G2494,n32508,n32509,n32510,n32511);
  nor U34259(n32511,n32512,n32513,n32514);
  nor U34260(n32514,n32449,n26883);
  nor U34261(n32513,n32450,n32515);
  nor U34262(n32512,n29438,n32452);
  nand U34263(n32510,n32453,G58893);
  nand U34264(n32509,n32516,n32455);
  nand U34265(n32508,n32456,n32517);
  nand U34266(G2493,n32518,n32519,n32520,n32521);
  nor U34267(n32521,n32522,n32523,n32524);
  nor U34268(n32524,n32449,n26913);
  and U34269(n32449,n32525,n32526);
  nand U34270(n32526,n32527,n29966,n32417);
  nand U34271(n32527,n32528,n32529);
  nand U34272(n32525,n32456,n32530);
  nor U34273(n32523,n32450,n32531);
  and U34274(n32450,n32532,n32533);
  or U34275(n32533,n32529,n29174);
  nand U34276(n32532,n32534,G58977);
  nor U34277(n32522,n29965,n32452);
  nand U34278(n32452,n32535,n32536);
  nand U34279(n32536,n32537,n32423,n32538);
  nand U34280(n32538,n32530,n32529);
  nand U34281(n32537,n32539,n31457);
  nand U34282(n32539,n32540,n27929);
  nand U34283(n32540,n32529,n29966);
  nand U34284(n32529,n32541,n32439);
  nand U34285(n32535,n32456,n32428);
  nand U34286(n32520,n32453,G58894);
  and U34287(n32453,n32417,n32534);
  not U34288(n32534,n31457);
  nand U34289(n32519,n32542,n32455);
  not U34290(n32455,n29966);
  nand U34291(n29966,n32543,n32441);
  nand U34292(n32518,n32456,n32544);
  not U34293(n32456,n32528);
  nand U34294(n32528,n32545,n32437);
  nand U34295(G2492,n32546,n32547,n32548,n32549);
  nor U34296(n32549,n32550,n32551,n32552);
  nor U34297(n32552,n26769,n32553);
  nor U34298(n32551,n32342,n32554);
  nor U34299(n32550,n29964,n32344);
  nand U34300(n32548,n32555,G59091);
  nand U34301(n32547,n32346,n32556);
  nand U34302(n32546,G58871,n32557);
  nand U34303(G2491,n32558,n32559,n32560,n32561);
  nor U34304(n32561,n32562,n32563,n32564);
  nor U34305(n32564,n26792,n32553);
  nor U34306(n32563,n32356,n32554);
  nor U34307(n32562,n29964,n32357);
  nand U34308(n32560,n32555,G59090);
  nand U34309(n32559,n32358,n32556);
  nand U34310(n32558,G58872,n32557);
  nand U34311(G2490,n32565,n32566,n32567,n32568);
  nor U34312(n32568,n32569,n32570,n32571);
  nor U34313(n32571,n26809,n32553);
  nor U34314(n32570,n32366,n32554);
  nor U34315(n32569,n29964,n32367);
  nand U34316(n32567,n32555,G59089);
  nand U34317(n32566,n32368,n32556);
  nand U34318(n32565,G58873,n32557);
  nand U34319(G2489,n32572,n32573,n32574,n32575);
  nor U34320(n32575,n32576,n32577,n32578);
  nor U34321(n32578,n26826,n32553);
  nor U34322(n32577,n32376,n32554);
  nor U34323(n32576,n29964,n32377);
  nand U34324(n32574,n32555,G59088);
  nand U34325(n32573,n32378,n32556);
  nand U34326(n32572,G58874,n32557);
  nand U34327(G2488,n32579,n32580,n32581,n32582);
  nor U34328(n32582,n32583,n32584,n32585);
  nor U34329(n32585,n26843,n32553);
  nor U34330(n32584,n32386,n32554);
  nor U34331(n32583,n29964,n32387);
  nand U34332(n32581,n32555,G59087);
  nand U34333(n32580,n32388,n32556);
  nand U34334(n32579,G58875,n32557);
  nand U34335(G2487,n32586,n32587,n32588,n32589);
  nor U34336(n32589,n32590,n32591,n32592);
  nor U34337(n32592,n26860,n32553);
  nor U34338(n32591,n32396,n32554);
  nor U34339(n32590,n29964,n32397);
  nand U34340(n32588,n32555,G59086);
  nand U34341(n32587,n32398,n32556);
  nand U34342(n32586,G58876,n32557);
  nand U34343(G2486,n32593,n32594,n32595,n32596);
  nor U34344(n32596,n32597,n32598,n32599);
  nor U34345(n32599,n26878,n32553);
  nor U34346(n32598,n32406,n32554);
  nor U34347(n32597,n29964,n32407);
  nand U34348(n32595,n32555,G59085);
  nand U34349(n32594,n32408,n32556);
  nand U34350(n32593,G58877,n32557);
  nand U34351(G2485,n32600,n32601,n32602,n32603);
  nor U34352(n32603,n32604,n32605,n32606);
  nor U34353(n32606,n26905,n32553);
  nand U34354(n32553,n32607,n29964,n32417);
  nor U34355(n32605,n32418,n32554);
  nor U34356(n32604,n29964,n32419);
  nand U34357(n32602,n32555,G59084);
  and U34358(n32555,n32608,n32609);
  nand U34359(n32609,n32610,n32423,n32611);
  nand U34360(n32611,G58977,n31433);
  nand U34361(n32610,n32612,n32613);
  nand U34362(n32608,n32614,n32428);
  nand U34363(n32601,n32429,n32556);
  nand U34364(n32556,n32615,n32616);
  or U34365(n32616,n32613,n29174);
  nand U34366(n32615,n32607,G58977);
  not U34367(n32607,n31433);
  nand U34368(n32600,G58878,n32557);
  nand U34369(n32557,n32617,n32618);
  nand U34370(n32618,n32614,n32612);
  nand U34371(n32612,n32434,n32619);
  not U34372(n32614,n32554);
  nand U34373(n32554,n32620,n32437);
  or U34374(n32617,n32619,n32613);
  nand U34375(n32613,n32621,n32439);
  nand U34376(n32619,n29964,n31433,n32417);
  nand U34377(n29964,n32622,n32440);
  nand U34378(G2484,n32623,n32624,n32625,n32626);
  nor U34379(n32626,n32627,n32628,n32629);
  nor U34380(n32629,n32342,n32630);
  nor U34381(n32628,n29962,n32344);
  nor U34382(n32627,n26769,n32631);
  nand U34383(n32625,n32632,G59083);
  nand U34384(n32624,n32346,n32633);
  nand U34385(n32623,G58871,n32634);
  nand U34386(G2483,n32635,n32636,n32637,n32638);
  nor U34387(n32638,n32639,n32640,n32641);
  nor U34388(n32641,n32356,n32630);
  nor U34389(n32640,n29962,n32357);
  nor U34390(n32639,n26792,n32631);
  nand U34391(n32637,n32632,G59082);
  nand U34392(n32636,n32358,n32633);
  nand U34393(n32635,G58872,n32634);
  nand U34394(G2482,n32642,n32643,n32644,n32645);
  nor U34395(n32645,n32646,n32647,n32648);
  nor U34396(n32648,n32366,n32630);
  nor U34397(n32647,n29962,n32367);
  nor U34398(n32646,n26809,n32631);
  nand U34399(n32644,n32632,G59081);
  nand U34400(n32643,n32368,n32633);
  nand U34401(n32642,G58873,n32634);
  nand U34402(G2481,n32649,n32650,n32651,n32652);
  nor U34403(n32652,n32653,n32654,n32655);
  nor U34404(n32655,n32376,n32630);
  nor U34405(n32654,n29962,n32377);
  nor U34406(n32653,n26826,n32631);
  nand U34407(n32651,n32632,G59080);
  nand U34408(n32650,n32378,n32633);
  nand U34409(n32649,G58874,n32634);
  nand U34410(G2480,n32656,n32657,n32658,n32659);
  nor U34411(n32659,n32660,n32661,n32662);
  nor U34412(n32662,n32386,n32630);
  nor U34413(n32661,n29962,n32387);
  nor U34414(n32660,n26843,n32631);
  nand U34415(n32658,n32632,G59079);
  nand U34416(n32657,n32388,n32633);
  nand U34417(n32656,G58875,n32634);
  nand U34418(G2479,n32663,n32664,n32665,n32666);
  nor U34419(n32666,n32667,n32668,n32669);
  nor U34420(n32669,n32396,n32630);
  nor U34421(n32668,n29962,n32397);
  nor U34422(n32667,n26860,n32631);
  nand U34423(n32665,n32632,G59078);
  nand U34424(n32664,n32398,n32633);
  nand U34425(n32663,G58876,n32634);
  nand U34426(G2478,n32670,n32671,n32672,n32673);
  nor U34427(n32673,n32674,n32675,n32676);
  nor U34428(n32676,n32406,n32630);
  nor U34429(n32675,n29962,n32407);
  nor U34430(n32674,n26878,n32631);
  nand U34431(n32672,n32632,G59077);
  nand U34432(n32671,n32408,n32633);
  nand U34433(n32670,G58877,n32634);
  nand U34434(G2477,n32677,n32678,n32679,n32680);
  nor U34435(n32680,n32681,n32682,n32683);
  nor U34436(n32683,n32418,n32630);
  nor U34437(n32682,n29962,n32419);
  nor U34438(n32681,n26905,n32631);
  nand U34439(n32631,n32417,n32684);
  nand U34440(n32679,n32632,G59076);
  and U34441(n32632,n32685,n32686);
  nand U34442(n32686,n32687,n32423,n32688);
  nand U34443(n32688,G58977,n31434);
  nand U34444(n32687,n32689,n32690);
  nand U34445(n32685,n32691,n32428);
  nand U34446(n32678,n32429,n32633);
  nand U34447(n32633,n32692,n32693);
  nand U34448(n32693,n32694,n29226);
  nand U34449(n32692,n32684,G58977);
  not U34450(n32684,n31434);
  nand U34451(n32677,G58878,n32634);
  nand U34452(n32634,n32695,n32696);
  nand U34453(n32696,n32417,n29962,n32694);
  not U34454(n32694,n32690);
  nand U34455(n32690,n32697,n32439);
  nor U34456(n32439,n32698,n32699);
  nand U34457(n32695,n32691,n32689);
  nand U34458(n32689,n32434,n32700);
  nand U34459(n32700,n29962,n31434,n32417);
  nand U34460(n29962,n32622,n32543);
  not U34461(n32691,n32630);
  nand U34462(n32630,n32437,n32701);
  nor U34463(n32437,G59115,G59114);
  nand U34464(G2476,n32702,n32703,n32704,n32705);
  nor U34465(n32705,n32706,n32707,n32708);
  nor U34466(n32708,n26769,n32709);
  nor U34467(n32707,n32342,n32710);
  nor U34468(n32706,n29980,n32344);
  nand U34469(n32704,n32711,G59075);
  nand U34470(n32703,n32346,n32712);
  nand U34471(n32702,G58871,n32713);
  nand U34472(G2475,n32714,n32715,n32716,n32717);
  nor U34473(n32717,n32718,n32719,n32720);
  nor U34474(n32720,n26792,n32709);
  nor U34475(n32719,n32356,n32710);
  nor U34476(n32718,n29980,n32357);
  nand U34477(n32716,n32711,G59074);
  nand U34478(n32715,n32358,n32712);
  nand U34479(n32714,G58872,n32713);
  nand U34480(G2474,n32721,n32722,n32723,n32724);
  nor U34481(n32724,n32725,n32726,n32727);
  nor U34482(n32727,n26809,n32709);
  nor U34483(n32726,n32366,n32710);
  nor U34484(n32725,n29980,n32367);
  nand U34485(n32723,n32711,G59073);
  nand U34486(n32722,n32368,n32712);
  nand U34487(n32721,G58873,n32713);
  nand U34488(G2473,n32728,n32729,n32730,n32731);
  nor U34489(n32731,n32732,n32733,n32734);
  nor U34490(n32734,n26826,n32709);
  nor U34491(n32733,n32376,n32710);
  nor U34492(n32732,n29980,n32377);
  nand U34493(n32730,n32711,G59072);
  nand U34494(n32729,n32378,n32712);
  nand U34495(n32728,G58874,n32713);
  nand U34496(G2472,n32735,n32736,n32737,n32738);
  nor U34497(n32738,n32739,n32740,n32741);
  nor U34498(n32741,n26843,n32709);
  nor U34499(n32740,n32386,n32710);
  nor U34500(n32739,n29980,n32387);
  nand U34501(n32737,n32711,G59071);
  nand U34502(n32736,n32388,n32712);
  nand U34503(n32735,G58875,n32713);
  nand U34504(G2471,n32742,n32743,n32744,n32745);
  nor U34505(n32745,n32746,n32747,n32748);
  nor U34506(n32748,n26860,n32709);
  nor U34507(n32747,n32396,n32710);
  nor U34508(n32746,n29980,n32397);
  nand U34509(n32744,n32711,G59070);
  nand U34510(n32743,n32398,n32712);
  nand U34511(n32742,G58876,n32713);
  nand U34512(G2470,n32749,n32750,n32751,n32752);
  nor U34513(n32752,n32753,n32754,n32755);
  nor U34514(n32755,n26878,n32709);
  nor U34515(n32754,n32406,n32710);
  nor U34516(n32753,n29980,n32407);
  nand U34517(n32751,n32711,G59069);
  nand U34518(n32750,n32408,n32712);
  nand U34519(n32749,G58877,n32713);
  nand U34520(G2469,n32756,n32757,n32758,n32759);
  nor U34521(n32759,n32760,n32761,n32762);
  nor U34522(n32762,n26905,n32709);
  nand U34523(n32709,n32763,n29980,n32417);
  nor U34524(n32761,n32418,n32710);
  nor U34525(n32760,n29980,n32419);
  nand U34526(n32758,n32711,G59068);
  and U34527(n32711,n32764,n32765);
  nand U34528(n32765,n32766,n32423,n32767);
  nand U34529(n32767,G58977,n31435);
  nand U34530(n32766,n32768,n32769);
  nand U34531(n32764,n32770,n32428);
  nand U34532(n32757,n32429,n32712);
  nand U34533(n32712,n32771,n32772);
  or U34534(n32772,n32769,n29174);
  nand U34535(n32771,n32763,G58977);
  not U34536(n32763,n31435);
  nand U34537(n32756,G58878,n32713);
  nand U34538(n32713,n32773,n32774);
  nand U34539(n32774,n32770,n32768);
  nand U34540(n32768,n32434,n32775);
  not U34541(n32770,n32710);
  nand U34542(n32710,n32436,n32776);
  or U34543(n32773,n32775,n32769);
  nand U34544(n32769,n32777,n32438);
  nand U34545(n32775,n29980,n31435,n32417);
  nand U34546(n29980,n32778,n32441);
  nand U34547(G2468,n32779,n32780,n32781,n32782);
  nor U34548(n32782,n32783,n32784,n32785);
  nor U34549(n32785,n32342,n32786);
  nor U34550(n32784,n29978,n32344);
  nor U34551(n32783,n26769,n32787);
  nand U34552(n32781,n32788,G59067);
  nand U34553(n32780,n32346,n32789);
  nand U34554(n32779,G58871,n32790);
  nand U34555(G2467,n32791,n32792,n32793,n32794);
  nor U34556(n32794,n32795,n32796,n32797);
  nor U34557(n32797,n32356,n32786);
  nor U34558(n32796,n29978,n32357);
  nor U34559(n32795,n26792,n32787);
  nand U34560(n32793,n32788,G59066);
  nand U34561(n32792,n32358,n32789);
  nand U34562(n32791,G58872,n32790);
  nand U34563(G2466,n32798,n32799,n32800,n32801);
  nor U34564(n32801,n32802,n32803,n32804);
  nor U34565(n32804,n32366,n32786);
  nor U34566(n32803,n29978,n32367);
  nor U34567(n32802,n26809,n32787);
  nand U34568(n32800,n32788,G59065);
  nand U34569(n32799,n32368,n32789);
  nand U34570(n32798,G58873,n32790);
  nand U34571(G2465,n32805,n32806,n32807,n32808);
  nor U34572(n32808,n32809,n32810,n32811);
  nor U34573(n32811,n32376,n32786);
  nor U34574(n32810,n29978,n32377);
  nor U34575(n32809,n26826,n32787);
  nand U34576(n32807,n32788,G59064);
  nand U34577(n32806,n32378,n32789);
  nand U34578(n32805,G58874,n32790);
  nand U34579(G2464,n32812,n32813,n32814,n32815);
  nor U34580(n32815,n32816,n32817,n32818);
  nor U34581(n32818,n32386,n32786);
  nor U34582(n32817,n29978,n32387);
  nor U34583(n32816,n26843,n32787);
  nand U34584(n32814,n32788,G59063);
  nand U34585(n32813,n32388,n32789);
  nand U34586(n32812,G58875,n32790);
  nand U34587(G2463,n32819,n32820,n32821,n32822);
  nor U34588(n32822,n32823,n32824,n32825);
  nor U34589(n32825,n32396,n32786);
  nor U34590(n32824,n29978,n32397);
  nor U34591(n32823,n26860,n32787);
  nand U34592(n32821,n32788,G59062);
  nand U34593(n32820,n32398,n32789);
  nand U34594(n32819,G58876,n32790);
  nand U34595(G2462,n32826,n32827,n32828,n32829);
  nor U34596(n32829,n32830,n32831,n32832);
  nor U34597(n32832,n32406,n32786);
  nor U34598(n32831,n29978,n32407);
  nor U34599(n32830,n26878,n32787);
  nand U34600(n32828,n32788,G59061);
  nand U34601(n32827,n32408,n32789);
  nand U34602(n32826,G58877,n32790);
  nand U34603(G2461,n32833,n32834,n32835,n32836);
  nor U34604(n32836,n32837,n32838,n32839);
  nor U34605(n32839,n32418,n32786);
  nor U34606(n32838,n29978,n32419);
  nor U34607(n32837,n26905,n32787);
  nand U34608(n32787,n32417,n32840);
  nand U34609(n32835,n32788,G59060);
  and U34610(n32788,n32841,n32842);
  nand U34611(n32842,n32843,n32423,n32844);
  nand U34612(n32844,G58977,n31458);
  nand U34613(n32843,n32845,n32846);
  nand U34614(n32841,n32847,n32428);
  nand U34615(n32834,n32429,n32789);
  nand U34616(n32789,n32848,n32849);
  nand U34617(n32849,n32850,n29226);
  nand U34618(n32848,n32840,G58977);
  not U34619(n32840,n31458);
  nand U34620(n32833,G58878,n32790);
  nand U34621(n32790,n32851,n32852);
  nand U34622(n32852,n32417,n29978,n32850);
  not U34623(n32850,n32846);
  nand U34624(n32846,n32777,n32541);
  nand U34625(n32851,n32847,n32845);
  nand U34626(n32845,n32434,n32853);
  nand U34627(n32853,n29978,n31458,n32417);
  nand U34628(n29978,n32854,n32441);
  nor U34629(n32441,n32855,n32856);
  not U34630(n32847,n32786);
  nand U34631(n32786,n32545,n32776);
  nand U34632(G2460,n32857,n32858,n32859,n32860);
  nor U34633(n32860,n32861,n32862,n32863);
  nor U34634(n32863,n26769,n32864);
  nor U34635(n32862,n32342,n32865);
  nor U34636(n32861,n29976,n32344);
  nand U34637(n32859,n32866,G59059);
  nand U34638(n32858,n32346,n32867);
  nand U34639(n32857,G58871,n32868);
  nand U34640(G2459,n32869,n32870,n32871,n32872);
  nor U34641(n32872,n32873,n32874,n32875);
  nor U34642(n32875,n26792,n32864);
  nor U34643(n32874,n32356,n32865);
  nor U34644(n32873,n29976,n32357);
  nand U34645(n32871,n32866,G59058);
  nand U34646(n32870,n32358,n32867);
  nand U34647(n32869,G58872,n32868);
  nand U34648(G2458,n32876,n32877,n32878,n32879);
  nor U34649(n32879,n32880,n32881,n32882);
  nor U34650(n32882,n26809,n32864);
  nor U34651(n32881,n32366,n32865);
  nor U34652(n32880,n29976,n32367);
  nand U34653(n32878,n32866,G59057);
  nand U34654(n32877,n32368,n32867);
  nand U34655(n32876,G58873,n32868);
  nand U34656(G2457,n32883,n32884,n32885,n32886);
  nor U34657(n32886,n32887,n32888,n32889);
  nor U34658(n32889,n26826,n32864);
  nor U34659(n32888,n32376,n32865);
  nor U34660(n32887,n29976,n32377);
  nand U34661(n32885,n32866,G59056);
  nand U34662(n32884,n32378,n32867);
  nand U34663(n32883,G58874,n32868);
  nand U34664(G2456,n32890,n32891,n32892,n32893);
  nor U34665(n32893,n32894,n32895,n32896);
  nor U34666(n32896,n26843,n32864);
  nor U34667(n32895,n32386,n32865);
  nor U34668(n32894,n29976,n32387);
  nand U34669(n32892,n32866,G59055);
  nand U34670(n32891,n32388,n32867);
  nand U34671(n32890,G58875,n32868);
  nand U34672(G2455,n32897,n32898,n32899,n32900);
  nor U34673(n32900,n32901,n32902,n32903);
  nor U34674(n32903,n26860,n32864);
  nor U34675(n32902,n32396,n32865);
  nor U34676(n32901,n29976,n32397);
  nand U34677(n32899,n32866,G59054);
  nand U34678(n32898,n32398,n32867);
  nand U34679(n32897,G58876,n32868);
  nand U34680(G2454,n32904,n32905,n32906,n32907);
  nor U34681(n32907,n32908,n32909,n32910);
  nor U34682(n32910,n26878,n32864);
  nor U34683(n32909,n32406,n32865);
  nor U34684(n32908,n29976,n32407);
  nand U34685(n32906,n32866,G59053);
  nand U34686(n32905,n32408,n32867);
  nand U34687(n32904,G58877,n32868);
  nand U34688(G2453,n32911,n32912,n32913,n32914);
  nor U34689(n32914,n32915,n32916,n32917);
  nor U34690(n32917,n26905,n32864);
  nand U34691(n32864,n32918,n29976,n32417);
  nor U34692(n32916,n32418,n32865);
  nor U34693(n32915,n29976,n32419);
  nand U34694(n32913,n32866,G59052);
  and U34695(n32866,n32919,n32920);
  nand U34696(n32920,n32921,n32423,n32922);
  nand U34697(n32922,G58977,n31436);
  nand U34698(n32921,n32923,n32924);
  nand U34699(n32919,n32925,n32428);
  nand U34700(n32912,n32429,n32867);
  nand U34701(n32867,n32926,n32927);
  or U34702(n32927,n32924,n29174);
  nand U34703(n32926,n32918,G58977);
  not U34704(n32918,n31436);
  nand U34705(n32911,G58878,n32868);
  nand U34706(n32868,n32928,n32929);
  nand U34707(n32929,n32925,n32923);
  nand U34708(n32923,n32434,n32930);
  not U34709(n32925,n32865);
  nand U34710(n32865,n32620,n32776);
  or U34711(n32928,n32930,n32924);
  nand U34712(n32924,n32777,n32621);
  nand U34713(n32930,n29976,n31436,n32417);
  nand U34714(n29976,n32778,n32622);
  nand U34715(G2452,n32931,n32932,n32933,n32934);
  nor U34716(n32934,n32935,n32936,n32937);
  nor U34717(n32937,n26769,n32938);
  nor U34718(n32936,n29974,n32344);
  nor U34719(n32935,n32342,n32939);
  nand U34720(n32933,n32940,G59051);
  nand U34721(n32932,n32346,n32941);
  nand U34722(n32931,G58871,n32942);
  nand U34723(G2451,n32943,n32944,n32945,n32946);
  nor U34724(n32946,n32947,n32948,n32949);
  nor U34725(n32949,n26792,n32938);
  nor U34726(n32948,n29974,n32357);
  nor U34727(n32947,n32356,n32939);
  nand U34728(n32945,n32940,G59050);
  nand U34729(n32944,n32358,n32941);
  nand U34730(n32943,G58872,n32942);
  nand U34731(G2450,n32950,n32951,n32952,n32953);
  nor U34732(n32953,n32954,n32955,n32956);
  nor U34733(n32956,n26809,n32938);
  nor U34734(n32955,n29974,n32367);
  nor U34735(n32954,n32366,n32939);
  nand U34736(n32952,n32940,G59049);
  nand U34737(n32951,n32368,n32941);
  nand U34738(n32950,G58873,n32942);
  nand U34739(G2449,n32957,n32958,n32959,n32960);
  nor U34740(n32960,n32961,n32962,n32963);
  nor U34741(n32963,n26826,n32938);
  nor U34742(n32962,n29974,n32377);
  nor U34743(n32961,n32376,n32939);
  nand U34744(n32959,n32940,G59048);
  nand U34745(n32958,n32378,n32941);
  nand U34746(n32957,G58874,n32942);
  nand U34747(G2448,n32964,n32965,n32966,n32967);
  nor U34748(n32967,n32968,n32969,n32970);
  nor U34749(n32970,n26843,n32938);
  nor U34750(n32969,n29974,n32387);
  nor U34751(n32968,n32386,n32939);
  nand U34752(n32966,n32940,G59047);
  nand U34753(n32965,n32388,n32941);
  nand U34754(n32964,G58875,n32942);
  nand U34755(G2447,n32971,n32972,n32973,n32974);
  nor U34756(n32974,n32975,n32976,n32977);
  nor U34757(n32977,n26860,n32938);
  nor U34758(n32976,n29974,n32397);
  nor U34759(n32975,n32396,n32939);
  nand U34760(n32973,n32940,G59046);
  nand U34761(n32972,n32398,n32941);
  nand U34762(n32971,G58876,n32942);
  nand U34763(G2446,n32978,n32979,n32980,n32981);
  nor U34764(n32981,n32982,n32983,n32984);
  nor U34765(n32984,n26878,n32938);
  nor U34766(n32983,n29974,n32407);
  nor U34767(n32982,n32406,n32939);
  nand U34768(n32980,n32940,G59045);
  nand U34769(n32979,n32408,n32941);
  nand U34770(n32978,G58877,n32942);
  nand U34771(G2445,n32985,n32986,n32987,n32988);
  nor U34772(n32988,n32989,n32990,n32991);
  nor U34773(n32991,n26905,n32938);
  nand U34774(n32938,n32417,n32992);
  nor U34775(n32990,n29974,n32419);
  nor U34776(n32989,n32418,n32939);
  nand U34777(n32987,n32940,G59044);
  and U34778(n32940,n32993,n32994);
  nand U34779(n32994,n32995,n32423,n32996);
  nand U34780(n32996,G58977,n31441);
  nand U34781(n32995,n32997,n32998);
  nand U34782(n32993,n32999,n32428);
  nand U34783(n32986,n32429,n32941);
  nand U34784(n32941,n33000,n33001);
  nand U34785(n33001,n33002,n29226);
  nand U34786(n33000,n32992,G58977);
  not U34787(n32992,n31441);
  nand U34788(n32985,G58878,n32942);
  nand U34789(n32942,n33003,n33004);
  nand U34790(n33004,n32417,n29974,n33002);
  not U34791(n33002,n32998);
  nand U34792(n32998,n32777,n32697);
  nor U34793(n32777,n32698,n33005);
  nand U34794(n33003,n32999,n32997);
  nand U34795(n32997,n32434,n33006);
  nand U34796(n33006,n29974,n31441,n32417);
  nand U34797(n29974,n32854,n32622);
  nor U34798(n32622,n32856,n33007);
  nand U34799(G2444,n33008,n33009,n33010,n33011);
  nor U34800(n33011,n33012,n33013,n33014);
  nor U34801(n33014,n26769,n33015);
  nor U34802(n33013,n32342,n33016);
  nor U34803(n33012,n29988,n32344);
  nand U34804(n33010,n33017,G59043);
  nand U34805(n33009,n32346,n33018);
  nand U34806(n33008,G58871,n33019);
  nand U34807(G2443,n33020,n33021,n33022,n33023);
  nor U34808(n33023,n33024,n33025,n33026);
  nor U34809(n33026,n26792,n33015);
  nor U34810(n33025,n32356,n33016);
  nor U34811(n33024,n29988,n32357);
  nand U34812(n33022,n33017,G59042);
  nand U34813(n33021,n32358,n33018);
  nand U34814(n33020,G58872,n33019);
  nand U34815(G2442,n33027,n33028,n33029,n33030);
  nor U34816(n33030,n33031,n33032,n33033);
  nor U34817(n33033,n26809,n33015);
  nor U34818(n33032,n32366,n33016);
  nor U34819(n33031,n29988,n32367);
  nand U34820(n33029,n33017,G59041);
  nand U34821(n33028,n32368,n33018);
  nand U34822(n33027,G58873,n33019);
  nand U34823(G2441,n33034,n33035,n33036,n33037);
  nor U34824(n33037,n33038,n33039,n33040);
  nor U34825(n33040,n26826,n33015);
  nor U34826(n33039,n32376,n33016);
  nor U34827(n33038,n29988,n32377);
  nand U34828(n33036,n33017,G59040);
  nand U34829(n33035,n32378,n33018);
  nand U34830(n33034,G58874,n33019);
  nand U34831(G2440,n33041,n33042,n33043,n33044);
  nor U34832(n33044,n33045,n33046,n33047);
  nor U34833(n33047,n26843,n33015);
  nor U34834(n33046,n32386,n33016);
  nor U34835(n33045,n29988,n32387);
  nand U34836(n33043,n33017,G59039);
  nand U34837(n33042,n32388,n33018);
  nand U34838(n33041,G58875,n33019);
  nand U34839(G2439,n33048,n33049,n33050,n33051);
  nor U34840(n33051,n33052,n33053,n33054);
  nor U34841(n33054,n26860,n33015);
  nor U34842(n33053,n32396,n33016);
  nor U34843(n33052,n29988,n32397);
  nand U34844(n33050,n33017,G59038);
  nand U34845(n33049,n32398,n33018);
  nand U34846(n33048,G58876,n33019);
  nand U34847(G2438,n33055,n33056,n33057,n33058);
  nor U34848(n33058,n33059,n33060,n33061);
  nor U34849(n33061,n26878,n33015);
  nor U34850(n33060,n32406,n33016);
  nor U34851(n33059,n29988,n32407);
  nand U34852(n33057,n33017,G59037);
  nand U34853(n33056,n32408,n33018);
  nand U34854(n33055,G58877,n33019);
  nand U34855(G2437,n33062,n33063,n33064,n33065);
  nor U34856(n33065,n33066,n33067,n33068);
  nor U34857(n33068,n26905,n33015);
  nand U34858(n33015,n33069,n29988,n32417);
  nor U34859(n33067,n32418,n33016);
  nor U34860(n33066,n29988,n32419);
  nand U34861(n33064,n33017,G59036);
  and U34862(n33017,n33070,n33071);
  nand U34863(n33071,n33072,n32423,n33073);
  nand U34864(n33073,G58977,n31442);
  nand U34865(n33072,n33074,n33075);
  nand U34866(n33070,n33076,n32428);
  nand U34867(n33063,n32429,n33018);
  nand U34868(n33018,n33077,n33078);
  or U34869(n33078,n33075,n29174);
  nand U34870(n33077,n33069,G58977);
  not U34871(n33069,n31442);
  nand U34872(n33062,G58878,n33019);
  nand U34873(n33019,n33079,n33080);
  nand U34874(n33080,n33076,n33074);
  nand U34875(n33074,n32434,n33081);
  not U34876(n33076,n33016);
  nand U34877(n33016,n33082,n32436);
  or U34878(n33079,n33081,n33075);
  nand U34879(n33075,n33083,n32438);
  nand U34880(n33081,n29988,n31442,n32417);
  nand U34881(n29988,n33084,n32440);
  nand U34882(G2436,n33085,n33086,n33087,n33088);
  nor U34883(n33088,n33089,n33090,n33091);
  nor U34884(n33091,n33092,n26779);
  nor U34885(n33090,n33093,n32451);
  nor U34886(n33089,n29926,n33094);
  nand U34887(n33087,n33095,G58887);
  nand U34888(n33086,n32454,n33096);
  nand U34889(n33085,n33097,n32457);
  nand U34890(G2435,n33098,n33099,n33100,n33101);
  nor U34891(n33101,n33102,n33103,n33104);
  nor U34892(n33104,n33092,n26797);
  nor U34893(n33103,n33093,n32465);
  nor U34894(n33102,n29840,n33094);
  nand U34895(n33100,n33095,G58888);
  nand U34896(n33099,n32466,n33096);
  nand U34897(n33098,n33097,n32467);
  nand U34898(G2434,n33105,n33106,n33107,n33108);
  nor U34899(n33108,n33109,n33110,n33111);
  nor U34900(n33111,n33092,n26814);
  nor U34901(n33110,n33093,n32475);
  nor U34902(n33109,n29744,n33094);
  nand U34903(n33107,n33095,G58889);
  nand U34904(n33106,n32476,n33096);
  nand U34905(n33105,n33097,n32477);
  nand U34906(G2433,n33112,n33113,n33114,n33115);
  nor U34907(n33115,n33116,n33117,n33118);
  nor U34908(n33118,n33092,n26831);
  nor U34909(n33117,n33093,n32485);
  nor U34910(n33116,n29675,n33094);
  nand U34911(n33114,n33095,G58890);
  nand U34912(n33113,n32486,n33096);
  nand U34913(n33112,n33097,n32487);
  nand U34914(G2432,n33119,n33120,n33121,n33122);
  nor U34915(n33122,n33123,n33124,n33125);
  nor U34916(n33125,n33092,n26848);
  nor U34917(n33124,n33093,n32495);
  nor U34918(n33123,n29599,n33094);
  nand U34919(n33121,n33095,G58891);
  nand U34920(n33120,n32496,n33096);
  nand U34921(n33119,n33097,n32497);
  nand U34922(G2431,n33126,n33127,n33128,n33129);
  nor U34923(n33129,n33130,n33131,n33132);
  nor U34924(n33132,n33092,n26866);
  nor U34925(n33131,n33093,n32505);
  nor U34926(n33130,n29520,n33094);
  nand U34927(n33128,n33095,G58892);
  nand U34928(n33127,n32506,n33096);
  nand U34929(n33126,n33097,n32507);
  nand U34930(G2430,n33133,n33134,n33135,n33136);
  nor U34931(n33136,n33137,n33138,n33139);
  nor U34932(n33139,n33092,n26883);
  nor U34933(n33138,n33093,n32515);
  nor U34934(n33137,n29416,n33094);
  nand U34935(n33135,n33095,G58893);
  nand U34936(n33134,n32516,n33096);
  nand U34937(n33133,n33097,n32517);
  nand U34938(G2429,n33140,n33141,n33142,n33143);
  nor U34939(n33143,n33144,n33145,n33146);
  nor U34940(n33146,n33092,n26913);
  and U34941(n33092,n33147,n33148);
  nand U34942(n33148,n33149,n29987,n32417);
  nand U34943(n33149,n33150,n33151);
  nand U34944(n33147,n33097,n32530);
  nor U34945(n33145,n33093,n32531);
  and U34946(n33093,n33152,n33153);
  or U34947(n33153,n33151,n29174);
  nand U34948(n33152,n33154,G58977);
  nor U34949(n33144,n29345,n33094);
  nand U34950(n33094,n33155,n33156);
  nand U34951(n33156,n33157,n32423,n33158);
  nand U34952(n33158,n32530,n33151);
  nand U34953(n33157,n33159,n31459);
  nand U34954(n33159,n33160,n27929);
  nand U34955(n33160,n33151,n29987);
  nand U34956(n33151,n33083,n32541);
  nand U34957(n33155,n33097,n32428);
  nand U34958(n33142,n33095,G58894);
  and U34959(n33095,n32417,n33154);
  not U34960(n33154,n31459);
  nand U34961(n33141,n32542,n33096);
  not U34962(n33096,n29987);
  nand U34963(n29987,n33084,n32543);
  nand U34964(n33140,n33097,n32544);
  not U34965(n33097,n33150);
  nand U34966(n33150,n33082,n32545);
  nand U34967(G2428,n33161,n33162,n33163,n33164);
  nor U34968(n33164,n33165,n33166,n33167);
  nor U34969(n33167,n26769,n33168);
  nor U34970(n33166,n32342,n33169);
  nor U34971(n33165,n29986,n32344);
  nand U34972(n33163,n33170,G59027);
  nand U34973(n33162,n32346,n33171);
  nand U34974(n33161,G58871,n33172);
  nand U34975(G2427,n33173,n33174,n33175,n33176);
  nor U34976(n33176,n33177,n33178,n33179);
  nor U34977(n33179,n26792,n33168);
  nor U34978(n33178,n32356,n33169);
  nor U34979(n33177,n29986,n32357);
  nand U34980(n33175,n33170,G59026);
  nand U34981(n33174,n32358,n33171);
  nand U34982(n33173,G58872,n33172);
  nand U34983(G2426,n33180,n33181,n33182,n33183);
  nor U34984(n33183,n33184,n33185,n33186);
  nor U34985(n33186,n26809,n33168);
  nor U34986(n33185,n32366,n33169);
  nor U34987(n33184,n29986,n32367);
  nand U34988(n33182,n33170,G59025);
  nand U34989(n33181,n32368,n33171);
  nand U34990(n33180,G58873,n33172);
  nand U34991(G2425,n33187,n33188,n33189,n33190);
  nor U34992(n33190,n33191,n33192,n33193);
  nor U34993(n33193,n26826,n33168);
  nor U34994(n33192,n32376,n33169);
  nor U34995(n33191,n29986,n32377);
  nand U34996(n33189,n33170,G59024);
  nand U34997(n33188,n32378,n33171);
  nand U34998(n33187,G58874,n33172);
  nand U34999(G2424,n33194,n33195,n33196,n33197);
  nor U35000(n33197,n33198,n33199,n33200);
  nor U35001(n33200,n26843,n33168);
  nor U35002(n33199,n32386,n33169);
  nor U35003(n33198,n29986,n32387);
  nand U35004(n33196,n33170,G59023);
  nand U35005(n33195,n32388,n33171);
  nand U35006(n33194,G58875,n33172);
  nand U35007(G2423,n33201,n33202,n33203,n33204);
  nor U35008(n33204,n33205,n33206,n33207);
  nor U35009(n33207,n26860,n33168);
  nor U35010(n33206,n32396,n33169);
  nor U35011(n33205,n29986,n32397);
  nand U35012(n33203,n33170,G59022);
  nand U35013(n33202,n32398,n33171);
  nand U35014(n33201,G58876,n33172);
  nand U35015(G2422,n33208,n33209,n33210,n33211);
  nor U35016(n33211,n33212,n33213,n33214);
  nor U35017(n33214,n26878,n33168);
  nor U35018(n33213,n32406,n33169);
  nor U35019(n33212,n29986,n32407);
  nand U35020(n33210,n33170,G59021);
  nand U35021(n33209,n32408,n33171);
  nand U35022(n33208,G58877,n33172);
  nand U35023(G2421,n33215,n33216,n33217,n33218);
  nor U35024(n33218,n33219,n33220,n33221);
  nor U35025(n33221,n26905,n33168);
  nand U35026(n33168,n33222,n29986,n32417);
  nor U35027(n33220,n32418,n33169);
  nor U35028(n33219,n29986,n32419);
  nand U35029(n33217,n33170,G59020);
  and U35030(n33170,n33223,n33224);
  nand U35031(n33224,n33225,n32423,n33226);
  nand U35032(n33226,G58977,n31443);
  nand U35033(n33225,n33227,n33228);
  nand U35034(n33223,n33229,n32428);
  nand U35035(n33216,n32429,n33171);
  nand U35036(n33171,n33230,n33231);
  or U35037(n33231,n33228,n29174);
  nand U35038(n33230,n33222,G58977);
  not U35039(n33222,n31443);
  nand U35040(n33215,G58878,n33172);
  nand U35041(n33172,n33232,n33233);
  nand U35042(n33233,n33229,n33227);
  nand U35043(n33227,n32434,n33234);
  not U35044(n33229,n33169);
  nand U35045(n33169,n33082,n32620);
  or U35046(n33232,n33234,n33228);
  nand U35047(n33228,n33083,n32621);
  nand U35048(n33234,n29986,n31443,n32417);
  nand U35049(n29986,n33235,n32440);
  and U35050(n32440,n33236,n33237);
  nand U35051(G2420,n33238,n33239,n33240,n33241);
  nor U35052(n33241,n33242,n33243,n33244);
  nor U35053(n33244,n32342,n33245);
  nor U35054(n33243,n29985,n32344);
  nor U35055(n33242,n26769,n33246);
  nand U35056(n33240,n33247,G59019);
  nand U35057(n33239,n32346,n33248);
  nand U35058(n33238,G58871,n33249);
  nand U35059(G2419,n33250,n33251,n33252,n33253);
  nor U35060(n33253,n33254,n33255,n33256);
  nor U35061(n33256,n32356,n33245);
  nor U35062(n33255,n29985,n32357);
  nor U35063(n33254,n26792,n33246);
  nand U35064(n33252,n33247,G59018);
  nand U35065(n33251,n32358,n33248);
  nand U35066(n33250,G58872,n33249);
  nand U35067(G2418,n33257,n33258,n33259,n33260);
  nor U35068(n33260,n33261,n33262,n33263);
  nor U35069(n33263,n32366,n33245);
  nor U35070(n33262,n29985,n32367);
  nor U35071(n33261,n26809,n33246);
  nand U35072(n33259,n33247,G59017);
  nand U35073(n33258,n32368,n33248);
  nand U35074(n33257,G58873,n33249);
  nand U35075(G2417,n33264,n33265,n33266,n33267);
  nor U35076(n33267,n33268,n33269,n33270);
  nor U35077(n33270,n32376,n33245);
  nor U35078(n33269,n29985,n32377);
  nor U35079(n33268,n26826,n33246);
  nand U35080(n33266,n33247,G59016);
  nand U35081(n33265,n32378,n33248);
  nand U35082(n33264,G58874,n33249);
  nand U35083(G2416,n33271,n33272,n33273,n33274);
  nor U35084(n33274,n33275,n33276,n33277);
  nor U35085(n33277,n32386,n33245);
  nor U35086(n33276,n29985,n32387);
  nor U35087(n33275,n26843,n33246);
  nand U35088(n33273,n33247,G59015);
  nand U35089(n33272,n32388,n33248);
  nand U35090(n33271,G58875,n33249);
  nand U35091(G2415,n33278,n33279,n33280,n33281);
  nor U35092(n33281,n33282,n33283,n33284);
  nor U35093(n33284,n32396,n33245);
  nor U35094(n33283,n29985,n32397);
  nor U35095(n33282,n26860,n33246);
  nand U35096(n33280,n33247,G59014);
  nand U35097(n33279,n32398,n33248);
  nand U35098(n33278,G58876,n33249);
  nand U35099(G2414,n33285,n33286,n33287,n33288);
  nor U35100(n33288,n33289,n33290,n33291);
  nor U35101(n33291,n32406,n33245);
  nor U35102(n33290,n29985,n32407);
  nor U35103(n33289,n26878,n33246);
  nand U35104(n33287,n33247,G59013);
  nand U35105(n33286,n32408,n33248);
  nand U35106(n33285,G58877,n33249);
  nand U35107(G2413,n33292,n33293,n33294,n33295);
  nor U35108(n33295,n33296,n33297,n33298);
  nor U35109(n33298,n32418,n33245);
  nor U35110(n33297,n29985,n32419);
  nor U35111(n33296,n26905,n33246);
  nand U35112(n33246,n32417,n33299);
  nand U35113(n33294,n33247,G59012);
  and U35114(n33247,n33300,n33301);
  nand U35115(n33301,n33302,n32423,n33303);
  nand U35116(n33303,G58977,n31444);
  nand U35117(n33302,n33304,n33305);
  nand U35118(n33300,n33306,n32428);
  nand U35119(n33293,n32429,n33248);
  nand U35120(n33248,n33307,n33308);
  nand U35121(n33308,n33309,n29226);
  nand U35122(n33307,n33299,G58977);
  not U35123(n33299,n31444);
  nand U35124(n33292,G58878,n33249);
  nand U35125(n33249,n33310,n33311);
  nand U35126(n33311,n32417,n29985,n33309);
  not U35127(n33309,n33305);
  nand U35128(n33305,n33083,n32697);
  nor U35129(n33083,n32699,n33312);
  nand U35130(n33310,n33306,n33304);
  nand U35131(n33304,n32434,n33313);
  nand U35132(n33313,n29985,n31444,n32417);
  nand U35133(n29985,n33235,n32543);
  and U35134(n32543,n33314,n33236);
  not U35135(n33306,n33245);
  nand U35136(n33245,n33082,n32701);
  nand U35137(G2412,n33315,n33316,n33317,n33318);
  nor U35138(n33318,n33319,n33320,n33321);
  nor U35139(n33321,n26769,n33322);
  nor U35140(n33320,n32342,n33323);
  nor U35141(n33319,n29996,n32344);
  nand U35142(n33317,n33324,G59011);
  nand U35143(n33316,n32346,n33325);
  nand U35144(n33315,G58871,n33326);
  nand U35145(G2411,n33327,n33328,n33329,n33330);
  nor U35146(n33330,n33331,n33332,n33333);
  nor U35147(n33333,n26792,n33322);
  nor U35148(n33332,n32356,n33323);
  nor U35149(n33331,n29996,n32357);
  nand U35150(n33329,n33324,G59010);
  nand U35151(n33328,n32358,n33325);
  nand U35152(n33327,G58872,n33326);
  nand U35153(G2410,n33334,n33335,n33336,n33337);
  nor U35154(n33337,n33338,n33339,n33340);
  nor U35155(n33340,n26809,n33322);
  nor U35156(n33339,n32366,n33323);
  nor U35157(n33338,n29996,n32367);
  nand U35158(n33336,n33324,G59009);
  nand U35159(n33335,n32368,n33325);
  nand U35160(n33334,G58873,n33326);
  nand U35161(G2409,n33341,n33342,n33343,n33344);
  nor U35162(n33344,n33345,n33346,n33347);
  nor U35163(n33347,n26826,n33322);
  nor U35164(n33346,n32376,n33323);
  nor U35165(n33345,n29996,n32377);
  nand U35166(n33343,n33324,G59008);
  nand U35167(n33342,n32378,n33325);
  nand U35168(n33341,G58874,n33326);
  nand U35169(G2408,n33348,n33349,n33350,n33351);
  nor U35170(n33351,n33352,n33353,n33354);
  nor U35171(n33354,n26843,n33322);
  nor U35172(n33353,n32386,n33323);
  nor U35173(n33352,n29996,n32387);
  nand U35174(n33350,n33324,G59007);
  nand U35175(n33349,n32388,n33325);
  nand U35176(n33348,G58875,n33326);
  nand U35177(G2407,n33355,n33356,n33357,n33358);
  nor U35178(n33358,n33359,n33360,n33361);
  nor U35179(n33361,n26860,n33322);
  nor U35180(n33360,n32396,n33323);
  nor U35181(n33359,n29996,n32397);
  nand U35182(n33357,n33324,G59006);
  nand U35183(n33356,n32398,n33325);
  nand U35184(n33355,G58876,n33326);
  nand U35185(G2406,n33362,n33363,n33364,n33365);
  nor U35186(n33365,n33366,n33367,n33368);
  nor U35187(n33368,n26878,n33322);
  nor U35188(n33367,n32406,n33323);
  nor U35189(n33366,n29996,n32407);
  nand U35190(n33364,n33324,G59005);
  nand U35191(n33363,n32408,n33325);
  nand U35192(n33362,G58877,n33326);
  nand U35193(G2405,n33369,n33370,n33371,n33372);
  nor U35194(n33372,n33373,n33374,n33375);
  nor U35195(n33375,n26905,n33322);
  nand U35196(n33322,n33376,n29996,n32417);
  nor U35197(n33374,n32418,n33323);
  nor U35198(n33373,n29996,n32419);
  nand U35199(n33371,n33324,G59004);
  and U35200(n33324,n33377,n33378);
  nand U35201(n33378,n33379,n32423,n33380);
  nand U35202(n33380,G58977,n31449);
  nand U35203(n33379,n33381,n33382);
  nand U35204(n33377,n33383,n32428);
  nand U35205(n33370,n32429,n33325);
  nand U35206(n33325,n33384,n33385);
  or U35207(n33385,n33382,n29174);
  nand U35208(n33384,n33376,G58977);
  not U35209(n33376,n31449);
  nand U35210(n33369,G58878,n33326);
  nand U35211(n33326,n33386,n33387);
  nand U35212(n33387,n33383,n33381);
  nand U35213(n33381,n32434,n33388);
  not U35214(n33383,n33323);
  nand U35215(n33323,n33389,n32436);
  nor U35216(n32436,G59117,G59116);
  or U35217(n33386,n33388,n33382);
  nand U35218(n33382,n33390,n32438);
  nor U35219(n32438,n33391,n33392);
  nand U35220(n33388,n29996,n31449,n32417);
  nand U35221(n29996,n33084,n32778);
  nand U35222(G2404,n33393,n33394,n33395,n33396);
  nor U35223(n33396,n33397,n33398,n33399);
  nor U35224(n33399,n33400,n26779);
  nor U35225(n33398,n33401,n32451);
  nor U35226(n33397,n29913,n33402);
  nand U35227(n33395,n33403,G58887);
  nand U35228(n33394,n32454,n33404);
  not U35229(n32454,n32344);
  nand U35230(n33393,n33405,n32457);
  nand U35231(G2403,n33406,n33407,n33408,n33409);
  nor U35232(n33409,n33410,n33411,n33412);
  nor U35233(n33412,n33400,n26797);
  nor U35234(n33411,n33401,n32465);
  nor U35235(n33410,n29832,n33402);
  nand U35236(n33408,n33403,G58888);
  nand U35237(n33407,n32466,n33404);
  not U35238(n32466,n32357);
  nand U35239(n33406,n33405,n32467);
  nand U35240(G2402,n33413,n33414,n33415,n33416);
  nor U35241(n33416,n33417,n33418,n33419);
  nor U35242(n33419,n33400,n26814);
  nor U35243(n33418,n33401,n32475);
  nor U35244(n33417,n29736,n33402);
  nand U35245(n33415,n33403,G58889);
  nand U35246(n33414,n32476,n33404);
  not U35247(n32476,n32367);
  nand U35248(n33413,n33405,n32477);
  nand U35249(G2401,n33420,n33421,n33422,n33423);
  nor U35250(n33423,n33424,n33425,n33426);
  nor U35251(n33426,n33400,n26831);
  nor U35252(n33425,n33401,n32485);
  nor U35253(n33424,n29667,n33402);
  nand U35254(n33422,n33403,G58890);
  nand U35255(n33421,n32486,n33404);
  not U35256(n32486,n32377);
  nand U35257(n33420,n33405,n32487);
  nand U35258(G2400,n33427,n33428,n33429,n33430);
  nor U35259(n33430,n33431,n33432,n33433);
  nor U35260(n33433,n33400,n26848);
  nor U35261(n33432,n33401,n32495);
  nor U35262(n33431,n29591,n33402);
  nand U35263(n33429,n33403,G58891);
  nand U35264(n33428,n32496,n33404);
  not U35265(n32496,n32387);
  nand U35266(n33427,n33405,n32497);
  nand U35267(G2399,n33434,n33435,n33436,n33437);
  nor U35268(n33437,n33438,n33439,n33440);
  nor U35269(n33440,n33400,n26866);
  nor U35270(n33439,n33401,n32505);
  nor U35271(n33438,n29512,n33402);
  nand U35272(n33436,n33403,G58892);
  nand U35273(n33435,n32506,n33404);
  not U35274(n32506,n32397);
  nand U35275(n33434,n33405,n32507);
  nand U35276(G2398,n33441,n33442,n33443,n33444);
  nor U35277(n33444,n33445,n33446,n33447);
  nor U35278(n33447,n33400,n26883);
  nor U35279(n33446,n33401,n32515);
  nor U35280(n33445,n29408,n33402);
  nand U35281(n33443,n33403,G58893);
  nand U35282(n33442,n32516,n33404);
  not U35283(n32516,n32407);
  nand U35284(n33441,n33405,n32517);
  nand U35285(G2397,n33448,n33449,n33450,n33451);
  nor U35286(n33451,n33452,n33453,n33454);
  nor U35287(n33454,n33400,n26913);
  and U35288(n33400,n33455,n33456);
  nand U35289(n33456,n33457,n29995,n32417);
  nand U35290(n33457,n33458,n33459);
  nand U35291(n33455,n33405,n32530);
  nor U35292(n33453,n33401,n32531);
  and U35293(n33401,n33460,n33461);
  or U35294(n33461,n33459,n29174);
  nand U35295(n33460,n33462,G58977);
  nor U35296(n33452,n29333,n33402);
  nand U35297(n33402,n33463,n33464);
  nand U35298(n33464,n33465,n32423,n33466);
  nand U35299(n33466,n32530,n33459);
  nand U35300(n33465,n33467,n31460);
  nand U35301(n33467,n33468,n27929);
  nand U35302(n33468,n33459,n29995);
  nand U35303(n33459,n33390,n32541);
  nor U35304(n32541,n33391,G59117);
  nand U35305(n33463,n33405,n32428);
  nand U35306(n33450,n33403,G58894);
  and U35307(n33403,n32417,n33462);
  not U35308(n33462,n31460);
  nand U35309(n33449,n32542,n33404);
  not U35310(n33404,n29995);
  nand U35311(n29995,n33084,n32854);
  nor U35312(n33084,n32855,n33469);
  not U35313(n32542,n32419);
  nand U35314(n33448,n33405,n32544);
  not U35315(n33405,n33458);
  nand U35316(n33458,n33389,n32545);
  nand U35317(G2396,n33470,n33471,n33472,n33473);
  nor U35318(n33473,n33474,n33475,n33476);
  nor U35319(n33476,n26769,n33477);
  not U35320(n26769,G58887);
  nor U35321(n33475,n32342,n33478);
  nor U35322(n33474,n29994,n32344);
  nand U35323(n33472,n33479,G58995);
  nand U35324(n33471,n32346,n33480);
  nand U35325(n33470,G58871,n33481);
  nand U35326(G2395,n33482,n33483,n33484,n33485);
  nor U35327(n33485,n33486,n33487,n33488);
  nor U35328(n33488,n26792,n33477);
  not U35329(n26792,G58888);
  nor U35330(n33487,n32356,n33478);
  nor U35331(n33486,n29994,n32357);
  nand U35332(n33484,n33479,G58994);
  nand U35333(n33483,n32358,n33480);
  nand U35334(n33482,G58872,n33481);
  nand U35335(G2394,n33489,n33490,n33491,n33492);
  nor U35336(n33492,n33493,n33494,n33495);
  nor U35337(n33495,n26809,n33477);
  not U35338(n26809,G58889);
  nor U35339(n33494,n32366,n33478);
  nor U35340(n33493,n29994,n32367);
  nand U35341(n33491,n33479,G58993);
  nand U35342(n33490,n32368,n33480);
  nand U35343(n33489,G58873,n33481);
  nand U35344(G2393,n33496,n33497,n33498,n33499);
  nor U35345(n33499,n33500,n33501,n33502);
  nor U35346(n33502,n26826,n33477);
  not U35347(n26826,G58890);
  nor U35348(n33501,n32376,n33478);
  nor U35349(n33500,n29994,n32377);
  nand U35350(n33498,n33479,G58992);
  nand U35351(n33497,n32378,n33480);
  nand U35352(n33496,G58874,n33481);
  nand U35353(G2392,n33503,n33504,n33505,n33506);
  nor U35354(n33506,n33507,n33508,n33509);
  nor U35355(n33509,n26843,n33477);
  not U35356(n26843,G58891);
  nor U35357(n33508,n32386,n33478);
  nor U35358(n33507,n29994,n32387);
  nand U35359(n33505,n33479,G58991);
  nand U35360(n33504,n32388,n33480);
  nand U35361(n33503,G58875,n33481);
  nand U35362(G2391,n33510,n33511,n33512,n33513);
  nor U35363(n33513,n33514,n33515,n33516);
  nor U35364(n33516,n26860,n33477);
  not U35365(n26860,G58892);
  nor U35366(n33515,n32396,n33478);
  nor U35367(n33514,n29994,n32397);
  nand U35368(n33512,n33479,G58990);
  nand U35369(n33511,n32398,n33480);
  nand U35370(n33510,G58876,n33481);
  nand U35371(G2390,n33517,n33518,n33519,n33520);
  nor U35372(n33520,n33521,n33522,n33523);
  nor U35373(n33523,n26878,n33477);
  not U35374(n26878,G58893);
  nor U35375(n33522,n32406,n33478);
  nor U35376(n33521,n29994,n32407);
  nand U35377(n33519,n33479,G58989);
  nand U35378(n33518,n32408,n33480);
  nand U35379(n33517,G58877,n33481);
  nand U35380(G2389,n33524,n33525,n33526,n33527);
  nor U35381(n33527,n33528,n33529,n33530);
  nor U35382(n33530,n26905,n33477);
  nand U35383(n33477,n33531,n29994,n32417);
  not U35384(n26905,G58894);
  nor U35385(n33529,n32418,n33478);
  nor U35386(n33528,n29994,n32419);
  nand U35387(n33526,n33479,G58988);
  and U35388(n33479,n33532,n33533);
  nand U35389(n33533,n33534,n32423,n33535);
  nand U35390(n33535,G58977,n31450);
  nand U35391(n33534,n33536,n33537);
  nand U35392(n33532,n33538,n32428);
  nand U35393(n33525,n32429,n33480);
  nand U35394(n33480,n33539,n33540);
  or U35395(n33540,n33537,n29174);
  nand U35396(n33539,n33531,G58977);
  not U35397(n33531,n31450);
  nand U35398(n33524,G58878,n33481);
  nand U35399(n33481,n33541,n33542);
  nand U35400(n33542,n33538,n33536);
  nand U35401(n33536,n32434,n33543);
  not U35402(n33538,n33478);
  nand U35403(n33478,n33389,n32620);
  or U35404(n33541,n33543,n33537);
  nand U35405(n33537,n33390,n32621);
  nor U35406(n32621,n33392,n33544);
  nand U35407(n33543,n29994,n31450,n32417);
  nand U35408(n29994,n33235,n32778);
  nor U35409(n32778,n33236,n33314);
  nand U35410(G2388,n33545,n33546,n33547,n33548);
  nor U35411(n33548,n33549,n33550,n33551);
  nor U35412(n33551,n33552,n32451);
  not U35413(n32451,n32346);
  nor U35414(n33550,n32342,n33553);
  not U35415(n32342,n32457);
  nand U35416(n32457,n33554,n33555);
  nand U35417(n33555,n33556,n28689);
  nand U35418(n33554,n32346,G58977);
  nor U35419(n32346,n26779,n32332);
  not U35420(n26779,G58871);
  nor U35421(n33549,n29993,n32344);
  nand U35422(n32344,n32417,G58895);
  nand U35423(n33547,n33557,G58887);
  nand U35424(n33546,G58871,n33558);
  nand U35425(n33545,n33559,G58987);
  nand U35426(G2387,n33560,n33561,n33562,n33563);
  nor U35427(n33563,n33564,n33565,n33566);
  nor U35428(n33566,n33552,n32465);
  not U35429(n32465,n32358);
  nor U35430(n33565,n32356,n33553);
  not U35431(n32356,n32467);
  nand U35432(n32467,n33567,n33568);
  nand U35433(n33568,n33556,n27942);
  nand U35434(n33567,n32358,G58977);
  nor U35435(n32358,n26797,n32332);
  not U35436(n26797,G58872);
  nor U35437(n33564,n29993,n32357);
  nand U35438(n32357,n32417,G58896);
  nand U35439(n33562,n33557,G58888);
  nand U35440(n33561,G58872,n33558);
  nand U35441(n33560,n33559,G58986);
  nand U35442(G2386,n33569,n33570,n33571,n33572);
  nor U35443(n33572,n33573,n33574,n33575);
  nor U35444(n33575,n33552,n32475);
  not U35445(n32475,n32368);
  nor U35446(n33574,n32366,n33553);
  not U35447(n32366,n32477);
  nand U35448(n32477,n33576,n33577);
  nand U35449(n33577,n33556,n32006);
  nand U35450(n33576,n32368,G58977);
  nor U35451(n32368,n26814,n32332);
  not U35452(n26814,G58873);
  nor U35453(n33573,n29993,n32367);
  nand U35454(n32367,n32417,G58897);
  nand U35455(n33571,n33557,G58889);
  nand U35456(n33570,G58873,n33558);
  nand U35457(n33569,n33559,G58985);
  nand U35458(G2385,n33578,n33579,n33580,n33581);
  nor U35459(n33581,n33582,n33583,n33584);
  nor U35460(n33584,n33552,n32485);
  not U35461(n32485,n32378);
  nor U35462(n33583,n32376,n33553);
  not U35463(n32376,n32487);
  nand U35464(n32487,n33585,n33586);
  nand U35465(n33586,n33556,n28572);
  nand U35466(n33585,n32378,G58977);
  nor U35467(n32378,n26831,n32332);
  not U35468(n26831,G58874);
  nor U35469(n33582,n29993,n32377);
  nand U35470(n32377,n32417,G58898);
  nand U35471(n33580,n33557,G58890);
  nand U35472(n33579,G58874,n33558);
  nand U35473(n33578,n33559,G58984);
  nand U35474(G2384,n33587,n33588,n33589,n33590);
  nor U35475(n33590,n33591,n33592,n33593);
  nor U35476(n33593,n33552,n32495);
  not U35477(n32495,n32388);
  nor U35478(n33592,n32386,n33553);
  not U35479(n32386,n32497);
  nand U35480(n32497,n33594,n33595);
  nand U35481(n33595,n33556,n32316);
  nand U35482(n33594,n32388,G58977);
  nor U35483(n32388,n26848,n32332);
  not U35484(n26848,G58875);
  nor U35485(n33591,n29993,n32387);
  nand U35486(n32387,n32417,G58899);
  nand U35487(n33589,n33557,G58891);
  nand U35488(n33588,G58875,n33558);
  nand U35489(n33587,n33559,G58983);
  nand U35490(G2383,n33596,n33597,n33598,n33599);
  nor U35491(n33599,n33600,n33601,n33602);
  nor U35492(n33602,n33552,n32505);
  not U35493(n32505,n32398);
  nor U35494(n33601,n32396,n33553);
  not U35495(n32396,n32507);
  nand U35496(n32507,n33603,n33604);
  nand U35497(n33604,n33556,n33605);
  nand U35498(n33603,n32398,G58977);
  nor U35499(n32398,n26866,n32332);
  not U35500(n26866,G58876);
  nor U35501(n33600,n29993,n32397);
  nand U35502(n32397,n32417,G58900);
  nand U35503(n33598,n33557,G58892);
  nand U35504(n33597,G58876,n33558);
  nand U35505(n33596,n33559,G58982);
  nand U35506(G2382,n33606,n33607,n33608,n33609);
  nor U35507(n33609,n33610,n33611,n33612);
  nor U35508(n33612,n33552,n32515);
  not U35509(n32515,n32408);
  nor U35510(n33611,n32406,n33553);
  not U35511(n32406,n32517);
  nand U35512(n32517,n33613,n33614);
  nand U35513(n33614,n33556,n28419);
  nand U35514(n33613,n32408,G58977);
  nor U35515(n32408,n26883,n32332);
  not U35516(n26883,G58877);
  nor U35517(n33610,n29993,n32407);
  nand U35518(n32407,n32417,G58901);
  nand U35519(n33608,n33557,G58893);
  nand U35520(n33607,G58877,n33558);
  nand U35521(n33606,n33559,G58981);
  nand U35522(G2381,n33615,n33616,n33617,n33618);
  nor U35523(n33618,n33619,n33620,n33621);
  nor U35524(n33621,n32418,n33553);
  not U35525(n32418,n32544);
  nand U35526(n32544,n33622,n33623);
  nand U35527(n33623,n33556,n33624);
  nor U35528(n33556,n27932,n32332);
  nand U35529(n33622,n32429,G58977);
  nor U35530(n33620,n33552,n32531);
  not U35531(n32531,n32429);
  nor U35532(n32429,n26913,n32332);
  not U35533(n26913,G58878);
  and U35534(n33552,n33625,n33626);
  nand U35535(n33626,n33627,n29226);
  nand U35536(n33625,n33628,G58977);
  nor U35537(n33619,n29993,n32419);
  nand U35538(n32419,n32417,G58902);
  nand U35539(n33617,n33557,G58894);
  and U35540(n33557,n32417,n33628);
  not U35541(n33628,n31451);
  nand U35542(n33616,G58878,n33558);
  nand U35543(n33558,n33629,n33630);
  nand U35544(n33630,n32417,n29993,n33627);
  not U35545(n33627,n33631);
  nand U35546(n33629,n33632,n33633);
  nand U35547(n33615,n33559,G58980);
  and U35548(n33559,n33634,n33635);
  nand U35549(n33635,n33636,n32423,n33637);
  nand U35550(n33637,G58977,n31451);
  nor U35551(n32423,n32332,n27960);
  nand U35552(n33636,n33633,n33631);
  nand U35553(n33631,n33390,n32697);
  nor U35554(n32697,G59117,n33544);
  nor U35555(n33390,n33005,n33312);
  not U35556(n33005,n32699);
  nand U35557(n33633,n33638,n32434);
  not U35558(n32434,n32530);
  nor U35559(n32530,n29174,n32332);
  nand U35560(n33638,n29993,n31451,n32417);
  nand U35561(n29993,n33235,n32854);
  nor U35562(n32854,n33236,n33237);
  nor U35563(n33235,n33469,n33007);
  nand U35564(n33634,n33632,n32428);
  nand U35565(n32428,n33640,n33641,n33642);
  or U35566(n33642,n27904,n27916);
  nand U35567(n33641,n27931,n33643);
  nand U35568(n33640,n27929,n28416,G58978);
  not U35569(n33632,n33553);
  nand U35570(n33553,n33389,n32701);
  nor U35571(n33389,n33644,n33645);
  nand U35572(G2380,n28440,n33646,n33647,n33648);
  nand U35573(n33648,n33649,G58979);
  nand U35574(n33647,n33650,n33651);
  nand U35575(n33650,n33652,n33653,n33654);
  nand U35576(n33654,n33655,n27965);
  nand U35577(n33653,n33656,n28416);
  nand U35578(n33656,G58976,n27965,n27960);
  nand U35579(n33652,n27870,n33657);
  nand U35580(n28440,G58976,G58979,n27960);
  nand U35581(G2379,n33658,n28439,n33659);
  nand U35582(n33659,G58978,n33660);
  nand U35583(n33660,n33651,n33646);
  nand U35584(n33646,G58979,n27929,n28770);
  nand U35585(n28439,n27929,n28416,n29226);
  nand U35586(n33658,n33661,n33651);
  nand U35587(n33661,n28448,n33662);
  nand U35588(n33662,n27930,n27928,n29176);
  not U35589(n28448,n27907);
  nor U35590(n27907,n28962,n28416);
  nand U35591(G2378,n28962,n32327,n33663,n33664);
  or U35592(n33664,n33639,G58979);
  nand U35593(n33663,n27930,n27929,G58978,G58979);
  nand U35594(G2377,n33665,n27904,n33666);
  nand U35595(n33666,n33649,G58976);
  not U35596(n33649,n33651);
  nand U35597(n33651,n33667,n33668,n33669);
  nand U35598(n33669,n33670,n28416);
  nand U35599(n33670,n28770,G58978);
  nand U35600(n33668,n28961,n27945,n28423);
  nor U35601(n28423,G59348,n28770);
  nand U35602(n33667,n33671,n32327);
  or U35603(n33671,n33657,n28962);
  not U35604(n28962,n27870);
  nor U35605(n27870,n27929,G58978);
  nand U35606(n33657,n33672,n33673,n33674,n33675);
  nor U35607(n33675,n33676,n33677,n33678,n33679);
  and U35608(n33679,n27871,n27872);
  xnor U35609(n27871,n33680,n31650);
  and U35610(n31650,n33681,n33682);
  nand U35611(n33681,n33683,n33684);
  nand U35612(n33680,n31651,n31648);
  nand U35613(n31648,n33685,n33686);
  or U35614(n31651,n33686,n33685);
  nor U35615(n33685,n27999,n30221);
  xor U35616(n33686,n33687,n29226);
  nand U35617(n33687,n33688,n33689,n33690,n33691);
  nor U35618(n33691,n33692,n33693);
  nor U35619(n33693,n29173,n29145);
  nor U35620(n33692,n28963,n31664);
  not U35621(n31664,G59313);
  nand U35622(n33690,G59122,n29287);
  nand U35623(n33689,G59108,n33694);
  nand U35624(n33694,n28769,n33695);
  nand U35625(n33695,n28875,G58979);
  nand U35626(n33688,n28559,n29288);
  not U35627(n28559,n28369);
  xnor U35628(n28369,n31644,n31643);
  xnor U35629(n31644,n27993,n33696);
  nor U35630(n33696,n33697,n33698,n33699,n33700);
  and U35631(n33700,n29228,G59249);
  nor U35632(n33699,n29486,n31514);
  not U35633(n31514,G59122);
  nor U35634(n33698,n29174,n29145);
  not U35635(n29145,G59154);
  nor U35636(n33697,n31034,n28370);
  not U35637(n28370,G59281);
  not U35638(n31034,n29225);
  nor U35639(n33678,n31673,n27908);
  nor U35640(n33677,n32306,n32286);
  nor U35641(n33676,n33701,n33702);
  nor U35642(n33674,n29177,n33703);
  nor U35643(n33703,n33704,n27986);
  nand U35644(n27986,n27976,n33705);
  nand U35645(n33705,n33706,n27930);
  nand U35646(n33706,n33707,n27944,n33708);
  nand U35647(n33708,n28959,n32006);
  and U35648(n27976,n33709,n33710,n33711,n33712);
  nand U35649(n33711,n28691,n33713);
  nand U35650(n33713,n33714,n33715);
  nor U35651(n33709,n33716,n33717);
  nor U35652(n33717,n32311,n27965);
  nor U35653(n33716,n32306,n33707);
  not U35654(n32306,n27990);
  nor U35655(n33704,G59346,G59347);
  nand U35656(n33673,n33718,n32330);
  nand U35657(n33718,n33719,n33720);
  nand U35658(n33720,n33721,n33644,n33722);
  not U35659(n33722,n33702);
  nand U35660(n33719,n33723,n33645);
  nand U35661(n33723,n33702,n33724);
  nand U35662(n33724,n33725,n33721);
  nand U35663(n33721,n33726,n33727,n33728,n33729);
  nand U35664(n33729,n33730,n33731);
  nand U35665(n33731,n33732,n33733);
  nand U35666(n33733,G59111,n33734);
  nand U35667(n33728,n33735,n27898,n27908);
  nand U35668(n27898,n33736,n33737,n33738,n33739);
  nor U35669(n33739,n33740,n33741,n33742);
  nor U35670(n33742,n33743,n33007);
  nor U35671(n33741,n33744,n33745);
  nor U35672(n33744,n31162,n29948);
  not U35673(n29948,n29945);
  nor U35674(n29945,n33746,n31155);
  nor U35675(n33746,n31181,n27943);
  nor U35676(n33740,n32189,n32285);
  nor U35677(n32189,n31155,n31162);
  nand U35678(n33738,n28406,n33747);
  nand U35679(n33737,n27900,n33748);
  not U35680(n27900,n28405);
  xnor U35681(n28405,n33749,n33750);
  and U35682(n33750,n33751,n33752);
  nand U35683(n33736,n27899,n33753);
  or U35684(n33735,n27912,n33734);
  not U35685(n33734,n32701);
  nand U35686(n33727,n33754,n33755);
  nand U35687(n33754,n33756,n33757,G59117);
  nand U35688(n33757,n33730,G59112);
  nand U35689(n33756,n27912,n27908);
  nand U35690(n27912,n33758,n33759,n33760,n33761);
  nor U35691(n33761,n33762,n33763);
  nor U35692(n33763,n33764,n32275);
  not U35693(n32275,n27969);
  nor U35694(n33762,n33765,n27914);
  nand U35695(n33760,n27915,n33748);
  xor U35696(n27915,n33766,n29174);
  nand U35697(n33766,n33767,n33768);
  nand U35698(n33759,n33769,n29944);
  nand U35699(n33758,n33314,n33770);
  or U35700(n33726,n33701,G59115);
  nand U35701(n33725,G59115,n33701);
  nand U35702(n33701,n33771,n33772);
  nand U35703(n33772,n33730,n33773);
  or U35704(n33771,n27889,n33730);
  nand U35705(n27889,n33774,n33775,n33776,n33777);
  nor U35706(n33777,n33778,n33779,n33780);
  nor U35707(n33780,n32285,n32197);
  xor U35708(n32197,n33781,n33732);
  not U35709(n33732,n31154);
  nor U35710(n33779,n33743,n33236);
  nor U35711(n33778,n33765,n33782);
  nand U35712(n33776,n29917,n32148);
  xor U35713(n29917,G59110,n33783);
  nand U35714(n33775,n28395,n33747);
  nand U35715(n33774,n27891,n33748);
  not U35716(n27891,n28393);
  nand U35717(n28393,n33784,n33785);
  nand U35718(n33785,n33786,n33787);
  not U35719(n33786,n33788);
  nand U35720(n33784,n33789,n33752,n33790);
  nand U35721(n33789,n33791,n33787);
  nand U35722(n33702,n33792,n33793);
  nand U35723(n33793,n33730,n31791);
  or U35724(n33792,n27882,n33730);
  not U35725(n33730,n27908);
  nand U35726(n27908,n33794,n33795,n32302);
  and U35727(n32302,n33796,n33797,n33798,n33799);
  nor U35728(n33799,n33800,n33801);
  xnor U35729(n33801,n33715,n33802);
  not U35730(n33800,n33710);
  nor U35731(n33710,n33803,n33804,n32162,n33805);
  and U35732(n33803,n33806,n32006);
  nand U35733(n33806,n33807,n28419,n27943);
  not U35734(n33797,n33808);
  nand U35735(n33796,n28759,n33809);
  nand U35736(n33809,n28959,n32316);
  nand U35737(n33795,n33810,n27930);
  nand U35738(n33810,n33811,n33812);
  nand U35739(n33812,n33813,n27965);
  nand U35740(n33813,n32291,n33814);
  nand U35741(n33814,n27945,n33815);
  nand U35742(n33815,n28447,n32290);
  not U35743(n32290,n28875);
  not U35744(n27945,n27944);
  nand U35745(n27944,n28876,n32159);
  or U35746(n33811,n32286,n27990);
  nand U35747(n27990,n33816,n33817);
  nand U35748(n33817,n33818,n33819,n33820,n33821);
  nand U35749(n33821,n33822,n33823,n33824);
  or U35750(n33824,n33825,n27942);
  nand U35751(n33823,n33826,n33827,n33828);
  not U35752(n33828,n33829);
  not U35753(n33827,n32031);
  nand U35754(n33826,n33830,n33831);
  or U35755(n33822,n33831,n33830);
  nand U35756(n33820,n33825,n27942);
  not U35757(n33818,n33832);
  nand U35758(n33794,n33769,n27965);
  nand U35759(n27882,n33833,n33834,n33835,n33836);
  nor U35760(n33836,n33837,n33838,n33839);
  nor U35761(n33839,n32285,n32188);
  nand U35762(n32188,n33840,n33841,n33842);
  nand U35763(n33842,n33843,n28689);
  or U35764(n33841,n33844,n31791);
  nand U35765(n33840,n33845,n33844);
  nand U35766(n33844,n33781,n31154);
  xnor U35767(n33781,n27943,G59110);
  nand U35768(n33845,n33846,n33847);
  nand U35769(n33847,n27943,n31791);
  nor U35770(n33838,n33764,n29152);
  not U35771(n29152,n28383);
  not U35772(n33764,n33747);
  nand U35773(n33747,n33848,n32295,n33849,n32293);
  nand U35774(n32293,n33850,n32316);
  nor U35775(n33849,n32299,n33851);
  nor U35776(n33851,n28959,n33852);
  nor U35777(n32299,n28761,n32316);
  not U35778(n28761,n29264);
  not U35779(n33848,n32297);
  nand U35780(n32297,n28447,n33853,n33854,n33855);
  nand U35781(n33855,n32031,n27943);
  nand U35782(n33854,n33856,n28689);
  nand U35783(n33856,n33857,n33858);
  nand U35784(n33858,n28573,n33859);
  nand U35785(n33859,n33805,n33860);
  nand U35786(n33860,n33707,n27942);
  nand U35787(n33857,n32162,n33707);
  not U35788(n33707,n32311);
  nor U35789(n32311,n32006,n28959);
  nand U35790(n33853,n32162,n33861);
  nand U35791(n33861,n32281,n33802);
  nor U35792(n33837,n33765,n33862);
  not U35793(n33765,n33753);
  nand U35794(n33753,n33863,n32286);
  nand U35795(n33835,n27881,n33748);
  nand U35796(n33748,n32288,n32289,n32284,n32291);
  not U35797(n32291,n27872);
  not U35798(n32289,n33864);
  xnor U35799(n27881,n33683,n33865);
  and U35800(n33865,n33684,n33682);
  nand U35801(n33682,n33866,n33867,n33868);
  nand U35802(n33868,n28576,G59104);
  nand U35803(n33684,G59104,n33869,n28576);
  nand U35804(n33869,n33866,n33867);
  or U35805(n33867,n33870,n29174);
  nand U35806(n33866,n33870,n29174);
  nand U35807(n33870,n33871,n33872,n33873,n33874);
  nor U35808(n33874,n33875,n33876);
  nor U35809(n33876,n29173,n28379);
  nor U35810(n33875,n28963,n28382);
  not U35811(n28382,G59312);
  nand U35812(n33873,G59109,n33877);
  nand U35813(n33872,n28383,n29288);
  nor U35814(n28383,n33878,n31643);
  nor U35815(n31643,n33879,n33880);
  and U35816(n33878,n33880,n33879);
  xor U35817(n33880,n33881,n28963);
  nand U35818(n33881,n33882,n33883,n33884,n33885);
  nor U35819(n33885,n33886,n33887,n33888,n33889);
  nor U35820(n33889,n29174,n28379);
  not U35821(n28379,G59153);
  and U35822(n33888,n29225,G59280);
  nor U35823(n33887,n33890,n31791);
  nor U35824(n33886,n33469,n33639);
  not U35825(n33469,n32856);
  nor U35826(n33884,n33891,n33892);
  and U35827(n33892,n29228,G59248);
  nor U35828(n33891,n29486,n31663);
  not U35829(n31663,G59121);
  nand U35830(n33883,n27960,G59114);
  nand U35831(n33882,n32329,n27931);
  nand U35832(n33871,G59121,n29287);
  and U35833(n33683,n33787,n33788);
  nand U35834(n33788,n33791,n33893);
  nand U35835(n33893,n33790,n33752);
  nand U35836(n33752,n33894,n33895);
  nand U35837(n33895,n33896,n33897);
  nand U35838(n33790,n33749,n33751);
  nand U35839(n33751,n33896,n33897,n33898);
  not U35840(n33898,n33894);
  nand U35841(n33894,n28963,n32327,n33899,n33900);
  nor U35842(n33900,n33901,n33902,n33903);
  nor U35843(n33903,n28959,n33904);
  nor U35844(n33902,n29857,n27999);
  nand U35845(n33899,n32030,n33905,n33714,G58979);
  and U35846(n32030,n32159,n28689,n33715);
  or U35847(n33897,n33906,n29174);
  nand U35848(n33896,n29174,n33906);
  nand U35849(n33906,n33907,n33908,n33909,n33910);
  nor U35850(n33910,n33911,n33912);
  nor U35851(n33912,n29173,n28404);
  nor U35852(n33911,n28963,n28015);
  not U35853(n28015,G59310);
  nand U35854(n33909,n28406,n29288);
  not U35855(n28406,n29166);
  xor U35856(n29166,n33913,n33914);
  nand U35857(n33913,n33915,n33916);
  nand U35858(n33908,G59119,n29287);
  nand U35859(n33907,G59111,n33877);
  nand U35860(n33749,n33768,n33917);
  nand U35861(n33917,n29226,n33767);
  nand U35862(n33767,n33918,n33919,n33920);
  not U35863(n33920,n33921);
  nand U35864(n33768,n33921,n33922);
  nand U35865(n33922,n33918,n33919);
  or U35866(n33919,n33923,n29174);
  nand U35867(n33918,n33923,n29174);
  nand U35868(n33923,n33924,n33925,n33926,n33927);
  nor U35869(n33927,n33928,n33929);
  nor U35870(n33929,n29173,n28415);
  nor U35871(n33928,n28963,n28013);
  not U35872(n28013,G59309);
  nand U35873(n33926,G59112,n33877);
  nand U35874(n33925,n27969,n29288);
  nand U35875(n27969,n33930,n33931);
  nand U35876(n33931,n33932,n33933);
  nand U35877(n33932,n33934,n33935);
  nand U35878(n33935,n33936,n28963);
  or U35879(n33930,n33933,n28963);
  nand U35880(n33924,G59118,n29287);
  nand U35881(n33921,n33937,n33938,n33939,n27932);
  nand U35882(n33938,G58979,n33940);
  nand U35883(n33940,n33941,n33624,n33942,n33943);
  nor U35884(n33943,n33944,n33945,n33946,n33947);
  nor U35885(n33945,n33948,n33949);
  nor U35886(n33949,n33950,n33951);
  nor U35887(n33951,n28573,n33605);
  nor U35888(n33950,n28959,n27965);
  nor U35889(n33944,n28572,n28419);
  nand U35890(n33942,n28759,n33807);
  not U35891(n33941,n33850);
  nand U35892(n33937,n28576,G59107);
  nand U35893(n33791,n33952,n33953,n33939,n33639);
  xnor U35894(n33952,n29226,n33954);
  nand U35895(n33787,n33955,n33956);
  nand U35896(n33956,n33939,n33639,n33953);
  nand U35897(n33953,n28576,G59105);
  xnor U35898(n33955,n33954,n29174);
  nand U35899(n33954,n33957,n33958,n33959,n33960);
  nand U35900(n33960,G59110,n33877);
  nand U35901(n33877,n28769,n28765,n27932,n33961);
  nor U35902(n33961,n33962,n33963,n33964);
  nor U35903(n33964,n28959,n28416,n32283,n27965);
  not U35904(n32283,n29177);
  nor U35905(n33963,n33965,n28416);
  nor U35906(n33965,n28875,n33864);
  nor U35907(n33864,n33966,n28689);
  nor U35908(n33962,n28416,n32288);
  not U35909(n28765,n29228);
  nor U35910(n33959,n33967,n33968);
  nor U35911(n33968,n29237,n31775);
  not U35912(n29237,n29287);
  and U35913(n33970,n33971,n33972,n33939);
  nand U35914(n33939,G58979,n28419,n32310,n33973);
  and U35915(n33973,n33905,n31324);
  nor U35916(n31324,n27954,n27943);
  nand U35917(n33969,G58979,n32298);
  nand U35918(n32298,n33863,n33974);
  and U35919(n33863,n33975,n33976);
  nand U35920(n33976,n33850,n33977,n33805);
  or U35921(n33975,n33966,n27943);
  and U35922(n33967,n29288,n28395);
  not U35923(n28395,n29159);
  nand U35924(n29159,n33978,n33879);
  nand U35925(n33879,n33979,n33980);
  nand U35926(n33980,n33981,n33915);
  xnor U35927(n33979,n33982,n28963);
  nand U35928(n33978,n33981,n33915,n33983);
  xnor U35929(n33983,n27993,n33982);
  nand U35930(n33982,n33984,n33985,n33986,n33987);
  nor U35931(n33987,n33988,n33989,n33990,n33991);
  nor U35932(n33991,n33782,n32327);
  nor U35933(n33990,n33639,n33236);
  nand U35934(n33236,n33992,n33993);
  nand U35935(n33993,n33994,n33995);
  nand U35936(n33994,n33996,n33997);
  nand U35937(n33992,n33998,n27946);
  xor U35938(n33998,n33999,n34000);
  nor U35939(n33989,n33644,n27932);
  and U35940(n33988,n29228,G59247);
  nor U35941(n33986,n34001,n34002);
  nor U35942(n34002,n29486,n31775);
  not U35943(n31775,G59120);
  nor U35944(n34001,n29174,n28392);
  not U35945(n28392,G59152);
  nand U35946(n33985,G59110,n34003);
  nand U35947(n33984,G59279,n29225);
  nand U35948(n33915,n34004,n34005);
  nand U35949(n34005,n33972,n29174,n27998,n34006);
  and U35950(n34006,n34007,n34008);
  xnor U35951(n34004,n34009,n28963);
  nand U35952(n33981,n33916,n33914);
  nand U35953(n33914,n33933,n34010);
  nand U35954(n34010,n27993,n33934);
  nand U35955(n33934,n34011,n34012);
  not U35956(n34011,n33936);
  nand U35957(n33933,n34013,n33936);
  nand U35958(n33936,n29173,n34014,n27998,n27932);
  nand U35959(n34014,G58979,n34015);
  nand U35960(n34015,n34016,n34017,n34018,n34019);
  nor U35961(n34019,n34020,n34021,n34022);
  nor U35962(n34022,n28573,n34023);
  nor U35963(n34021,n32310,n34024,n34025);
  nor U35964(n34025,n28573,n33715);
  nor U35965(n34024,n33948,n33605);
  nor U35966(n34020,n32006,n32281);
  not U35967(n34018,n33946);
  nand U35968(n33946,n34026,n34027,n34028,n34029);
  nor U35969(n34029,n33808,n33804);
  nand U35970(n34028,n33715,n32006);
  nand U35971(n34027,n28573,n28689);
  nand U35972(n34026,n33714,n27943);
  nand U35973(n34017,n28759,n27942);
  nand U35974(n34016,n33805,n28959);
  not U35975(n29173,n30080);
  xnor U35976(n34013,n34012,n28963);
  nand U35977(n34012,n34030,n34031);
  nor U35978(n34031,n34032,n34033,n34034,n34035);
  nor U35979(n34035,n33639,n33237);
  not U35980(n33237,n33314);
  nor U35981(n33314,n34036,n34037);
  nor U35982(n34037,n27958,n34038);
  and U35983(n34038,G59112,n34039);
  nor U35984(n34034,n29174,n28415);
  not U35985(n28415,G59150);
  and U35986(n34033,n29225,G59277);
  nor U35987(n34032,n33890,n29944);
  nor U35988(n34030,n34040,n34041,n34042,n34043);
  nor U35989(n34043,n32327,n27914);
  nor U35990(n34042,n33392,n27932);
  and U35991(n34041,n29228,G59245);
  nor U35992(n34040,n29486,n32018);
  nand U35993(n33916,n34044,n34007,n34008,n34045);
  not U35994(n28877,n33972);
  not U35995(n34008,n33901);
  nand U35996(n33901,n28769,n34046);
  nand U35997(n34046,G58979,n28419,n34047);
  nand U35998(n34007,n33850,n33977,G58979,n32159);
  xnor U35999(n34044,n27993,n34009);
  nand U36000(n34009,n34048,n34049);
  nor U36001(n34049,n34050,n34051,n34052,n34053);
  nor U36002(n34053,n29174,n28404);
  not U36003(n28404,G59151);
  and U36004(n34052,n29225,G59278);
  nand U36005(n29225,n28963,n34054);
  nand U36006(n34054,n28577,G58979);
  nor U36007(n34051,n33890,n31181);
  not U36008(n33890,n34003);
  nand U36009(n34003,n27998,n33971,n33972,n33904);
  nand U36010(n33904,G58979,n27965,n29177);
  nand U36011(n33972,G58979,n32159,n28961);
  not U36012(n28961,n28447);
  nand U36013(n33971,G58979,n34055);
  nand U36014(n34055,n34056,n34057,n32295,n34058);
  nor U36015(n34058,n34059,n34060,n34061);
  nor U36016(n34061,n27943,n34062);
  nor U36017(n34062,n34063,n34064,n34065);
  nor U36018(n34065,n33605,n33805,n33948);
  nor U36019(n34064,n33715,n28572);
  nor U36020(n34063,n27942,n28760);
  nor U36021(n34060,n34066,n33712);
  not U36022(n33712,n28759);
  nor U36023(n28759,n28689,n32006);
  nor U36024(n34066,n34067,n33714);
  nor U36025(n34067,n33948,n27954);
  nor U36026(n34059,n34068,n34069);
  and U36027(n32295,n34070,n34071,n34072,n34073);
  nor U36028(n34073,n33804,n34074,n33808);
  nor U36029(n33808,n27942,n31941);
  not U36030(n31941,n32161);
  and U36031(n34074,n32006,n34023);
  nor U36032(n33804,n28573,n28691);
  not U36033(n34072,n33947);
  nand U36034(n33947,n34075,n34076);
  nand U36035(n34076,n34077,n33605);
  nand U36036(n34077,n33802,n33798);
  nand U36037(n33798,n32316,n28419);
  not U36038(n33802,n33714);
  nand U36039(n34075,n32316,n28572,n33715);
  nand U36040(n34071,n28760,n28419,n33715);
  nand U36041(n34070,n34078,n34079);
  nand U36042(n34079,n32310,n28573,n34080,n27954);
  nand U36043(n34078,n34081,n33624);
  nand U36044(n34081,n34047,n32310);
  not U36045(n34047,n34080);
  nand U36046(n34057,n34082,n29264);
  nand U36047(n34056,n33850,n32162);
  not U36048(n27998,n29349);
  nor U36049(n29349,n33745,n28416);
  nor U36050(n34050,n33007,n33639);
  not U36051(n33007,n32855);
  xor U36052(n32855,n34083,n34084);
  xnor U36053(n34083,n34036,n34085);
  nor U36054(n34048,n34086,n34087,n34088,n34089);
  nor U36055(n34089,n34090,n32327);
  nor U36056(n34088,n33755,n27932);
  not U36057(n27932,n27960);
  nor U36058(n27960,G58978,G58977);
  and U36059(n34087,n29228,G59246);
  nor U36060(n29228,n32284,n28416);
  nand U36061(n32284,n32160,n27943,n34091);
  nor U36062(n34086,n29486,n32020);
  not U36063(n29486,n29227);
  nand U36064(n29227,n28769,n34092);
  nand U36065(n34092,G58979,n34093);
  nand U36066(n34093,n34094,n34095,n32288,n33966);
  nand U36067(n33966,n28433,n33715,n33805,n34096);
  nor U36068(n34096,n32316,n28691,n28572);
  nand U36069(n32288,n32316,n34097);
  nand U36070(n34097,n34098,n34080);
  nand U36071(n34080,n32160,n34099);
  nor U36072(n32160,n33605,n27942);
  nand U36073(n34098,n34099,n28433);
  nor U36074(n34099,n28689,n33805,n28760);
  nand U36075(n34095,n33977,n32159,n33850);
  nand U36076(n34094,n27916,n29177);
  nor U36077(n29177,n33852,n34100);
  not U36078(n33852,n34082);
  nor U36079(n34082,n32281,n32006,n33948,n33805);
  nand U36080(n28769,n27872,G58979);
  nor U36081(n27872,n28446,n27942);
  nand U36082(n29288,n29174,n27999);
  not U36083(n27999,n28576);
  nand U36084(n33958,G59311,n27993);
  nand U36085(n32286,n33905,n32031,n33714,n28689);
  nor U36086(n33714,n28419,n32316);
  nand U36087(n33957,G59152,n30080);
  nand U36088(n30080,n32327,n33639);
  nand U36089(n33639,G59348,G58978);
  not U36090(n32327,n27931);
  nand U36091(n33834,n32856,n33770);
  not U36092(n33770,n33743);
  nor U36093(n33743,n28875,n28577);
  not U36094(n28577,n33974);
  nand U36095(n33974,n32031,n28689,n34091);
  nor U36096(n34091,n33624,n28760,n32316,n33948);
  not U36097(n28760,n32162);
  nor U36098(n32162,n28572,n32006);
  nor U36099(n28875,n28446,n28959);
  nand U36100(n32856,n34101,n34102);
  nand U36101(n34102,n34103,n34104);
  nand U36102(n34103,n33996,n34105);
  nand U36103(n34105,n33997,n33995);
  nand U36104(n34101,n34106,n34107);
  nand U36105(n34107,n33997,n34108);
  nand U36106(n34108,n27946,n33996);
  or U36107(n33996,n34000,n33999);
  nand U36108(n33997,n33999,n34000);
  nand U36109(n34000,n34109,n34110);
  nand U36110(n34110,G59110,n34039);
  nand U36111(n34109,n27890,n27929);
  nand U36112(n33999,n34111,n34112);
  nand U36113(n34112,n34113,n34114);
  or U36114(n34114,n34084,n34036);
  not U36115(n34113,n34085);
  nand U36116(n34111,n34084,n34036);
  nand U36117(n34036,n34115,n34116);
  nand U36118(n34116,n27958,n34039,G59112);
  nand U36119(n27958,n27943,G58977);
  nand U36120(n34115,n27971,n27929);
  nand U36121(n34084,n34117,n34118);
  nand U36122(n34118,G59111,n34039);
  nand U36123(n34117,n27899,n27929);
  not U36124(n34106,n34104);
  nand U36125(n34104,n34119,n34120);
  nand U36126(n34120,G59109,n34039);
  nand U36127(n34039,n34085,n33995,n34121);
  nand U36128(n34121,G58977,n28689);
  not U36129(n33995,n27946);
  nor U36130(n27946,n27942,n27929);
  nand U36131(n34085,G58977,n34122);
  nand U36132(n34122,n34100,n34123);
  nand U36133(n34123,n33850,n32159);
  nand U36134(n32159,n34124,n34125);
  nand U36135(n34125,G58941,n27982);
  nor U36136(n33850,n28689,n28959);
  not U36137(n34100,n34068);
  nor U36138(n34068,n28573,n27943);
  nand U36139(n34119,n32329,n27929);
  nand U36140(n33833,n32148,n29918);
  nand U36141(n29918,n34126,n34127);
  nand U36142(n34127,n33846,n33773,n33783);
  not U36143(n33846,n34128);
  nand U36144(n34126,n34129,n31791);
  nand U36145(n34129,n34128,n33783);
  nand U36146(n33783,n27943,n31154);
  not U36147(n32148,n33745);
  nand U36148(n33672,n27916,n34130);
  nand U36149(n34130,n28447,n28446,n34131);
  not U36150(n34131,n33769);
  nand U36151(n33769,n32285,n33745);
  nand U36152(n33745,n29264,n34023,n34132);
  nor U36153(n34132,n27954,n32310,n32006);
  not U36154(n27954,n33830);
  nor U36155(n34023,n28419,n33805);
  nand U36156(n32285,n28424,n33905,n32161,n33605);
  nand U36157(n28446,n27943,n33624,n33977);
  nor U36158(n33977,n32281,n28572,n28691,n33948);
  not U36159(n32281,n33807);
  nor U36160(n33807,n32316,n33715);
  nand U36161(n28447,n32310,n28689,n33715,n34133);
  and U36162(n34133,n33905,n28433);
  nor U36163(n28433,n28419,n27942);
  nor U36164(n33905,n28573,n33805,n32006);
  not U36165(n33805,n33624);
  nand U36166(n33624,n34134,n34135,n34136,n34137);
  nor U36167(n34137,n34138,n34139,n34140,n34141);
  nor U36168(n34141,n34142,n29963);
  nor U36169(n34140,n34143,n29961);
  nor U36170(n34139,n34144,n29979);
  nor U36171(n34138,n34145,n29975);
  nor U36172(n34136,n34146,n34147,n34148,n34149);
  nor U36173(n34149,n34150,n29973);
  nor U36174(n34148,n34151,n29347);
  nor U36175(n34147,n34152,n29343);
  nor U36176(n34146,n34153,n29341);
  nor U36177(n34135,n34154,n34155,n34156,n34157);
  nor U36178(n34157,n34158,n29335);
  nor U36179(n34156,n34159,n29331);
  nor U36180(n34155,n34160,n29329);
  nor U36181(n34154,n34161,n29967);
  nor U36182(n34134,n34162,n34163,n34164,n34165);
  nor U36183(n34165,n34166,n29965);
  nor U36184(n34164,n34167,n29977);
  nor U36185(n34163,n34168,n29345);
  nor U36186(n34162,n34169,n29333);
  not U36187(n32310,n32316);
  nand U36188(n32316,n34170,n34171,n34172,n34173);
  nor U36189(n34173,n34174,n34175,n34176,n34177);
  nor U36190(n34177,n34142,n30219);
  not U36191(n30219,G59087);
  nor U36192(n34176,n34143,n30218);
  not U36193(n30218,G59079);
  nor U36194(n34175,n34144,n30229);
  not U36195(n30229,G59071);
  nor U36196(n34174,n34145,n30227);
  not U36197(n30227,G59055);
  nor U36198(n34172,n34178,n34179,n34180,n34181);
  nor U36199(n34181,n34150,n30226);
  not U36200(n30226,G59047);
  nor U36201(n34180,n34151,n29600);
  not U36202(n29600,G59039);
  nor U36203(n34179,n34152,n29598);
  not U36204(n29598,G59023);
  nor U36205(n34178,n34153,n29597);
  not U36206(n29597,G59015);
  nor U36207(n34171,n34182,n34183,n34184,n34185);
  nor U36208(n34185,n34158,n29592);
  not U36209(n29592,G59007);
  nor U36210(n34184,n34159,n29590);
  not U36211(n29590,G58991);
  nor U36212(n34183,n34160,n29589);
  not U36213(n29589,G58983);
  nor U36214(n34182,n34161,n30221);
  not U36215(n30221,G59103);
  nor U36216(n34170,n34186,n34187,n34188,n34189);
  nor U36217(n34189,n34166,n30220);
  not U36218(n30220,G59095);
  nor U36219(n34188,n34167,n30228);
  not U36220(n30228,G59063);
  nor U36221(n34187,n34168,n29599);
  not U36222(n29599,G59031);
  nor U36223(n34186,n34169,n29591);
  not U36224(n29591,G58999);
  not U36225(n27916,n27965);
  nand U36226(n27965,n34190,n34191);
  or U36227(n34191,n34192,n34193);
  nand U36228(n34190,n34194,n34192,n34195,n34196);
  nor U36229(n34196,n34197,n34198);
  nor U36230(n34198,n34199,n33816);
  nand U36231(n33816,n34200,n34201);
  nand U36232(n34201,G59113,n34202);
  nand U36233(n34202,G59108,n34203);
  or U36234(n34200,n34203,G59108);
  nor U36235(n34197,n31673,G59346,n33643);
  not U36236(n31673,G59108);
  nand U36237(n34195,n34204,n34205,n34206,n34207);
  nor U36238(n34207,n34208,n34209);
  nor U36239(n34209,n34199,n33819);
  xnor U36240(n33819,n34203,n34210);
  xnor U36241(n34210,n32330,G59108);
  not U36242(n32330,G59113);
  nand U36243(n34203,n34211,n34212);
  nand U36244(n34212,n34213,n33645);
  nand U36245(n34213,n34214,n31791);
  nand U36246(n34211,G59109,n34215);
  nor U36247(n34208,G59109,n34216);
  nand U36248(n34206,n34217,n33832);
  nand U36249(n33832,n34218,n34219);
  nand U36250(n34219,n34220,n34215);
  xnor U36251(n34220,G59114,G59109);
  nand U36252(n34218,n34221,n34214);
  not U36253(n34214,n34215);
  nand U36254(n34215,n34222,n34223);
  nand U36255(n34223,n34224,n33644);
  nand U36256(n34224,n33773,n34225);
  or U36257(n34222,n34225,n33773);
  xnor U36258(n34221,n33645,G59109);
  nand U36259(n34205,n34226,n34227);
  nand U36260(n34227,n34228,n34229);
  nand U36261(n34229,n34230,n34231);
  nand U36262(n34231,n27928,n34232,G59110);
  nand U36263(n34226,n34216,n34233);
  nand U36264(n34204,n34234,n34235,n34236);
  nand U36265(n34236,n34237,n34238);
  nand U36266(n34238,n34216,n34239);
  not U36267(n34237,n34240);
  nand U36268(n34235,n34233,n34228,n34216);
  nand U36269(n34228,n34217,n33825);
  xor U36270(n33825,n34241,n34225);
  nand U36271(n34225,n34242,n34243);
  nand U36272(n34243,G59116,n34244);
  or U36273(n34244,n34245,n31181);
  nand U36274(n34242,n34245,n31181);
  xnor U36275(n34241,G59115,G59110);
  nand U36276(n34234,n34246,n34247,n34248);
  nand U36277(n34248,n34230,n29944);
  nand U36278(n34247,n34249,n33643);
  nand U36279(n34249,n34250,n34233);
  nand U36280(n34233,n34069,n34251);
  nand U36281(n34251,n33948,n33605);
  nand U36282(n34250,n34239,n34240);
  nand U36283(n34240,n34252,n34253,n34254);
  nand U36284(n34254,n34217,n33831);
  xnor U36285(n33831,n34245,n34255);
  xnor U36286(n34255,n33755,G59111);
  not U36287(n34253,n34256);
  nand U36288(n34252,n34257,n34230);
  nand U36289(n34257,n34258,n34259,n27928);
  not U36290(n27928,G58976);
  nand U36291(n34259,n31181,n34232);
  not U36292(n34232,G59346);
  nand U36293(n34258,G59346,n34260);
  nand U36294(n34260,G59118,n27899);
  nand U36295(n34239,n34261,n34262);
  nand U36296(n34262,n33830,n33948);
  nor U36297(n33830,n27942,n33715);
  not U36298(n34261,n34193);
  nand U36299(n34246,n34217,n33829);
  nand U36300(n33829,n34245,n34263);
  nand U36301(n34263,G59117,n29944);
  nand U36302(n34245,G59112,n33392);
  not U36303(n34217,n34199);
  nand U36304(n34199,n34216,n34264);
  nand U36305(n34264,n34193,n34069);
  not U36306(n34069,n28424);
  nor U36307(n28424,n28419,n28959);
  nor U36308(n34193,n28573,n28959,n33715);
  not U36309(n33715,n33605);
  nand U36310(n34192,n34256,n31325);
  nand U36311(n31325,n34265,n34266,n34267,n34268);
  nor U36312(n34268,n34269,n34270,n34271,n34272);
  nor U36313(n34272,n29963,n31433);
  nand U36314(n31433,n34273,n34274);
  not U36315(n29963,G59084);
  nor U36316(n34271,n29961,n31434);
  nand U36317(n31434,n34273,n34275);
  not U36318(n29961,G59076);
  nor U36319(n34270,n29979,n31435);
  nand U36320(n31435,n34276,n34277);
  not U36321(n29979,G59068);
  nor U36322(n34269,n29975,n31436);
  nand U36323(n31436,n34277,n34274);
  not U36324(n29975,G59052);
  nor U36325(n34267,n34278,n34279,n34280,n34281);
  nor U36326(n34281,n29973,n31441);
  nand U36327(n31441,n34275,n34277);
  not U36328(n29973,G59044);
  nor U36329(n34280,n29347,n31442);
  nand U36330(n31442,n34282,n34276);
  not U36331(n29347,G59036);
  nor U36332(n34279,n29343,n31443);
  nand U36333(n31443,n34282,n34274);
  not U36334(n29343,G59020);
  nor U36335(n34278,n29341,n31444);
  nand U36336(n31444,n34282,n34275);
  not U36337(n29341,G59012);
  nor U36338(n34266,n34283,n34284,n34285,n34286);
  nor U36339(n34286,n29335,n31449);
  nand U36340(n31449,n34287,n34276);
  not U36341(n29335,G59004);
  nor U36342(n34285,n29331,n31450);
  nand U36343(n31450,n34287,n34274);
  nor U36344(n34274,n34090,n27971);
  not U36345(n29331,G58988);
  nor U36346(n34284,n29329,n31451);
  nand U36347(n31451,n34287,n34275);
  nor U36348(n34275,n27914,n34090);
  not U36349(n34090,n27899);
  not U36350(n29329,G58980);
  nor U36351(n34283,n29967,n31452);
  nand U36352(n31452,n34273,n34276);
  nor U36353(n34276,n27899,n27971);
  not U36354(n27971,n27914);
  not U36355(n29967,G59100);
  nor U36356(n34265,n34288,n34289,n34290,n34291);
  nor U36357(n34291,n29965,n31457);
  nand U36358(n31457,n34292,n34273);
  nor U36359(n34273,n27890,n32329);
  not U36360(n29965,G59092);
  nor U36361(n34290,n29977,n31458);
  nand U36362(n31458,n34292,n34277);
  nor U36363(n34277,n33782,n32329);
  not U36364(n32329,n33862);
  not U36365(n29977,G59060);
  nor U36366(n34289,n29345,n31459);
  nand U36367(n31459,n34292,n34282);
  nor U36368(n34282,n33862,n27890);
  not U36369(n29345,G59028);
  nor U36370(n34288,n29333,n31460);
  nand U36371(n31460,n34292,n34287);
  nor U36372(n34287,n33862,n33782);
  not U36373(n33782,n27890);
  xor U36374(n27890,n34293,n34294);
  xnor U36375(n33862,n34295,n34296);
  nor U36376(n34296,n34293,n34294);
  and U36377(n34294,n34297,n34298);
  nand U36378(n34298,n34299,n34300);
  or U36379(n34300,n34301,n34302);
  not U36380(n34299,n34303);
  nand U36381(n34297,n34302,n34301);
  and U36382(n34293,n34304,n34305,n34306);
  nand U36383(n34306,G59115,n27931);
  nand U36384(n34305,n32699,n27929);
  xnor U36385(n32699,n32701,n33644);
  nand U36386(n34304,n29176,G59110);
  nand U36387(n34295,n34307,n34308,n34309);
  nand U36388(n34309,n27929,n32698);
  not U36389(n32698,n33312);
  nor U36390(n33312,n32999,n33082,n34310);
  nor U36391(n34310,n33645,n32701);
  nor U36392(n33082,n33645,G59115);
  not U36393(n33645,G59114);
  not U36394(n32999,n32939);
  nand U36395(n32939,n32701,n32776);
  nor U36396(n32776,n33644,G59114);
  not U36397(n33644,G59115);
  nor U36398(n32701,n33392,n33755);
  nand U36399(n34308,G59114,n27931);
  nand U36400(n34307,n29176,G59109);
  nor U36401(n34292,n27914,n27899);
  xor U36402(n27899,n34311,n34302);
  nand U36403(n34302,n34312,n34313);
  nand U36404(n34313,n33655,n34314);
  xnor U36405(n34314,n32020,n34315);
  nor U36406(n34315,n28429,n32018);
  nand U36407(n28429,n34316,n34317);
  nand U36408(n34317,G58978,n29188);
  not U36409(n29188,G59149);
  or U36410(n34316,G58978,G59308);
  not U36411(n32020,G59119);
  nand U36412(n34312,n32031,n29176);
  xnor U36413(n34311,n34303,n34301);
  nand U36414(n34301,n34318,n34319,n34320);
  nand U36415(n34320,G59116,n27931);
  nand U36416(n34319,n33391,n27929);
  not U36417(n33391,n33544);
  nor U36418(n33544,n32620,n32545);
  nor U36419(n32545,n33392,G59116);
  nor U36420(n32620,n33755,G59117);
  not U36421(n33755,G59116);
  nand U36422(n34318,n29176,G59111);
  nand U36423(n27914,n34321,n34303);
  nand U36424(n34303,n34322,n34323);
  or U36425(n34321,n34323,n34322);
  nand U36426(n34322,n34324,n34325,G58977);
  nand U36427(n34325,n33643,n27955);
  nand U36428(n27955,n28691,n28689,n32031);
  nor U36429(n32031,n33605,n28959);
  not U36430(n28959,n27942);
  nand U36431(n27942,n34326,n34327,n34328,n34329);
  nor U36432(n34329,n34330,n34331,n34332,n34333);
  nor U36433(n34333,n34142,n29855);
  not U36434(n29855,G59090);
  nor U36435(n34332,n34143,n29854);
  not U36436(n29854,G59082);
  nor U36437(n34331,n34144,n29849);
  not U36438(n29849,G59074);
  nor U36439(n34330,n34145,n29847);
  not U36440(n29847,G59058);
  nor U36441(n34328,n34334,n34335,n34336,n34337);
  nor U36442(n34337,n34150,n29846);
  not U36443(n29846,G59050);
  nor U36444(n34336,n34151,n29841);
  not U36445(n29841,G59042);
  nor U36446(n34335,n34152,n29839);
  not U36447(n29839,G59026);
  nor U36448(n34334,n34153,n29838);
  not U36449(n29838,G59018);
  nor U36450(n34327,n34338,n34339,n34340,n34341);
  nor U36451(n34341,n34158,n29833);
  not U36452(n29833,G59010);
  nor U36453(n34340,n34159,n29831);
  not U36454(n29831,G58994);
  nor U36455(n34339,n34160,n29830);
  not U36456(n29830,G58986);
  nor U36457(n34338,n34161,n29857);
  not U36458(n29857,G59106);
  nor U36459(n34326,n34342,n34343,n34344,n34345);
  nor U36460(n34345,n34166,n29856);
  not U36461(n29856,G59098);
  nor U36462(n34344,n34167,n29848);
  not U36463(n29848,G59066);
  nor U36464(n34343,n34168,n29840);
  not U36465(n29840,G59034);
  nor U36466(n34342,n34169,n29832);
  not U36467(n29832,G59002);
  nand U36468(n33605,n34346,n34347,n34348,n34349);
  nor U36469(n34349,n34350,n34351,n34352,n34353);
  nor U36470(n34353,n34142,n30138);
  not U36471(n30138,G59086);
  nor U36472(n34352,n34143,n30137);
  not U36473(n30137,G59078);
  nor U36474(n34351,n34144,n30148);
  not U36475(n30148,G59070);
  nor U36476(n34350,n34145,n30146);
  not U36477(n30146,G59054);
  nor U36478(n34348,n34354,n34355,n34356,n34357);
  nor U36479(n34357,n34150,n30145);
  not U36480(n30145,G59046);
  nor U36481(n34356,n34151,n29521);
  not U36482(n29521,G59038);
  nor U36483(n34355,n34152,n29519);
  not U36484(n29519,G59022);
  nor U36485(n34354,n34153,n29518);
  not U36486(n29518,G59014);
  nor U36487(n34347,n34358,n34359,n34360,n34361);
  nor U36488(n34361,n34158,n29513);
  not U36489(n29513,G59006);
  nor U36490(n34360,n34159,n29511);
  not U36491(n29511,G58990);
  nor U36492(n34359,n34160,n29510);
  not U36493(n29510,G58982);
  nor U36494(n34358,n34161,n30140);
  not U36495(n30140,G59102);
  nor U36496(n34346,n34362,n34363,n34364,n34365);
  nor U36497(n34365,n34166,n30139);
  not U36498(n30139,G59094);
  nor U36499(n34364,n34167,n30147);
  not U36500(n30147,G59062);
  nor U36501(n34363,n34168,n29520);
  not U36502(n29520,G59030);
  nor U36503(n34362,n34169,n29512);
  not U36504(n29512,G58998);
  nor U36505(n34369,n34370,n34371,n34372,n34373);
  nor U36506(n34373,n34142,n29946);
  not U36507(n29946,G59091);
  nor U36508(n34372,n34143,n29942);
  not U36509(n29942,G59083);
  nor U36510(n34371,n34144,n29937);
  not U36511(n29937,G59075);
  nor U36512(n34370,n34145,n29935);
  not U36513(n29935,G59059);
  nor U36514(n34368,n34374,n34375,n34376,n34377);
  nor U36515(n34377,n34150,n29933);
  not U36516(n29933,G59051);
  nor U36517(n34376,n34151,n29927);
  not U36518(n29927,G59043);
  nor U36519(n34375,n34152,n29925);
  not U36520(n29925,G59027);
  nor U36521(n34374,n34153,n29923);
  not U36522(n29923,G59019);
  nor U36523(n34367,n34378,n34379,n34380,n34381);
  nor U36524(n34381,n34158,n29915);
  not U36525(n29915,G59011);
  nor U36526(n34380,n34159,n29911);
  not U36527(n29911,G58995);
  nor U36528(n34379,n34160,n29908);
  not U36529(n29908,G58987);
  nor U36530(n34378,n34161,n29949);
  not U36531(n29949,G59107);
  nor U36532(n34366,n34382,n34383,n34384,n34385);
  nor U36533(n34385,n34166,n29947);
  not U36534(n29947,G59099);
  nor U36535(n34384,n34167,n29936);
  not U36536(n29936,G59067);
  nor U36537(n34383,n34168,n29926);
  not U36538(n29926,G59035);
  nor U36539(n34382,n34169,n29913);
  not U36540(n29913,G59003);
  not U36541(n28691,n32006);
  nand U36542(n32006,n34386,n34387,n34388,n34389);
  nor U36543(n34389,n34390,n34391,n34392,n34393);
  nor U36544(n34393,n34142,n29759);
  not U36545(n29759,G59089);
  nor U36546(n34392,n34143,n29758);
  not U36547(n29758,G59081);
  nor U36548(n34391,n34144,n29753);
  not U36549(n29753,G59073);
  nor U36550(n34390,n34145,n29751);
  not U36551(n29751,G59057);
  nor U36552(n34388,n34394,n34395,n34396,n34397);
  nor U36553(n34397,n34150,n29750);
  not U36554(n29750,G59049);
  nor U36555(n34396,n34151,n29745);
  not U36556(n29745,G59041);
  nor U36557(n34395,n34152,n29743);
  not U36558(n29743,G59025);
  nor U36559(n34394,n34153,n29742);
  not U36560(n29742,G59017);
  nor U36561(n34387,n34398,n34399,n34400,n34401);
  nor U36562(n34401,n34158,n29737);
  not U36563(n29737,G59009);
  nor U36564(n34400,n34159,n29735);
  not U36565(n29735,G58993);
  nor U36566(n34399,n34160,n29734);
  not U36567(n29734,G58985);
  nor U36568(n34398,n34161,n29761);
  not U36569(n29761,G59105);
  nor U36570(n34386,n34402,n34403,n34404,n34405);
  nor U36571(n34405,n34166,n29760);
  not U36572(n29760,G59097);
  nor U36573(n34404,n34167,n29752);
  not U36574(n29752,G59065);
  nor U36575(n34403,n34168,n29744);
  not U36576(n29744,G59033);
  nor U36577(n34402,n34169,n29736);
  not U36578(n29736,G59001);
  nand U36579(n34324,n28445,n34406);
  nand U36580(n34406,G58979,n32018);
  not U36581(n32018,G59118);
  not U36582(n28445,n29176);
  nand U36583(n34323,n29175,n34407,n34408,n34409);
  nand U36584(n34409,n27929,n33392);
  not U36585(n33392,G59117);
  nand U36586(n34408,G59117,n27931);
  nor U36587(n27931,n27929,G58979);
  nand U36588(n34407,n29176,G59112);
  nor U36589(n29176,n28416,G58978);
  not U36590(n29333,G58996);
  nor U36591(n34256,n28573,n33948,n34230);
  not U36592(n34230,n34216);
  nor U36593(n34216,G58978,G58976);
  not U36594(n33948,n28419);
  nand U36595(n28419,n34410,n34411,n34412,n34413);
  nor U36596(n34413,n34414,n34415,n34416,n34417);
  nor U36597(n34417,n34142,n29436);
  not U36598(n29436,G59085);
  nor U36599(n34416,n34143,n29434);
  not U36600(n29434,G59077);
  nor U36601(n34415,n34144,n29428);
  not U36602(n29428,G59069);
  nor U36603(n34414,n34145,n29424);
  not U36604(n29424,G59053);
  nor U36605(n34412,n34418,n34419,n34420,n34421);
  nor U36606(n34421,n34150,n29422);
  not U36607(n29422,G59045);
  nor U36608(n34420,n34151,n29417);
  not U36609(n29417,G59037);
  nor U36610(n34419,n34152,n29415);
  not U36611(n29415,G59021);
  nor U36612(n34418,n34153,n29414);
  not U36613(n29414,G59013);
  nor U36614(n34411,n34422,n34423,n34424,n34425);
  nor U36615(n34425,n34158,n29409);
  not U36616(n29409,G59005);
  nor U36617(n34424,n34159,n29407);
  not U36618(n29407,G58989);
  nor U36619(n34423,n34160,n29406);
  not U36620(n29406,G58981);
  nor U36621(n34422,n34161,n29440);
  not U36622(n29440,G59101);
  nor U36623(n34410,n34426,n34427,n34428,n34429);
  nor U36624(n34429,n34166,n29438);
  not U36625(n29438,G59093);
  nor U36626(n34428,n34167,n29426);
  not U36627(n29426,G59061);
  nor U36628(n34427,n34168,n29416);
  not U36629(n29416,G59029);
  nor U36630(n34426,n34169,n29408);
  not U36631(n29408,G58997);
  not U36632(n28573,n28572);
  nand U36633(n28572,n34430,n34431,n34432,n34433);
  nor U36634(n34433,n34434,n34435,n34436,n34437);
  nor U36635(n34437,n34142,n30303);
  not U36636(n30303,G59088);
  nand U36637(n34142,n34128,n31155);
  nor U36638(n34436,n34143,n30302);
  not U36639(n30302,G59080);
  nand U36640(n34143,n31154,n34128);
  nor U36641(n34435,n34144,n30313);
  not U36642(n30313,G59072);
  nand U36643(n34144,n31163,n31182);
  nor U36644(n34434,n34145,n30311);
  not U36645(n30311,G59056);
  nand U36646(n34145,n31182,n31155);
  nor U36647(n34432,n34438,n34439,n34440,n34441);
  nor U36648(n34441,n34150,n30310);
  not U36649(n30310,G59048);
  nand U36650(n34150,n31154,n31182);
  nor U36651(n34440,n34151,n29676);
  not U36652(n29676,G59040);
  nand U36653(n34151,n31180,n31163);
  nor U36654(n34439,n34152,n29674);
  not U36655(n29674,G59024);
  nand U36656(n34152,n31180,n31155);
  nor U36657(n34438,n34153,n29673);
  not U36658(n29673,G59016);
  nand U36659(n34153,n31180,n31154);
  nor U36660(n34431,n34442,n34443,n34444,n34445);
  nor U36661(n34445,n34158,n29668);
  not U36662(n29668,G59008);
  nand U36663(n34158,n33843,n31163);
  nor U36664(n34444,n34159,n29666);
  not U36665(n29666,G58992);
  nand U36666(n34159,n33843,n31155);
  nor U36667(n31155,n31181,G59112);
  nor U36668(n34443,n34160,n29665);
  not U36669(n29665,G58984);
  nand U36670(n34160,n33843,n31154);
  nor U36671(n31154,n29944,n31181);
  not U36672(n31181,G59111);
  nor U36673(n34442,n34161,n30305);
  not U36674(n30305,G59104);
  nand U36675(n34161,n34128,n31163);
  nor U36676(n31163,G59111,G59112);
  nor U36677(n34430,n34446,n34447,n34448,n34449);
  nor U36678(n34449,n34166,n30304);
  not U36679(n30304,G59096);
  nand U36680(n34166,n31162,n34128);
  nor U36681(n34128,G59110,G59109);
  nor U36682(n34448,n34167,n30312);
  not U36683(n30312,G59064);
  nand U36684(n34167,n31162,n31182);
  nor U36685(n31182,n33773,G59109);
  nor U36686(n34447,n34168,n29675);
  not U36687(n29675,G59032);
  nand U36688(n34168,n31162,n31180);
  nor U36689(n31180,n31791,G59110);
  nor U36690(n34446,n34169,n29667);
  not U36691(n29667,G59000);
  nand U36692(n34169,n31162,n33843);
  nor U36693(n33843,n31791,n33773);
  not U36694(n33773,G59110);
  not U36695(n31791,G59109);
  nor U36696(n31162,n29944,G59111);
  not U36697(n29944,G59112);
  nand U36698(n34194,G59108,G58976);
  nand U36699(n27904,G58976,n28416);
  not U36700(n33665,n32333);
  nor U36701(n32333,n28416,n29175);
  not U36702(n29175,n33655);
  nor U36703(n33655,n33643,n27929);
  not U36704(n27929,G58977);
  not U36705(n33643,G58978);
  not U36706(n28416,G58979);
  nor U36707(G2376,n27862,n28043);
  not U36708(n28043,G58975);
  nor U36709(G2375,n27862,n28042);
  not U36710(n28042,G58974);
  nor U36711(G2374,n27862,n28041);
  not U36712(n28041,G58973);
  nor U36713(G2373,n27862,n28040);
  not U36714(n28040,G58972);
  nor U36715(G2372,n27862,n28039);
  not U36716(n28039,G58971);
  nor U36717(G2371,n27862,n28038);
  not U36718(n28038,G58970);
  nor U36719(G2370,n27862,n28037);
  not U36720(n28037,G58969);
  nor U36721(G2369,n27862,n28036);
  not U36722(n28036,G58968);
  nor U36723(G2368,n27862,n28035);
  not U36724(n28035,G58967);
  nor U36725(G2367,n27862,n28034);
  not U36726(n28034,G58966);
  nor U36727(G2366,n27862,n28033);
  not U36728(n28033,G58965);
  nor U36729(G2365,n27862,n28032);
  not U36730(n28032,G58964);
  nor U36731(G2364,n27862,n28031);
  not U36732(n28031,G58963);
  nor U36733(G2363,n27862,n28030);
  not U36734(n28030,G58962);
  nor U36735(G2362,n27862,n28029);
  not U36736(n28029,G58961);
  nor U36737(G2361,n27862,n28028);
  not U36738(n28028,G58960);
  and U36739(G2360,n27863,G58959);
  and U36740(G2359,n27863,G58958);
  and U36741(G2358,n27863,G58957);
  and U36742(G2357,n27863,G58956);
  and U36743(G2356,n27863,G58955);
  and U36744(G2355,n27863,G58954);
  and U36745(G2354,n27863,G58953);
  and U36746(G2353,n27863,G58952);
  nor U36747(G2352,n27862,n28049);
  not U36748(n28049,G58951);
  nor U36749(G2351,n27862,n28048);
  not U36750(n28048,G58950);
  nor U36751(G2350,n27862,n28047);
  not U36752(n28047,G58949);
  nor U36753(G2349,n27862,n28046);
  not U36754(n28046,G58948);
  and U36755(G2348,n27863,G58947);
  and U36756(G2347,n27863,G58946);
  not U36757(n27863,n27862);
  nand U36758(n27862,n34450,n34451);
  nand U36759(n34451,G58943,n34452);
  nand U36760(G2346,n34453,n34454,n34455,n34456);
  nor U36761(n34456,n34457,n27867,n34458);
  nor U36762(n34458,n34124,n27930);
  not U36763(n34124,n34452);
  nor U36764(n27867,G58943,G58941);
  nor U36765(n34457,n27739,n34450);
  nand U36766(n34455,n27851,n27922);
  nand U36767(n34454,n34459,n27982);
  nand U36768(n34453,G58943,G33,G58942);
  nand U36769(G2345,n34460,n34461,n34462,n34463);
  nand U36770(n34463,n34452,G33);
  nor U36771(n34452,n27982,G58941);
  nor U36772(n34462,n34464,n34465);
  nor U36773(n34465,n27922,n34459,n28876);
  nor U36774(n34459,n34466,n27747);
  or U36775(n34461,n34450,n34466);
  nand U36776(n34450,n27982,n28876);
  nand U36777(n34460,n28770,G58942);
  nand U36778(G2344,n34467,n34468,n34469,n34470);
  nand U36779(n34470,G58941,n27739,n28876);
  not U36780(n28876,G58943);
  nand U36781(n34469,G33,n34471,G58943);
  nand U36782(n34471,n34466,n34472);
  nand U36783(n34472,n27982,n27922);
  not U36784(n34468,n34473);
  nand U36785(n34467,G58942,n34474,n28770);
  not U36786(n28770,n27930);
  nand U36787(n27930,G58905,G37);
  nand U36788(n34474,n34466,n34475);
  nand U36789(n34475,n34476,n27739,G58943);
  nand U36790(n34476,n27922,n27747);
  not U36791(n27922,G59349);
  nand U36792(G2343,n34477,n34478,n34479);
  nand U36793(n34479,G58940,n27851);
  nand U36794(n34478,n34473,G59310);
  nand U36795(n34477,n34464,G59311);
  nand U36796(G2342,n34480,n34481,n34482);
  nand U36797(n34482,G58939,n27851);
  nand U36798(n34481,n34473,G59311);
  nand U36799(n34480,n34464,G59312);
  nand U36800(G2341,n34483,n34484,n34485);
  nand U36801(n34485,G58938,n27851);
  nand U36802(n34484,n34473,G59312);
  nand U36803(n34483,n34464,G59313);
  nand U36804(G2340,n34486,n34487,n34488);
  nand U36805(n34488,G58937,n27851);
  nand U36806(n34487,n34473,G59313);
  nand U36807(n34486,n34464,G59314);
  nand U36808(G2339,n34489,n34490,n34491);
  nand U36809(n34491,G58936,n27851);
  nand U36810(n34490,n34473,G59314);
  nand U36811(n34489,n34464,G59315);
  nand U36812(G2338,n34492,n34493,n34494);
  nand U36813(n34494,G58935,n27851);
  nand U36814(n34493,n34473,G59315);
  nand U36815(n34492,n34464,G59316);
  nand U36816(G2337,n34495,n34496,n34497);
  nand U36817(n34497,G58934,n27851);
  nand U36818(n34496,n34473,G59316);
  nand U36819(n34495,n34464,G59317);
  nand U36820(G2336,n34498,n34499,n34500);
  nand U36821(n34500,G58933,n27851);
  nand U36822(n34499,n34473,G59317);
  nand U36823(n34498,n34464,G59318);
  nand U36824(G2335,n34501,n34502,n34503);
  nand U36825(n34503,G58932,n27851);
  nand U36826(n34502,n34473,G59318);
  nand U36827(n34501,n34464,G59319);
  nand U36828(G2334,n34504,n34505,n34506);
  nand U36829(n34506,G58931,n27851);
  nand U36830(n34505,n34473,G59319);
  nand U36831(n34504,n34464,G59320);
  nand U36832(G2333,n34507,n34508,n34509);
  nand U36833(n34509,G58930,n27851);
  nand U36834(n34508,n34473,G59320);
  nand U36835(n34507,n34464,G59321);
  nand U36836(G2332,n34510,n34511,n34512);
  nand U36837(n34512,G58929,n27851);
  nand U36838(n34511,n34473,G59321);
  nand U36839(n34510,n34464,G59322);
  nand U36840(G2331,n34513,n34514,n34515);
  nand U36841(n34515,G58928,n27851);
  nand U36842(n34514,n34473,G59322);
  nand U36843(n34513,n34464,G59323);
  nand U36844(G2330,n34516,n34517,n34518);
  nand U36845(n34518,G58927,n27851);
  nand U36846(n34517,n34473,G59323);
  nand U36847(n34516,n34464,G59324);
  nand U36848(G2329,n34519,n34520,n34521);
  nand U36849(n34521,G58926,n27851);
  nand U36850(n34520,n34473,G59324);
  nand U36851(n34519,n34464,G59325);
  nand U36852(G2328,n34522,n34523,n34524);
  nand U36853(n34524,G58925,n27851);
  nand U36854(n34523,n34473,G59325);
  nand U36855(n34522,n34464,G59326);
  nand U36856(G2327,n34525,n34526,n34527);
  nand U36857(n34527,G58924,n27851);
  nand U36858(n34526,n34473,G59326);
  nand U36859(n34525,n34464,G59327);
  nand U36860(G2326,n34528,n34529,n34530);
  nand U36861(n34530,G58923,n27851);
  nand U36862(n34529,n34473,G59327);
  nand U36863(n34528,n34464,G59328);
  nand U36864(G2325,n34531,n34532,n34533);
  nand U36865(n34533,G58922,n27851);
  nand U36866(n34532,n34473,G59328);
  nand U36867(n34531,n34464,G59329);
  nand U36868(G2324,n34534,n34535,n34536);
  nand U36869(n34536,G58921,n27851);
  nand U36870(n34535,n34473,G59329);
  nand U36871(n34534,n34464,G59330);
  nand U36872(G2323,n34537,n34538,n34539);
  nand U36873(n34539,G58920,n27851);
  nand U36874(n34538,n34473,G59330);
  nand U36875(n34537,n34464,G59331);
  nand U36876(G2322,n34540,n34541,n34542);
  nand U36877(n34542,G58919,n27851);
  nand U36878(n34541,n34473,G59331);
  nand U36879(n34540,n34464,G59332);
  nand U36880(G2321,n34543,n34544,n34545);
  nand U36881(n34545,G58918,n27851);
  nand U36882(n34544,n34473,G59332);
  nand U36883(n34543,n34464,G59333);
  nand U36884(G2320,n34546,n34547,n34548);
  nand U36885(n34548,G58917,n27851);
  nand U36886(n34547,n34473,G59333);
  nand U36887(n34546,n34464,G59334);
  nand U36888(G2319,n34549,n34550,n34551);
  nand U36889(n34551,G58916,n27851);
  nand U36890(n34550,n34473,G59334);
  nand U36891(n34549,n34464,G59335);
  nand U36892(G2318,n34552,n34553,n34554);
  nand U36893(n34554,G58915,n27851);
  nand U36894(n34553,n34473,G59335);
  nand U36895(n34552,n34464,G59336);
  nand U36896(G2317,n34555,n34556,n34557);
  nand U36897(n34557,G58914,n27851);
  nand U36898(n34556,n34473,G59336);
  nand U36899(n34555,n34464,G59337);
  nand U36900(G2316,n34558,n34559,n34560);
  nand U36901(n34560,G58913,n27851);
  nand U36902(n34559,n34473,G59337);
  nand U36903(n34558,n34464,G59338);
  nand U36904(G2315,n34561,n34562,n34563);
  nand U36905(n34563,G58912,n27851);
  nand U36906(n34562,n34473,G59338);
  nand U36907(n34561,n34464,G59339);
  nand U36908(G2314,n34564,n34565,n34566);
  nand U36909(n34566,G58911,n27851);
  nand U36910(n34565,n34473,G59339);
  not U36911(n34466,G58941);
  nand U36912(n34564,n34464,G59340);
  nor U36913(n27852,n27982,G58943);
  not U36914(n27982,G58942);
  nand U36915(G1721,n34567,n34568);
  nand U36916(n34568,G59389,n34569);
  nand U36917(n34567,n34570,G58940);
  nand U36918(G1720,n34571,n34572);
  nand U36919(n34572,G59379,n34569);
  nand U36920(n34571,n34570,G58930);
  nand U36921(G1719,n34573,n34574);
  nand U36922(n34574,G59378,n34569);
  nand U36923(n34573,n34570,G58929);
  nand U36924(G1718,n34575,n34576);
  nand U36925(n34576,G59377,n34569);
  nand U36926(n34575,n34570,G58928);
  nand U36927(G1717,n34577,n34578);
  nand U36928(n34578,G59376,n34569);
  nand U36929(n34577,n34570,G58927);
  nand U36930(G1716,n34579,n34580);
  nand U36931(n34580,G59375,n34569);
  nand U36932(n34579,n34570,G58926);
  nand U36933(G1715,n34581,n34582);
  nand U36934(n34582,G59374,n34569);
  nand U36935(n34581,n34570,G58925);
  nand U36936(G1714,n34583,n34584);
  nand U36937(n34584,G59373,n34569);
  nand U36938(n34583,n34570,G58924);
  nand U36939(G1713,n34585,n34586);
  nand U36940(n34586,G59372,n34569);
  nand U36941(n34585,n34570,G58923);
  nand U36942(G1712,n34587,n34588);
  nand U36943(n34588,G59371,n34569);
  nand U36944(n34587,n34570,G58922);
  nand U36945(G1711,n34589,n34590);
  nand U36946(n34590,G59370,n34569);
  nand U36947(n34589,n34570,G58921);
  nand U36948(G1710,n34591,n34592);
  nand U36949(n34592,G59388,n34569);
  nand U36950(n34591,n34570,G58939);
  nand U36951(G1709,n34593,n34594);
  nand U36952(n34594,G59369,n34569);
  nand U36953(n34593,n34570,G58920);
  nand U36954(G1708,n34595,n34596);
  nand U36955(n34596,G59368,n34569);
  nand U36956(n34595,n34570,G58919);
  nand U36957(G1707,n34597,n34598);
  nand U36958(n34598,G59367,n34569);
  nand U36959(n34597,n34570,G58918);
  nand U36960(G1706,n34599,n34600);
  nand U36961(n34600,G59366,n34569);
  nand U36962(n34599,n34570,G58917);
  nand U36963(G1705,n34601,n34602);
  nand U36964(n34602,G59365,n34569);
  nand U36965(n34601,n34570,G58916);
  nand U36966(G1704,n34603,n34604);
  nand U36967(n34604,G59364,n34569);
  nand U36968(n34603,n34570,G58915);
  nand U36969(G1703,n34605,n34606);
  nand U36970(n34606,G59363,n34569);
  nand U36971(n34605,n34570,G58914);
  nand U36972(G1702,n34607,n34608);
  nand U36973(n34608,G59362,n34569);
  nand U36974(n34607,n34570,G58913);
  nand U36975(G1701,n34609,n34610);
  nand U36976(n34610,G59361,n34569);
  nand U36977(n34609,n34570,G58912);
  nand U36978(G1700,n34611,n34612);
  nand U36979(n34612,G59360,n34569);
  nand U36980(n34611,n34570,G58911);
  nand U36981(G1699,n34613,n34614);
  nand U36982(n34614,G59387,n34569);
  nand U36983(n34613,n34570,G58938);
  nand U36984(G1698,n34615,n34616);
  nand U36985(n34616,G59386,n34569);
  nand U36986(n34615,n34570,G58937);
  nand U36987(G1697,n34617,n34618);
  nand U36988(n34618,G59385,n34569);
  nand U36989(n34617,n34570,G58936);
  nand U36990(G1696,n34619,n34620);
  nand U36991(n34620,G59384,n34569);
  nand U36992(n34619,n34570,G58935);
  nand U36993(G1695,n34621,n34622);
  nand U36994(n34622,G59383,n34569);
  nand U36995(n34621,n34570,G58934);
  nand U36996(G1694,n34623,n34624);
  nand U36997(n34624,G59382,n34569);
  nand U36998(n34623,n34570,G58933);
  nand U36999(G1693,n34625,n34626);
  nand U37000(n34626,G59381,n34569);
  nand U37001(n34625,n34570,G58932);
  nand U37002(G1692,n34627,n34628);
  nand U37003(n34628,G59380,n34569);
  nand U37004(n34627,n34570,G58931);
  nand U37005(n34631,G60141,n34632);
  nand U37006(n34630,G59243,n28772);
  not U37007(n28772,G59244);
  nand U37008(n34629,G59692,n21946);
  not U37009(n21946,G59693);
  nand U37010(G1627,n34633,n34634);
  nand U37011(n34634,G58902,G1731);
  nand U37012(n34633,G59693,n34635);
  nand U37013(G1626,n34636,n34637);
  nand U37014(n34637,G58901,G1731);
  nand U37015(n34636,G59692,n34635);
  nand U37016(G1625,n34638,n34639);
  nand U37017(n34639,G58900,G1731);
  nand U37018(n34638,G59691,n34635);
  nand U37019(G1624,n34640,n34641);
  nand U37020(n34641,G58899,G1731);
  nand U37021(n34640,G59690,n34635);
  nand U37022(G1623,n34642,n34643);
  nand U37023(n34643,G58898,G1731);
  nand U37024(n34642,G59689,n34635);
  nand U37025(G1622,n34644,n34645);
  nand U37026(n34645,G58897,G1731);
  nand U37027(n34644,G59688,n34635);
  nand U37028(G1621,n34646,n34647);
  nand U37029(n34647,G58896,G1731);
  nand U37030(n34646,G59687,n34635);
  nand U37031(G1620,n34648,n34649);
  nand U37032(n34649,G58895,G1731);
  nand U37033(n34648,G59686,n34635);
  nand U37034(G1619,n34650,n34651);
  nand U37035(n34651,G58894,G1731);
  nand U37036(n34650,G59685,n34635);
  nand U37037(G1618,n34652,n34653);
  nand U37038(n34653,G58893,G1731);
  nand U37039(n34652,G59684,n34635);
  nand U37040(G1617,n34654,n34655);
  nand U37041(n34655,G58892,G1731);
  nand U37042(n34654,G59683,n34635);
  nand U37043(G1616,n34656,n34657);
  nand U37044(n34657,G58891,G1731);
  nand U37045(n34656,G59682,n34635);
  nand U37046(G1615,n34658,n34659);
  nand U37047(n34659,G58890,G1731);
  nand U37048(n34658,G59681,n34635);
  nand U37049(G1614,n34660,n34661);
  nand U37050(n34661,G58889,G1731);
  nand U37051(n34660,G59680,n34635);
  nand U37052(G1613,n34662,n34663);
  nand U37053(n34663,G58888,G1731);
  nand U37054(n34662,G59679,n34635);
  nand U37055(G1612,n34664,n34665);
  nand U37056(n34665,G58887,G1731);
  nand U37057(n34664,G59678,n34635);
  nand U37058(G1611,n34666,n34667);
  nand U37059(n34667,G58886,G1731);
  nand U37060(n34666,G59677,n34635);
  nand U37061(G1610,n34668,n34669);
  nand U37062(n34669,G58885,G1731);
  nand U37063(n34668,G59676,n34635);
  nand U37064(G1609,n34670,n34671);
  nand U37065(n34671,G58884,G1731);
  nand U37066(n34670,G59675,n34635);
  nand U37067(G1608,n34672,n34673);
  nand U37068(n34673,G58883,G1731);
  nand U37069(n34672,G59674,n34635);
  nand U37070(G1607,n34674,n34675);
  nand U37071(n34675,G58882,G1731);
  nand U37072(n34674,G59673,n34635);
  nand U37073(G1606,n34676,n34677);
  nand U37074(n34677,G58881,G1731);
  nand U37075(n34676,G59672,n34635);
  nand U37076(G1605,n34678,n34679);
  nand U37077(n34679,G58880,G1731);
  nand U37078(n34678,G59671,n34635);
  nand U37079(G1604,n34680,n34681);
  nand U37080(n34681,G58879,G1731);
  nand U37081(n34680,G59670,n34635);
  nand U37082(G1603,n34682,n34683);
  nand U37083(n34683,G58878,G1731);
  nand U37084(n34682,G59669,n34635);
  nand U37085(G1602,n34684,n34685);
  nand U37086(n34685,G58877,G1731);
  nand U37087(n34684,G59668,n34635);
  nand U37088(G1601,n34686,n34687);
  nand U37089(n34687,G58876,G1731);
  nand U37090(n34686,G59667,n34635);
  nand U37091(G1600,n34688,n34689);
  nand U37092(n34689,G58875,G1731);
  nand U37093(n34688,G59666,n34635);
  nand U37094(G1599,n34690,n34691);
  nand U37095(n34691,G58874,G1731);
  nand U37096(n34690,G59665,n34635);
  nand U37097(G1598,n34692,n34693);
  nand U37098(n34693,G58873,G1731);
  nand U37099(n34692,G59664,n34635);
  nand U37100(G1597,n34694,n34695);
  nand U37101(n34695,G58872,G1731);
  nand U37102(n34694,G59663,n34635);
  nand U37103(G1596,n34696,n34697);
  nand U37104(n34697,G58871,G1731);
  nand U37105(n34696,G59662,n34635);
  nand U37106(G1587,n34698,n34699,n34700);
  nand U37107(n34700,G60142,n20962);
  nand U37108(n34699,n20961,G59693);
  nand U37109(n34698,n34701,G58870);
  nand U37110(G1586,n34702,n34703,n34704);
  nand U37111(n34704,G60141,n20962);
  nand U37112(n34703,n20961,G59692);
  nand U37113(n34702,n34701,G58869);
  nand U37114(G1585,n34705,n34706,n34707);
  nand U37115(n34707,G60140,n20962);
  nand U37116(n34706,n20961,G59691);
  nand U37117(n34705,n34701,G58868);
  nand U37118(G1584,n34708,n34709,n34710);
  nand U37119(n34710,G60139,n20962);
  nand U37120(n34709,n20961,G59690);
  nand U37121(n34708,n34701,G58867);
  nand U37122(G1583,n34711,n34712,n34713);
  nand U37123(n34713,G60138,n20962);
  nand U37124(n34712,n20961,G59689);
  nand U37125(n34711,n34701,G58866);
  nand U37126(G1582,n34714,n34715,n34716);
  nand U37127(n34716,G60137,n20962);
  nand U37128(n34715,n20961,G59688);
  nand U37129(n34714,n34701,G58865);
  nand U37130(G1581,n34717,n34718,n34719);
  nand U37131(n34719,G60136,n20962);
  nand U37132(n34718,n20961,G59687);
  nand U37133(n34717,n34701,G58864);
  nand U37134(G1580,n34720,n34721,n34722);
  nand U37135(n34722,G60135,n20962);
  nand U37136(n34721,n20961,G59686);
  nand U37137(n34720,n34701,G58863);
  nand U37138(G1579,n34723,n34724,n34725);
  nand U37139(n34725,G60134,n20962);
  nand U37140(n34724,n20961,G59685);
  nand U37141(n34723,G58862,n34701);
  nand U37142(G1578,n34726,n34727,n34728);
  nand U37143(n34728,G60133,n20962);
  nand U37144(n34727,n20961,G59684);
  nand U37145(n34726,G58861,n34701);
  nand U37146(G1577,n34729,n34730,n34731);
  nand U37147(n34731,G60132,n20962);
  nand U37148(n34730,n20961,G59683);
  nand U37149(n34729,G58860,n34701);
  nand U37150(G1576,n34732,n34733,n34734);
  nand U37151(n34734,G60131,n20962);
  nand U37152(n34733,n20961,G59682);
  nand U37153(n34732,G58859,n34701);
  nand U37154(G1575,n34735,n34736,n34737);
  nand U37155(n34737,G60130,n20962);
  nand U37156(n34736,n20961,G59681);
  nand U37157(n34735,G58858,n34701);
  nand U37158(G1574,n34738,n34739,n34740);
  nand U37159(n34740,G60129,n20962);
  nand U37160(n34739,n20961,G59680);
  nand U37161(n34738,G58857,n34701);
  nand U37162(G1573,n34741,n34742,n34743);
  nand U37163(n34743,G60128,n20962);
  nand U37164(n34742,n20961,G59679);
  nand U37165(n34741,G58856,n34701);
  nand U37166(G1572,n34744,n34745,n34746);
  nand U37167(n34746,G60127,n20962);
  nand U37168(n34745,n20961,G59678);
  nand U37169(n34744,G58855,n34701);
  nand U37170(G1571,n34747,n34748,n34749);
  nand U37171(n34749,G60126,n20962);
  nand U37172(n34748,n20961,G59677);
  nand U37173(n34747,n34701,G58854);
  nand U37174(G1570,n34750,n34751,n34752);
  nand U37175(n34752,G60125,n20962);
  nand U37176(n34751,n20961,G59676);
  nand U37177(n34750,G58853,n34701);
  nand U37178(G1569,n34753,n34754,n34755);
  nand U37179(n34755,G60124,n20962);
  nand U37180(n34754,n20961,G59675);
  nand U37181(n34753,G58852,n34701);
  nand U37182(G1568,n34756,n34757,n34758);
  nand U37183(n34758,G60123,n20962);
  nand U37184(n34757,n20961,G59674);
  nand U37185(n34756,G58851,n34701);
  nand U37186(G1567,n34759,n34760,n34761);
  nand U37187(n34761,G60122,n20962);
  nand U37188(n34760,n20961,G59673);
  nand U37189(n34759,G58850,n34701);
  nand U37190(G1566,n34762,n34763,n34764);
  nand U37191(n34764,G60121,n20962);
  nand U37192(n34763,n20961,G59672);
  nand U37193(n34762,G58849,n34701);
  nand U37194(G1565,n34765,n34766,n34767);
  nand U37195(n34767,G60120,n20962);
  nand U37196(n34766,n20961,G59671);
  nand U37197(n34765,G58848,n34701);
  nand U37198(G1564,n34768,n34769,n34770);
  nand U37199(n34770,G60119,n20962);
  nand U37200(n34769,n20961,G59670);
  nand U37201(n34768,G58847,n34701);
  nand U37202(G1563,n34771,n34772,n34773);
  nand U37203(n34773,G60118,n20962);
  nand U37204(n34772,n20961,G59669);
  nand U37205(n34771,G58846,n34701);
  nand U37206(G1562,n34774,n34775,n34776);
  nand U37207(n34776,G60117,n20962);
  nand U37208(n34775,n20961,G59668);
  nand U37209(n34774,G58845,n34701);
  nand U37210(G1561,n34777,n34778,n34779);
  nand U37211(n34779,G60116,n20962);
  nand U37212(n34778,n20961,G59667);
  nand U37213(n34777,G58844,n34701);
  nand U37214(G1560,n34780,n34781,n34782);
  nand U37215(n34782,G60115,n20962);
  nand U37216(n34781,n20961,G59666);
  nand U37217(n34780,G58843,n34701);
  nand U37218(G1559,n34783,n34784,n34785);
  nand U37219(n34785,G60114,n20962);
  nand U37220(n34784,n20961,G59665);
  nand U37221(n34783,G58842,n34701);
  nand U37222(G1558,n34786,n34787,n34788);
  nand U37223(n34788,G60113,n20962);
  nand U37224(n34787,n20961,G59664);
  nand U37225(n34786,G58841,n34701);
  nand U37226(G1557,n34789,n34790,n34791);
  nand U37227(n34791,G60112,n20962);
  nand U37228(n34790,n20961,G59663);
  nand U37229(n34789,G58840,n34701);
  nand U37230(G1556,n34792,n34793,n34794);
  nand U37231(n34794,G60111,n20962);
  nand U37232(n34793,n20961,G59662);
  nand U37233(n34792,G58839,n34701);
  nand U37234(G1553,n34796,n34797,n34798,n34799);
  nor U37235(n34799,G58908,G58907,n34635,n34800);
  not U37236(n34800,G59351);
  nor U37237(n34798,G59345,G59353,G59350);
  not U37238(n34797,G58910);
  not U37239(n34796,G58909);
  nand U37240(G1552,n34795,G1730);
  nand U37241(n34803,n34804,n34805,G60243,G60249);
  not U37242(n34804,G59805);
  or U37243(n34802,G59808,G60251,G60248);
  nor U37244(n34795,n34801,n21776);
  nor U37245(n34810,n34811,n34812);
  or U37246(n34812,G59382,G59383,G59384,G59385);
  or U37247(n34811,G59386,G59387,G59388,G59389);
  nor U37248(n34809,n34813,G59375,G59377,G59376);
  or U37249(n34813,G59378,G59379,G59380,G59381);
  nor U37250(n34808,n34814,G59368,G59370,G59369);
  or U37251(n34814,G59371,G59372,G59373,G59374);
  nor U37252(n34807,n34815,G59361,G59363,G59362);
  or U37253(n34815,G59364,G59365,G59366,G59367);
  nand U37254(n34801,G59800,G59794,n34816,n34817);
  nor U37255(n34817,G59802,G59799,G59359,G59358);
  nor U37256(n34816,G59357,G59356);
  nand U37257(G15270,n34818,n34819);
  nand U37258(n34819,G59805,n34820);
  nand U37259(n34818,G60239,n34821);
  nand U37260(G15269,n34822,n34823);
  nand U37261(n34823,G59806,n34820);
  nand U37262(n34822,G60240,n34821);
  nand U37263(G15268,n34824,n34825);
  nand U37264(n34825,G59807,n34820);
  nand U37265(n34824,G60241,n34821);
  nand U37266(G15267,n34826,n34827);
  nand U37267(n34827,G59808,n34820);
  nand U37268(n34826,G60242,n34821);
  nand U37269(G15266,n34828,n34829);
  nand U37270(n34829,n34830,n20976,n34831);
  nand U37271(n34828,G59842,n34832);
  nand U37272(G15265,n34833,n34834);
  nand U37273(n34834,G59843,n34832);
  nand U37274(n34833,n34835,n34831);
  nand U37275(n34835,n20976,n34830);
  not U37276(n34830,n34836);
  not U37277(n20976,G35);
  nand U37278(G15264,n34837,n34838);
  nand U37279(n34838,n34839,n34840,n34841,n34842);
  nand U37280(n34837,n34843,G60006);
  nand U37281(G15263,n34844,n34845);
  nand U37282(n34845,n34843,G60007);
  nand U37283(n34844,n34846,n34842);
  nand U37284(n34846,n34847,n34848);
  nand U37285(n34848,n34849,n34850);
  nand U37286(n34847,n34839,n34851);
  nand U37287(G15262,n34852,n34853);
  nand U37288(n34853,n34843,G60008);
  nand U37289(n34852,n34854,n34842);
  nand U37290(n34854,n34855,n34856,n34857);
  nand U37291(n34857,n34839,n34858);
  nand U37292(n34856,G59876,n34859,G60016);
  nand U37293(n34855,n34860,n34849);
  nand U37294(G15260,n34861,n34862);
  nand U37295(n34862,n34843,G60009);
  nand U37296(n34861,n34863,n34842);
  nand U37297(n34863,n34864,n34865,n34866);
  nand U37298(n34866,n34839,n34867);
  nand U37299(n34865,G59876,n34868,G60016);
  nand U37300(n34864,n34869,n34849);
  nand U37301(G15259,n34870,n34871);
  nand U37302(n34871,n34843,G60010);
  not U37303(n34843,n34842);
  nand U37304(n34870,n34872,n34842);
  nand U37305(n34842,n34873,n34874,n34875);
  nand U37306(n34875,n34876,n34877);
  nand U37307(n34872,n34878,n34879,n34880);
  nand U37308(n34880,n34839,n34881);
  nand U37309(n34879,G59876,n34882);
  nand U37310(n34882,G60016,n34883);
  nand U37311(n34878,n34849,n34884);
  nor U37312(n34849,n34885,G59875);
  nand U37313(G15258,n34886,n34887);
  or U37314(n34887,n34820,G60252);
  nand U37315(n34886,G60243,n34820);
  nand U37316(G15257,n34888,n34889);
  or U37317(n34889,n34890,n34891);
  nand U37318(n34888,n34892,n34890);
  nand U37319(n34890,n34893,n34894,n34895,n34896);
  nand U37320(n34895,n34897,n34898);
  nand U37321(n34894,G59876,n34899,n34900);
  nand U37322(n34892,n34901,n34902);
  nand U37323(n34902,G59877,n34903);
  nand U37324(n34903,n34904,n34899);
  nand U37325(n34904,n34905,n34906);
  nand U37326(n34906,G59875,n34907);
  nand U37327(n34907,n34908,n34909);
  nand U37328(n34909,n34910,n34911);
  nand U37329(n34910,n34912,n34913);
  nand U37330(n34908,G60246,n34914);
  nand U37331(n34905,n34915,n34912);
  nand U37332(G15256,n34916,n34917);
  nand U37333(n34917,G60249,n34820);
  nand U37334(n34916,G60253,n34821);
  nand U37335(G15255,n34918,n34919);
  nand U37336(n34919,n34920,G60252);
  nand U37337(n34918,n34921,n34922);
  nand U37338(n34921,n34923,n34924,G59875);
  nand U37339(G15254,n34925,n34926);
  nand U37340(n34926,n34920,G60253);
  not U37341(n34920,n34922);
  nand U37342(n34925,n34922,n34927);
  nand U37343(n34922,n34893,n34928);
  nand U37344(n34928,n34929,n34897);
  nand U37345(G14741,n34930,n34931,n34932,n34933);
  nand U37346(n34933,G59877,n34934,n34935);
  nand U37347(n34932,n34936,G60015);
  nand U37348(n34931,n34937,n34938);
  nand U37349(n34930,n34939,n34940);
  nand U37350(G14739,n34832,n34941);
  nand U37351(n34941,G60251,G59841);
  nand U37352(G14738,n34942,n34943);
  nand U37353(n34943,G59877,n34897,n34929);
  nand U37354(n34942,G60250,n34944);
  nand U37355(n34944,n34945,n34876);
  nand U37356(G14737,n34946,n34947,n34948);
  or U37357(n34947,n34820,G60250);
  nand U37358(n34946,G60248,n34820);
  nand U37359(G14736,n34949,n34950,n34948);
  nand U37360(n34948,n34836,n34951);
  nand U37361(n34950,G35,n34831);
  nand U37362(n34949,G60246,n34832);
  nand U37363(G14735,n34952,n34953);
  nand U37364(n34953,n34954,n34955);
  nand U37365(n34954,n34956,n34957);
  nand U37366(n34957,n34958,n34959);
  nand U37367(n34958,n34960,n34961);
  nand U37368(n34961,n34962,n34839);
  nand U37369(n34956,n34885,n34963);
  nand U37370(n34963,n34964,n34965);
  nand U37371(n34965,n34839,n34966);
  nand U37372(n34966,n34967,n34968);
  nand U37373(n34952,G60245,n34969);
  nand U37374(G14734,n34970,n34971);
  nand U37375(n34971,G60244,n34969);
  nand U37376(n34969,n34876,n34955);
  nand U37377(G14733,n34972,n34973,n34974);
  nand U37378(n34973,G60242,n34975);
  nand U37379(n34972,n34976,G60207);
  nand U37380(G14732,n34974,n34977,n34978);
  nand U37381(n34978,G60241,n34975);
  nand U37382(G14731,n34979,n34980,n34981);
  or U37383(n34981,n34974,n34982);
  nand U37384(n34974,n34976,G60208);
  nand U37385(n34980,G60240,n34975);
  nand U37386(n34979,n34983,n34984,n34985,n34976);
  nand U37387(n34985,G60207,G59842);
  nand U37388(G14730,n34986,n34987,n34977);
  nand U37389(n34977,n34976,n34988,n34983,n34982);
  nand U37390(n34987,G60239,n34975);
  nand U37391(n34986,n34983,n34984,n34976);
  not U37392(n34976,n34975);
  nand U37393(n34975,n34989,n34990,n34991,n34992);
  nor U37394(n34992,n34993,n34994,n34995,n34996);
  nand U37395(n34996,n34997,n34998,n34999,n35000);
  nand U37396(n34995,n35001,n35002,n35003,n35004);
  nand U37397(n34994,n35005,n35006,n35007,n35008);
  nand U37398(n34993,n35009,n35010,n35011,n35012);
  nor U37399(n34991,n35013,n35014,G59845,G59844);
  nor U37400(n35014,n34988,n34983);
  not U37401(n34988,G59842);
  nand U37402(n35013,n35015,n35016,n35017,n35018);
  nor U37403(n34990,G59857,G59856,G59855,G59854);
  nor U37404(n34989,G59853,G59852,G59851,G59850);
  not U37405(n34983,G59843);
  nand U37406(G14729,n35019,n35020,n35021,n35022);
  nor U37407(n35022,n35023,n35024,n35025);
  nor U37408(n35025,n35026,n35027);
  and U37409(n35024,n35028,n35029);
  nor U37410(n35023,n35030,n35031);
  nand U37411(n35021,n35032,n35033);
  nand U37412(n35020,n35034,n35035);
  nand U37413(n35019,n35036,G60206);
  nand U37414(G14728,n35037,n35038,n35039,n35040);
  nor U37415(n35040,n35041,n35042,n35043);
  nor U37416(n35043,n35044,n35027);
  nor U37417(n35042,n35045,n35046);
  nor U37418(n35041,n35047,n35031);
  nand U37419(n35039,n35048,n35033);
  nand U37420(n35038,n35034,n35049);
  nand U37421(n35037,n35036,G60205);
  nand U37422(G14727,n35050,n35051,n35052,n35053);
  nor U37423(n35053,n35054,n35055,n35056);
  nor U37424(n35056,n35057,n35027);
  nor U37425(n35055,n35045,n35058);
  nor U37426(n35054,n35059,n35031);
  nand U37427(n35052,n35060,n35033);
  nand U37428(n35051,n35061,n35034);
  nand U37429(n35050,n35036,G60204);
  nand U37430(G14726,n35062,n35063,n35064,n35065);
  nor U37431(n35065,n35066,n35067,n35068);
  nor U37432(n35068,n35069,n35027);
  nor U37433(n35067,n35045,n35070);
  nor U37434(n35066,n35071,n35031);
  nand U37435(n35064,n35072,n35033);
  nand U37436(n35063,n35034,n35073);
  nand U37437(n35062,n35036,G60203);
  nand U37438(G14725,n35074,n35075,n35076,n35077);
  nor U37439(n35077,n35078,n35079,n35080);
  nor U37440(n35080,n35081,n35027);
  nor U37441(n35079,n35045,n35082);
  nor U37442(n35078,n35083,n35031);
  nand U37443(n35076,n35084,n35033);
  nand U37444(n35075,n35034,n35085);
  nand U37445(n35074,n35036,G60202);
  nand U37446(G14724,n35086,n35087,n35088,n35089);
  nor U37447(n35089,n35090,n35091,n35092);
  nor U37448(n35092,n35093,n35027);
  nor U37449(n35091,n35045,n35094);
  nor U37450(n35090,n35095,n35031);
  nand U37451(n35088,n35096,n35033);
  nand U37452(n35087,n35034,n35097);
  nand U37453(n35086,n35036,G60201);
  nand U37454(G14723,n35098,n35099,n35100,n35101);
  nor U37455(n35101,n35102,n35103,n35104);
  nor U37456(n35104,n35105,n35027);
  and U37457(n35103,n35028,n35106);
  nor U37458(n35102,n35107,n35031);
  nand U37459(n35100,n35108,n35033);
  nand U37460(n35099,n35034,n35109);
  nand U37461(n35098,n35036,G60200);
  nand U37462(G14722,n35110,n35111,n35112,n35113);
  nor U37463(n35113,n35114,n35115,n35116);
  nor U37464(n35116,n35117,n35027);
  nor U37465(n35115,n35045,n35118);
  nor U37466(n35114,n35119,n35031);
  nand U37467(n35112,n35120,n35033);
  nand U37468(n35111,n35034,n35121);
  nand U37469(n35110,n35036,G60199);
  nand U37470(G14721,n35122,n35123,n35124,n35125);
  nor U37471(n35125,n35126,n35127,n35128);
  nor U37472(n35128,n35129,n35027);
  nor U37473(n35127,n35045,n35130);
  nor U37474(n35126,n35131,n35031);
  nand U37475(n35124,n35132,n35033);
  nand U37476(n35123,n35034,n35133);
  nand U37477(n35122,n35036,G60198);
  nand U37478(G14720,n35134,n35135,n35136,n35137);
  nor U37479(n35137,n35138,n35139,n35140);
  nor U37480(n35140,n35141,n35027);
  and U37481(n35139,n35028,n35142);
  nor U37482(n35138,n35143,n35031);
  nand U37483(n35136,n35144,n35033);
  nand U37484(n35135,n35034,n35145);
  nand U37485(n35134,n35036,G60197);
  nand U37486(G14719,n35146,n35147,n35148,n35149);
  nor U37487(n35149,n35150,n35151,n35152);
  nor U37488(n35152,n35153,n35027);
  nor U37489(n35151,n35045,n35154);
  nor U37490(n35150,n35155,n35031);
  nand U37491(n35148,n35156,n35033);
  nand U37492(n35147,n35034,n35157);
  nand U37493(n35146,n35036,G60196);
  nand U37494(G14718,n35158,n35159,n35160,n35161);
  nor U37495(n35161,n35162,n35163,n35164);
  nor U37496(n35164,n35165,n35027);
  nor U37497(n35163,n35045,n35166);
  nor U37498(n35162,n35167,n35031);
  nand U37499(n35160,n35168,n35033);
  nand U37500(n35159,n35034,n35169);
  nand U37501(n35158,n35036,G60195);
  nand U37502(G14717,n35170,n35171,n35172,n35173);
  nor U37503(n35173,n35174,n35175,n35176,n35177);
  nor U37504(n35177,n35178,n35179);
  and U37505(n35176,G60194,n35036);
  and U37506(n35175,n35180,n35034);
  nand U37507(n35172,n35181,G60226);
  nand U37508(n35171,n35182,n35028);
  nand U37509(n35170,n35183,G60067);
  nand U37510(G14716,n35184,n35185,n35186,n35187);
  nor U37511(n35187,n35174,n35188,n35189,n35190);
  nor U37512(n35190,n35178,n35191);
  and U37513(n35189,G60193,n35036);
  and U37514(n35188,n35192,n35034);
  nand U37515(n35186,n35181,G60225);
  nand U37516(n35185,n35193,n35028);
  nand U37517(n35184,n35183,G60066);
  nand U37518(G14715,n35194,n35195,n35196,n35197);
  nor U37519(n35197,n35174,n35198,n35199,n35200);
  nor U37520(n35200,n35178,n35201);
  and U37521(n35199,G60192,n35036);
  and U37522(n35198,n35202,n35034);
  nand U37523(n35196,n35181,G60224);
  nand U37524(n35195,n35203,n35028);
  nand U37525(n35194,n35183,G60065);
  nand U37526(G14714,n35204,n35205,n35206,n35207);
  nor U37527(n35207,n35174,n35208,n35209,n35210);
  nor U37528(n35210,n35178,n35211);
  and U37529(n35209,G60191,n35036);
  and U37530(n35208,n35212,n35034);
  nand U37531(n35206,n35181,G60223);
  nand U37532(n35205,n35213,n35028);
  nand U37533(n35204,n35183,G60064);
  nand U37534(G14713,n35214,n35215,n35216,n35217);
  nor U37535(n35217,n35174,n35218,n35219,n35220);
  nor U37536(n35220,n35178,n35221);
  and U37537(n35219,G60190,n35036);
  and U37538(n35218,n35222,n35034);
  nand U37539(n35216,n35181,G60222);
  nand U37540(n35215,n35223,n35028);
  nand U37541(n35214,n35183,G60063);
  nand U37542(G14712,n35224,n35225,n35226,n35227);
  nor U37543(n35227,n35174,n35228,n35229,n35230);
  nor U37544(n35230,n35178,n35231);
  and U37545(n35229,G60189,n35036);
  and U37546(n35228,n35232,n35034);
  nand U37547(n35226,n35181,G60221);
  nand U37548(n35225,n35233,n35028);
  nand U37549(n35224,n35183,G60062);
  nand U37550(G14711,n35234,n35235,n35236,n35237);
  nor U37551(n35237,n35174,n35238,n35239,n35240);
  nor U37552(n35240,n35178,n35241);
  and U37553(n35239,G60188,n35036);
  and U37554(n35238,n35034,n35242);
  nand U37555(n35236,n35181,G60220);
  nand U37556(n35235,n35243,n35028);
  nand U37557(n35234,n35183,G60061);
  nand U37558(G14710,n35244,n35245,n35246,n35247);
  nor U37559(n35247,n35174,n35248,n35249,n35250);
  nor U37560(n35250,n35178,n35251);
  and U37561(n35249,G60187,n35036);
  and U37562(n35248,n35252,n35034);
  nand U37563(n35246,n35181,G60219);
  nand U37564(n35245,n35253,n35028);
  nand U37565(n35244,n35183,G60060);
  nand U37566(G14709,n35254,n35255,n35256,n35257);
  nor U37567(n35257,n35174,n35258,n35259,n35260);
  nor U37568(n35260,n35178,n35261);
  and U37569(n35259,G60186,n35036);
  and U37570(n35258,n35262,n35034);
  nand U37571(n35256,n35181,G60218);
  nand U37572(n35255,n35263,n35028);
  nand U37573(n35254,n35183,G60059);
  nand U37574(G14708,n35264,n35265,n35266,n35267);
  nor U37575(n35267,n35174,n35268,n35269,n35270);
  nor U37576(n35270,n35178,n35271);
  nor U37577(n35269,n35272,n35273);
  nor U37578(n35268,n35274,n35275);
  nand U37579(n35266,n35181,G60217);
  nand U37580(n35265,n35276,n35028);
  nand U37581(n35264,n35183,G60058);
  nand U37582(G14707,n35277,n35278,n35279,n35280);
  nor U37583(n35283,n35178,n35284);
  and U37584(n35282,G60184,n35036);
  and U37585(n35281,n35285,n35034);
  nand U37586(n35279,n35181,G60216);
  nand U37587(n35278,n35286,n35028);
  nand U37588(n35277,n35183,G60057);
  nand U37589(G14706,n35287,n35288,n35289,n35290);
  nor U37590(n35293,n35178,n35294);
  and U37591(n35292,G60183,n35036);
  and U37592(n35291,n35034,n35295);
  nand U37593(n35289,n35181,G60215);
  nand U37594(n35288,n35296,n35028);
  nand U37595(n35287,n35183,G60056);
  nand U37596(G14705,n35297,n35298,n35299,n35300);
  nor U37597(n35303,n35178,n35304);
  and U37598(n35302,G60182,n35036);
  and U37599(n35301,n35034,n35305);
  not U37600(n35034,n35274);
  nand U37601(n35299,n35181,G60214);
  nand U37602(n35298,n35306,n35028);
  nand U37603(n35297,n35183,G60055);
  nand U37604(G14704,n35307,n35308,n35309,n35310);
  nor U37605(n35310,n35174,n35311,n35312,n35313);
  nor U37606(n35313,n35178,n35314);
  nor U37607(n35312,n35315,n35273);
  nor U37608(n35311,n35274,n35316);
  nand U37609(n35309,n35181,G60213);
  nand U37610(n35308,n35317,n35028);
  nand U37611(n35307,n35183,G60054);
  nand U37612(G14703,n35318,n35319,n35320,n35321);
  nor U37613(n35321,n35174,n35322,n35323,n35324);
  nor U37614(n35324,n35178,n35325);
  nor U37615(n35323,n35326,n35273);
  and U37616(n35322,n35327,n35328);
  nand U37617(n35320,n35181,G60212);
  nand U37618(n35319,n35329,n35330);
  nand U37619(n35318,n35183,G60053);
  nand U37620(G14702,n35331,n35332,n35333,n35334);
  nor U37621(n35334,n35174,n35335,n35336,n35337);
  nor U37622(n35337,n35178,n35338);
  not U37623(n35178,n35033);
  nor U37624(n35336,n35339,n35273);
  and U37625(n35335,n35327,n35340);
  nor U37626(n35174,G59876,G59877,n35181);
  nand U37627(n35333,n35181,G60211);
  nand U37628(n35332,n34840,n35330);
  nand U37629(n35331,n35183,G60052);
  nand U37630(G14701,n35341,n35342,n35343,n35344);
  nor U37631(n35344,n35345,n35346,n35347);
  nor U37632(n35347,n35348,n35027);
  nor U37633(n35346,n35349,n35350);
  nor U37634(n35345,n35351,n35031);
  nand U37635(n35343,n35352,n35033);
  nand U37636(n35342,n35353,n35327);
  nand U37637(n35341,n35036,G60178);
  nand U37638(G14700,n35354,n35355,n35356,n35357);
  nor U37639(n35357,n35358,n35359,n35360);
  nor U37640(n35360,n35361,n35027);
  nor U37641(n35359,n35349,n35362);
  nor U37642(n35358,n35363,n35031);
  nand U37643(n35356,n35364,n35033);
  nand U37644(n35355,n35365,n35327);
  nand U37645(n35354,n35036,G60177);
  nand U37646(G14699,n35366,n35367,n35368,n35369);
  nor U37647(n35369,n35370,n35371,n35372);
  nor U37648(n35372,n35373,n35027);
  nor U37649(n35371,n35349,n35374);
  nor U37650(n35370,n34984,n35031);
  nand U37651(n35368,n35375,n35033);
  nand U37652(n35367,n35376,n35327);
  nand U37653(n35366,n35036,G60176);
  nand U37654(G14698,n35377,n35378,n35379,n35380);
  nor U37655(n35380,n35381,n35382,n35383);
  nor U37656(n35383,n35384,n35027);
  not U37657(n35027,n35183);
  nor U37658(n35183,n35181,G59875,n35385);
  nor U37659(n35382,n35349,n35386);
  not U37660(n35349,n35330);
  nand U37661(n35330,n35045,n35387);
  nand U37662(n35387,n35388,n34911,n35389);
  not U37663(n35045,n35028);
  nand U37664(n35028,n35390,n35391);
  nand U37665(n35391,n35032,n35031,G59876);
  nand U37666(n35390,n35392,n35393,n35389);
  nor U37667(n35381,n34982,n35031);
  nand U37668(n35379,n34938,n35033);
  nand U37669(n35033,n35394,n35395);
  nand U37670(n35395,n35389,n35393,n35396,n35397);
  not U37671(n35396,n35398);
  nand U37672(n35394,G59876,n35031,n35399);
  nand U37673(n35378,n35400,n35327);
  nand U37674(n35327,n35401,n35274);
  nand U37675(n35274,n35389,n35392,n34914,n35402);
  nand U37676(n35401,n35031,n35388,n34915);
  nand U37677(n35377,n35036,G60175);
  not U37678(n35036,n35273);
  nand U37679(n35273,n35389,n35403);
  nand U37680(n35403,n35404,n35405);
  nand U37681(n35405,n35398,n35397,n35393);
  not U37682(n35397,n35392);
  nand U37683(n35404,n35402,n35406);
  nand U37684(n35406,n35392,n34914);
  nor U37685(n35389,n34898,n35181);
  not U37686(n35181,n35031);
  nand U37687(n35031,n34893,n35407,n35408,n35409);
  nor U37688(n34893,n35410,n35411);
  nor U37689(n35411,n34964,n34885);
  nor U37690(n34964,n35412,n35413);
  nor U37691(n35413,n35414,n34898,n35415);
  nor U37692(n35412,n35416,n35417);
  nand U37693(G14697,n35418,n35419);
  nand U37694(n35419,n35420,n35032);
  nand U37695(n35418,n35421,G60206);
  nand U37696(G14696,n35422,n35423,n35424);
  nand U37697(n35424,n35421,G60205);
  nand U37698(n35423,n35420,n35048);
  nand U37699(n35422,n35425,n35426);
  nand U37700(G14695,n35427,n35428,n35429);
  nand U37701(n35429,n35421,G60204);
  nand U37702(n35428,n35420,n35060);
  nand U37703(n35427,n35425,n35430);
  nand U37704(G14694,n35431,n35432,n35433);
  nand U37705(n35433,n35421,G60203);
  nand U37706(n35432,n35420,n35072);
  nand U37707(n35431,n35425,n35434);
  nand U37708(G14693,n35435,n35436,n35437);
  nand U37709(n35437,n35421,G60202);
  nand U37710(n35436,n35420,n35084);
  nand U37711(n35435,n35425,n35438);
  nand U37712(G14692,n35439,n35440,n35441);
  nand U37713(n35441,n35421,G60201);
  nand U37714(n35440,n35420,n35096);
  nand U37715(n35439,n35425,n35442);
  nand U37716(G14691,n35443,n35444,n35445);
  nand U37717(n35445,n35421,G60200);
  nand U37718(n35444,n35420,n35108);
  nand U37719(n35443,n35425,n35106);
  nand U37720(G14690,n35446,n35447,n35448);
  nand U37721(n35448,n35421,G60199);
  nand U37722(n35447,n35420,n35120);
  nand U37723(n35446,n35425,n35449);
  nand U37724(G14689,n35450,n35451,n35452);
  nand U37725(n35452,n35421,G60198);
  nand U37726(n35451,n35420,n35132);
  nand U37727(n35450,n35425,n35453);
  nand U37728(G14688,n35454,n35455,n35456);
  nand U37729(n35456,n35421,G60197);
  nand U37730(n35455,n35420,n35144);
  nand U37731(n35454,n35425,n35142);
  nand U37732(G14687,n35457,n35458,n35459);
  nand U37733(n35459,n35421,G60196);
  nand U37734(n35458,n35420,n35156);
  nand U37735(n35457,n35425,n35460);
  nand U37736(G14686,n35461,n35462,n35463);
  nand U37737(n35463,n35421,G60195);
  nand U37738(n35462,n35420,n35168);
  nand U37739(n35461,n35425,n35464);
  nand U37740(G14685,n35465,n35466,n35467);
  nand U37741(n35467,n35421,G60194);
  nand U37742(n35466,n35420,n35468);
  nand U37743(n35465,n35425,n35182);
  nand U37744(G14684,n35469,n35470,n35471);
  nand U37745(n35471,n35421,G60193);
  nand U37746(n35470,n35420,n35472);
  nand U37747(n35469,n35425,n35193);
  nand U37748(G14683,n35473,n35474,n35475);
  nand U37749(n35475,n35421,G60192);
  nand U37750(n35474,n35420,n35476);
  nand U37751(n35473,n35425,n35203);
  nand U37752(G14682,n35477,n35478,n35479);
  nand U37753(n35479,n35421,G60191);
  nand U37754(n35478,n35420,n35480);
  nand U37755(n35477,n35425,n35213);
  nand U37756(G14681,n35481,n35482,n35483);
  nand U37757(n35483,n35421,G60190);
  nand U37758(n35482,n35420,n35484);
  nand U37759(n35481,n35425,n35223);
  nand U37760(G14680,n35485,n35486,n35487);
  nand U37761(n35487,n35421,G60189);
  nand U37762(n35486,n35420,n35488);
  nand U37763(n35485,n35425,n35233);
  nand U37764(G14679,n35489,n35490,n35491);
  nand U37765(n35491,n35421,G60188);
  nand U37766(n35490,n35420,n35492);
  nand U37767(n35489,n35425,n35243);
  nand U37768(G14678,n35493,n35494,n35495);
  nand U37769(n35495,n35421,G60187);
  nand U37770(n35494,n35420,n35496);
  nand U37771(n35493,n35425,n35253);
  nand U37772(G14677,n35497,n35498,n35499);
  nand U37773(n35499,n35421,G60186);
  nand U37774(n35498,n35420,n35500);
  nand U37775(n35497,n35425,n35263);
  nand U37776(G14676,n35501,n35502,n35503);
  nand U37777(n35503,n35421,G60185);
  nand U37778(n35502,n35420,n35504);
  nand U37779(n35501,n35425,n35276);
  nand U37780(G14675,n35505,n35506,n35507);
  nand U37781(n35507,n35421,G60184);
  nand U37782(n35506,n35420,n35508);
  nand U37783(n35505,n35425,n35286);
  nand U37784(G14674,n35509,n35510,n35511);
  nand U37785(n35511,n35421,G60183);
  nand U37786(n35510,n35420,n35512);
  nand U37787(n35509,n35425,n35296);
  nand U37788(G14673,n35513,n35514,n35515);
  nand U37789(n35515,n35421,G60182);
  nand U37790(n35514,n35420,n35516);
  nand U37791(n35513,n35425,n35306);
  nand U37792(G14672,n35517,n35518,n35519);
  nand U37793(n35519,n35421,G60181);
  nand U37794(n35518,n35420,n35520);
  nand U37795(n35517,n35425,n35317);
  nand U37796(G14671,n35521,n35522,n35523);
  nand U37797(n35523,n35421,G60180);
  nand U37798(n35522,n35420,n35524);
  nand U37799(n35521,n35425,n35329);
  nand U37800(G14670,n35525,n35526,n35527);
  nand U37801(n35527,n35421,G60179);
  nand U37802(n35526,n35420,n35528);
  nand U37803(n35525,n35425,n34840);
  nand U37804(G14669,n35529,n35530,n35531);
  nand U37805(n35531,n35421,G60178);
  nand U37806(n35530,n35420,n35352);
  nand U37807(n35529,n35425,n34850);
  nand U37808(G14668,n35532,n35533,n35534);
  nand U37809(n35534,n35421,G60177);
  nand U37810(n35533,n35420,n35364);
  nand U37811(n35532,n35425,n34860);
  nand U37812(G14667,n35535,n35536,n35537);
  nand U37813(n35537,n35421,G60176);
  nand U37814(n35536,n35420,n35375);
  nand U37815(n35535,n35425,n34869);
  nand U37816(G14666,n35538,n35539,n35540);
  nand U37817(n35540,n35421,G60175);
  nand U37818(n35539,n35420,n34938);
  nand U37819(n35538,n35425,n34884);
  nand U37820(n35543,n35546,n34876);
  nand U37821(G14665,n35547,n35548,n35549,n35550);
  nand U37822(n35550,G1,n35551);
  nand U37823(n35549,n35552,G58870);
  nand U37824(n35548,n35553,n35032);
  nand U37825(n35547,n35554,G60174);
  nand U37826(G14664,n35555,n35556,n35557,n35558);
  nor U37827(n35558,n35559,n35560,n35561);
  nor U37828(n35561,n21711,n35562);
  nor U37829(n35560,n35563,n35564);
  nor U37830(n35559,n35565,n35566);
  nand U37831(n35557,n35554,G60173);
  nand U37832(n35556,n35553,n35048);
  nand U37833(n35555,n35567,n35049);
  nand U37834(G14663,n35568,n35569,n35570,n35571);
  nor U37835(n35571,n35572,n35573,n35574);
  nor U37836(n35574,n21723,n35562);
  nor U37837(n35573,n35563,n35575);
  nor U37838(n35572,n35566,n35576);
  nand U37839(n35570,n35554,G60172);
  nand U37840(n35569,n35553,n35060);
  nand U37841(n35568,n35567,n35061);
  nand U37842(G14662,n35577,n35578,n35579,n35580);
  nor U37843(n35580,n35581,n35582,n35583);
  nor U37844(n35583,n21733,n35562);
  nor U37845(n35582,n35563,n35584);
  nor U37846(n35581,n35566,n35585);
  nand U37847(n35579,n35554,G60171);
  nand U37848(n35578,n35553,n35072);
  nand U37849(n35577,n35567,n35073);
  nand U37850(G14661,n35586,n35587,n35588,n35589);
  nor U37851(n35589,n35590,n35591,n35592);
  nor U37852(n35592,n21743,n35562);
  nor U37853(n35591,n35563,n35593);
  nor U37854(n35590,n35566,n35594);
  nand U37855(n35588,n35554,G60170);
  nand U37856(n35587,n35553,n35084);
  nand U37857(n35586,n35567,n35085);
  nand U37858(G14660,n35595,n35596,n35597,n35598);
  nor U37859(n35598,n35599,n35600,n35601);
  nor U37860(n35601,n21753,n35562);
  nor U37861(n35600,n35563,n35602);
  nor U37862(n35599,n35566,n35603);
  nand U37863(n35597,n35554,G60169);
  nand U37864(n35596,n35553,n35096);
  nand U37865(n35595,n35567,n35097);
  nand U37866(G14659,n35604,n35605,n35606,n35607);
  nor U37867(n35607,n35608,n35609,n35610);
  nor U37868(n35610,n21763,n35562);
  nor U37869(n35609,n35563,n35611);
  nor U37870(n35608,n35566,n35612);
  nand U37871(n35606,n35554,G60168);
  nand U37872(n35605,n35553,n35108);
  nand U37873(n35604,n35567,n35109);
  nand U37874(G14658,n35613,n35614,n35615,n35616);
  nor U37875(n35616,n35617,n35618,n35619);
  nor U37876(n35619,n21775,n35562);
  not U37877(n35562,n35552);
  nor U37878(n35552,n35620,n35621);
  nor U37879(n35618,n35563,n35622);
  not U37880(n35563,n35551);
  nor U37881(n35551,n35620,n34805);
  nor U37882(n35617,n35566,n35623);
  nand U37883(n35615,n35554,G60167);
  nand U37884(n35614,n35553,n35120);
  nand U37885(n35613,n35567,n35121);
  nand U37886(G14657,n35624,n35625,n35626);
  nor U37887(n35626,n35627,n35628,n35629);
  nor U37888(n35629,n35630,n35566);
  nor U37889(n35628,n35620,n35631);
  nor U37890(n35627,n35632,n35633);
  nand U37891(n35625,n35567,n35133);
  nand U37892(n35624,n35554,G60166);
  nand U37893(G14656,n35634,n35635,n35636);
  nor U37894(n35636,n35637,n35638,n35639);
  nor U37895(n35639,n35640,n35566);
  nor U37896(n35638,n35620,n35641);
  nor U37897(n35637,n35642,n35633);
  nand U37898(n35635,n35567,n35145);
  nand U37899(n35634,n35554,G60165);
  nand U37900(G14655,n35643,n35644,n35645);
  nor U37901(n35645,n35646,n35647,n35648);
  nor U37902(n35648,n35649,n35566);
  nor U37903(n35647,n35620,n35650);
  nor U37904(n35646,n35651,n35633);
  nand U37905(n35644,n35567,n35157);
  nand U37906(n35643,n35554,G60164);
  nand U37907(G14654,n35652,n35653,n35654);
  nor U37908(n35654,n35655,n35656,n35657);
  nor U37909(n35657,n35658,n35566);
  nor U37910(n35656,n35620,n35659);
  nor U37911(n35655,n35660,n35633);
  nand U37912(n35653,n35567,n35169);
  nand U37913(n35652,n35554,G60163);
  nand U37914(G14653,n35661,n35662,n35663);
  nor U37915(n35663,n35664,n35665,n35666);
  nor U37916(n35666,n35667,n35566);
  nor U37917(n35665,n35620,n35668);
  nor U37918(n35664,n35179,n35633);
  nand U37919(n35662,n35567,n35180);
  nand U37920(n35661,n35554,G60162);
  nand U37921(G14652,n35669,n35670,n35671);
  nor U37922(n35671,n35672,n35673,n35674);
  nor U37923(n35674,n35675,n35566);
  nor U37924(n35673,n35620,n35676);
  nor U37925(n35672,n35191,n35633);
  nand U37926(n35670,n35567,n35192);
  nand U37927(n35669,n35554,G60161);
  nand U37928(G14651,n35677,n35678,n35679);
  nor U37929(n35679,n35680,n35681,n35682);
  nor U37930(n35682,n35683,n35566);
  nor U37931(n35681,n35620,n35684);
  nor U37932(n35680,n35201,n35633);
  nand U37933(n35678,n35567,n35202);
  nand U37934(n35677,n35554,G60160);
  nand U37935(G14650,n35685,n35686,n35687);
  nor U37936(n35687,n35688,n35689,n35690);
  nor U37937(n35690,n35691,n35566);
  nand U37938(n35566,n35692,n35693);
  nor U37939(n35689,n35620,n35694);
  nand U37940(n35620,n35695,n35693);
  nor U37941(n35688,n35211,n35633);
  not U37942(n35633,n35553);
  nand U37943(n35686,n35567,n35212);
  nand U37944(n35685,n35554,G60159);
  nand U37945(G14649,n35696,n35697,n35698,n35699);
  nand U37946(n35699,n35700,n35701);
  nand U37947(n35698,n35553,n35484);
  nand U37948(n35697,n35567,n35222);
  nand U37949(n35696,n35554,G60158);
  nand U37950(G14648,n35702,n35703,n35704,n35705);
  nand U37951(n35705,n35700,n35706);
  nand U37952(n35704,n35553,n35488);
  nand U37953(n35703,n35567,n35232);
  nand U37954(n35702,n35554,G60157);
  nand U37955(G14647,n35707,n35708,n35709,n35710);
  nand U37956(n35710,n35700,n35711);
  nand U37957(n35709,n35553,n35492);
  nand U37958(n35708,n35567,n35242);
  nand U37959(n35707,n35554,G60156);
  nand U37960(G14646,n35712,n35713,n35714,n35715);
  nand U37961(n35715,n35700,n35716);
  nand U37962(n35714,n35553,n35496);
  nand U37963(n35713,n35567,n35252);
  nand U37964(n35712,n35554,G60155);
  nand U37965(G14645,n35717,n35718,n35719,n35720);
  nand U37966(n35720,n35700,n35721);
  nand U37967(n35719,n35553,n35500);
  nand U37968(n35718,n35567,n35262);
  nand U37969(n35717,n35554,G60154);
  nand U37970(G14644,n35722,n35723,n35724,n35725);
  nand U37971(n35725,n35700,n35726);
  nand U37972(n35724,n35553,n35504);
  nand U37973(n35723,n35567,n35727);
  nand U37974(n35722,n35554,G60153);
  nand U37975(G14643,n35728,n35729,n35730,n35731);
  nand U37976(n35731,n35700,n35732);
  nand U37977(n35730,n35553,n35508);
  nand U37978(n35729,n35567,n35285);
  nand U37979(n35728,n35554,G60152);
  nand U37980(G14642,n35733,n35734,n35735,n35736);
  nand U37981(n35736,n35700,n35737);
  nand U37982(n35735,n35553,n35512);
  nand U37983(n35734,n35567,n35295);
  nand U37984(n35733,n35554,G60151);
  nand U37985(G14641,n35738,n35739,n35740,n35741);
  nand U37986(n35741,n35700,n35742);
  nand U37987(n35740,n35553,n35516);
  nand U37988(n35739,n35567,n35305);
  nand U37989(n35738,n35554,G60150);
  nand U37990(G14640,n35743,n35744,n35745,n35746);
  nand U37991(n35746,n35700,n35747);
  nand U37992(n35745,n35553,n35520);
  nand U37993(n35744,n35567,n35748);
  nand U37994(n35743,n35554,G60149);
  nand U37995(G14639,n35749,n35750,n35751,n35752);
  nand U37996(n35752,n35700,n35753);
  nand U37997(n35751,n35553,n35524);
  nand U37998(n35750,n35567,n35328);
  nand U37999(n35749,n35554,G60148);
  nand U38000(G14638,n35754,n35755,n35756,n35757);
  nand U38001(n35757,n35700,n35758);
  nand U38002(n35756,n35553,n35528);
  nand U38003(n35755,n35567,n35340);
  nand U38004(n35754,n35554,G60147);
  nand U38005(G14637,n35759,n35760,n35761,n35762);
  nand U38006(n35762,n35700,n35763);
  nand U38007(n35761,n35553,n35352);
  nand U38008(n35760,n35567,n35353);
  nand U38009(n35759,n35554,G60146);
  nand U38010(G14636,n35764,n35765,n35766,n35767);
  nand U38011(n35767,n35700,n35768);
  nand U38012(n35766,n35553,n35364);
  nand U38013(n35765,n35567,n35365);
  nand U38014(n35764,n35554,G60145);
  nand U38015(G14635,n35769,n35770,n35771,n35772);
  nand U38016(n35772,n35700,n35773);
  nand U38017(n35771,n35553,n35375);
  nand U38018(n35770,n35567,n35376);
  nand U38019(n35769,n35554,G60144);
  nand U38020(G14634,n35774,n35775,n35776,n35777);
  nand U38021(n35777,n35700,n35778);
  nor U38022(n35700,n35554,n35779);
  nand U38023(n35776,n35553,n34938);
  nor U38024(n35553,n35780,n35554);
  nand U38025(n35775,n35567,n35400);
  nand U38026(n35774,n35554,G60143);
  nand U38027(n35693,n35782,n35783);
  nand U38028(n35783,n34839,n35784);
  nand U38029(n35784,n35785,n35786);
  nand U38030(n35786,n35787,n34934);
  nand U38031(n35787,n34967,n35788);
  or U38032(n35788,n35789,n35790);
  nor U38033(G14633,n34632,n35791);
  not U38034(n34632,G60142);
  nand U38035(G14632,n35792,n35793,n35794);
  nand U38036(n35794,n35795,G60141);
  nand U38037(n35793,n35796,G60173);
  nand U38038(n35792,G60096,n35797);
  nand U38039(G14631,n35798,n35799,n35800);
  nand U38040(n35800,n35795,G60140);
  nand U38041(n35799,n35796,G60172);
  nand U38042(n35798,G60097,n35797);
  nand U38043(G14630,n35801,n35802,n35803);
  nand U38044(n35803,n35795,G60139);
  nand U38045(n35802,n35796,G60171);
  nand U38046(n35801,G60098,n35797);
  nand U38047(G14629,n35804,n35805,n35806);
  nand U38048(n35806,n35795,G60138);
  nand U38049(n35805,n35796,G60170);
  nand U38050(n35804,G60099,n35797);
  nand U38051(G14628,n35807,n35808,n35809);
  nand U38052(n35809,n35795,G60137);
  nand U38053(n35808,n35796,G60169);
  nand U38054(n35807,G60100,n35797);
  nand U38055(G14627,n35810,n35811,n35812);
  nand U38056(n35812,n35795,G60136);
  nand U38057(n35811,n35796,G60168);
  nand U38058(n35810,G60101,n35797);
  nand U38059(G14626,n35813,n35814,n35815);
  nand U38060(n35815,n35795,G60135);
  nand U38061(n35814,n35796,G60167);
  nand U38062(n35813,G60102,n35797);
  nand U38063(G14625,n35816,n35817,n35818);
  nand U38064(n35818,n35795,G60134);
  nand U38065(n35817,n35796,G60166);
  nand U38066(n35816,G60103,n35797);
  nand U38067(G14624,n35819,n35820,n35821);
  nand U38068(n35821,n35795,G60133);
  nand U38069(n35820,n35796,G60165);
  nand U38070(n35819,G60104,n35797);
  nand U38071(G14623,n35822,n35823,n35824);
  nand U38072(n35824,n35795,G60132);
  nand U38073(n35823,n35796,G60164);
  nand U38074(n35822,G60105,n35797);
  nand U38075(G14622,n35825,n35826,n35827);
  nand U38076(n35827,n35795,G60131);
  nand U38077(n35826,n35796,G60163);
  nand U38078(n35825,G60106,n35797);
  nand U38079(G14621,n35828,n35829,n35830);
  nand U38080(n35830,n35795,G60130);
  nand U38081(n35829,n35796,G60162);
  nand U38082(n35828,G60107,n35797);
  nand U38083(G14620,n35831,n35832,n35833);
  nand U38084(n35833,n35795,G60129);
  nand U38085(n35832,n35796,G60161);
  nand U38086(n35831,G60108,n35797);
  nand U38087(G14619,n35834,n35835,n35836);
  nand U38088(n35836,n35795,G60128);
  nand U38089(n35835,n35796,G60160);
  nand U38090(n35834,G60109,n35797);
  nand U38091(G14618,n35837,n35838,n35839);
  nand U38092(n35839,n35795,G60127);
  nand U38093(n35838,n35796,G60159);
  and U38094(n35796,n35840,n35692);
  nand U38095(n35837,G60110,n35797);
  nand U38096(G14617,n35841,n35842,n35843);
  nand U38097(n35843,n35795,G60126);
  nand U38098(n35842,G60080,n35797);
  nand U38099(n35841,n35840,G60158);
  nand U38100(G14616,n35844,n35845,n35846);
  nand U38101(n35846,n35795,G60125);
  nand U38102(n35845,G60081,n35797);
  nand U38103(n35844,n35840,G60157);
  nand U38104(G14615,n35847,n35848,n35849);
  nand U38105(n35849,n35795,G60124);
  nand U38106(n35848,G60082,n35797);
  nand U38107(n35847,n35840,G60156);
  nand U38108(G14614,n35850,n35851,n35852);
  nand U38109(n35852,n35795,G60123);
  nand U38110(n35851,G60083,n35797);
  nand U38111(n35850,n35840,G60155);
  nand U38112(G14613,n35853,n35854,n35855);
  nand U38113(n35855,n35795,G60122);
  nand U38114(n35854,G60084,n35797);
  nand U38115(n35853,n35840,G60154);
  nand U38116(G14612,n35856,n35857,n35858);
  nand U38117(n35858,n35795,G60121);
  nand U38118(n35857,G60085,n35797);
  nand U38119(n35856,n35840,G60153);
  nand U38120(G14611,n35859,n35860,n35861);
  nand U38121(n35861,n35795,G60120);
  nand U38122(n35860,G60086,n35797);
  nand U38123(n35859,n35840,G60152);
  nand U38124(G14610,n35862,n35863,n35864);
  nand U38125(n35864,n35795,G60119);
  nand U38126(n35863,G60087,n35797);
  nand U38127(n35862,n35840,G60151);
  nand U38128(G14609,n35865,n35866,n35867);
  nand U38129(n35867,n35795,G60118);
  nand U38130(n35866,G60088,n35797);
  nand U38131(n35865,n35840,G60150);
  nand U38132(G14608,n35868,n35869,n35870);
  nand U38133(n35870,n35795,G60117);
  nand U38134(n35869,G60089,n35797);
  nand U38135(n35868,n35840,G60149);
  nand U38136(G14607,n35871,n35872,n35873);
  nand U38137(n35873,n35795,G60116);
  nand U38138(n35872,G60090,n35797);
  nand U38139(n35871,n35840,G60148);
  nand U38140(G14606,n35874,n35875,n35876);
  nand U38141(n35876,n35795,G60115);
  nand U38142(n35875,G60091,n35797);
  nand U38143(n35874,n35840,G60147);
  nand U38144(G14605,n35877,n35878,n35879);
  nand U38145(n35879,n35795,G60114);
  nand U38146(n35878,G60092,n35797);
  nand U38147(n35877,n35840,G60146);
  nand U38148(G14604,n35880,n35881,n35882);
  nand U38149(n35882,n35795,G60113);
  nand U38150(n35881,G60093,n35797);
  nand U38151(n35880,n35840,G60145);
  nand U38152(G14603,n35883,n35884,n35885);
  nand U38153(n35885,n35795,G60112);
  nand U38154(n35884,G60094,n35797);
  nand U38155(n35883,n35840,G60144);
  nand U38156(G14602,n35886,n35887,n35888);
  nand U38157(n35888,n35795,G60111);
  nand U38158(n35887,G60095,n35797);
  nand U38159(n35886,n35840,G60143);
  nor U38160(n35840,n35385,n35795);
  nand U38161(n35791,n35889,n35890);
  nand U38162(n35890,n35891,n34934);
  nand U38163(n35891,n35892,n35893);
  nand U38164(n35893,n34876,n34914,n35894);
  nand U38165(n35892,n34839,n35895,n35896);
  nand U38166(n35889,n34900,G59876);
  nand U38167(G14601,n35897,n35898,n35899);
  nand U38168(n35899,n35900,G60110);
  nand U38169(n35897,n35901,G60159);
  nand U38170(G14600,n35902,n35903,n35904);
  nand U38171(n35904,n35900,G60109);
  nand U38172(n35902,n35901,G60160);
  nand U38173(G14599,n35905,n35906,n35907);
  nand U38174(n35907,n35900,G60108);
  nand U38175(n35905,n35901,G60161);
  nand U38176(G14598,n35908,n35909,n35910);
  nand U38177(n35910,n35900,G60107);
  nand U38178(n35908,n35901,G60162);
  nand U38179(G14597,n35911,n35912,n35913);
  nand U38180(n35913,n35900,G60106);
  nand U38181(n35911,n35901,G60163);
  nand U38182(G14596,n35914,n35915,n35916);
  nand U38183(n35916,n35900,G60105);
  nand U38184(n35914,n35901,G60164);
  nand U38185(G14595,n35917,n35918,n35919);
  nand U38186(n35919,n35900,G60104);
  nand U38187(n35917,n35901,G60165);
  nand U38188(G14594,n35920,n35921,n35922);
  nand U38189(n35922,n35900,G60103);
  nand U38190(n35920,n35901,G60166);
  nand U38191(G14593,n35923,n35924,n35925);
  nand U38192(n35925,n35900,G60102);
  nand U38193(n35923,n35901,G60167);
  nand U38194(G14592,n35926,n35927,n35928);
  nand U38195(n35928,n35900,G60101);
  nand U38196(n35926,n35901,G60168);
  nand U38197(G14591,n35929,n35930,n35931);
  nand U38198(n35931,n35900,G60100);
  nand U38199(n35929,n35901,G60169);
  nand U38200(G14590,n35932,n35933,n35934);
  nand U38201(n35934,n35900,G60099);
  nand U38202(n35932,n35901,G60170);
  nand U38203(G14589,n35935,n35936,n35937);
  nand U38204(n35937,n35900,G60098);
  nand U38205(n35935,n35901,G60171);
  nand U38206(G14588,n35938,n35939,n35940);
  nand U38207(n35940,n35900,G60097);
  nand U38208(n35938,n35901,G60172);
  nand U38209(G14587,n35941,n35942,n35943);
  nand U38210(n35943,n35900,G60096);
  nand U38211(n35941,n35901,G60173);
  nand U38212(G14586,n35944,n35898,n35945);
  nand U38213(n35945,n35900,G60095);
  nand U38214(n35898,n35946,n35778);
  nand U38215(n35944,n35901,G60143);
  nand U38216(G14585,n35947,n35903,n35948);
  nand U38217(n35948,n35900,G60094);
  nand U38218(n35903,n35946,n35773);
  nand U38219(n35947,n35901,G60144);
  nand U38220(G14584,n35949,n35906,n35950);
  nand U38221(n35950,n35900,G60093);
  nand U38222(n35906,n35946,n35768);
  nand U38223(n35949,n35901,G60145);
  nand U38224(G14583,n35951,n35909,n35952);
  nand U38225(n35952,n35900,G60092);
  nand U38226(n35909,n35946,n35763);
  nand U38227(n35951,n35901,G60146);
  nand U38228(G14582,n35953,n35912,n35954);
  nand U38229(n35954,n35900,G60091);
  nand U38230(n35912,n35946,n35758);
  nand U38231(n35953,n35901,G60147);
  nand U38232(G14581,n35955,n35915,n35956);
  nand U38233(n35956,n35900,G60090);
  nand U38234(n35915,n35946,n35753);
  nand U38235(n35955,n35901,G60148);
  nand U38236(G14580,n35957,n35918,n35958);
  nand U38237(n35958,n35900,G60089);
  nand U38238(n35918,n35946,n35747);
  nand U38239(n35957,n35901,G60149);
  nand U38240(G14579,n35959,n35921,n35960);
  nand U38241(n35960,n35900,G60088);
  nand U38242(n35921,n35946,n35742);
  nand U38243(n35959,n35901,G60150);
  nand U38244(G14578,n35961,n35924,n35962);
  nand U38245(n35962,n35900,G60087);
  nand U38246(n35924,n35946,n35737);
  not U38247(n35737,n35623);
  nand U38248(n35623,n35963,n35964);
  nand U38249(n35964,n34805,n22120);
  not U38250(n22120,G58847);
  or U38251(n35963,G24,n34805);
  nand U38252(n35961,n35901,G60151);
  nand U38253(G14577,n35965,n35927,n35966);
  nand U38254(n35966,n35900,G60086);
  nand U38255(n35927,n35946,n35732);
  not U38256(n35732,n35612);
  nand U38257(n35612,n35967,n35968);
  nand U38258(n35968,n34805,n22126);
  not U38259(n22126,G58848);
  or U38260(n35967,G23,n34805);
  nand U38261(n35965,n35901,G60152);
  nand U38262(G14576,n35969,n35930,n35970);
  nand U38263(n35970,n35900,G60085);
  nand U38264(n35930,n35946,n35726);
  not U38265(n35726,n35603);
  nand U38266(n35603,n35971,n35972);
  nand U38267(n35972,n34805,n22132);
  not U38268(n22132,G58849);
  or U38269(n35971,G22,n34805);
  nand U38270(n35969,n35901,G60153);
  nand U38271(G14575,n35973,n35933,n35974);
  nand U38272(n35974,n35900,G60084);
  nand U38273(n35933,n35946,n35721);
  not U38274(n35721,n35594);
  nand U38275(n35594,n35975,n35976);
  nand U38276(n35976,n34805,n22138);
  not U38277(n22138,G58850);
  or U38278(n35975,G21,n34805);
  nand U38279(n35973,n35901,G60154);
  nand U38280(G14574,n35977,n35936,n35978);
  nand U38281(n35978,n35900,G60083);
  nand U38282(n35936,n35946,n35716);
  not U38283(n35716,n35585);
  nand U38284(n35585,n35979,n35980);
  nand U38285(n35980,n34805,n22144);
  not U38286(n22144,G58851);
  or U38287(n35979,G20,n34805);
  nand U38288(n35977,n35901,G60155);
  nand U38289(G14573,n35981,n35939,n35982);
  nand U38290(n35982,n35900,G60082);
  nand U38291(n35939,n35946,n35711);
  not U38292(n35711,n35576);
  nand U38293(n35576,n35983,n35984);
  nand U38294(n35984,n34805,n22150);
  not U38295(n22150,G58852);
  or U38296(n35983,G19,n34805);
  nand U38297(n35981,n35901,G60156);
  nand U38298(G14572,n35985,n35942,n35986);
  nand U38299(n35986,n35900,G60081);
  nand U38300(n35942,n35946,n35706);
  not U38301(n35706,n35565);
  nand U38302(n35565,n35987,n35988);
  nand U38303(n35988,n34805,n22156);
  not U38304(n22156,G58853);
  or U38305(n35987,G18,n34805);
  nand U38306(n35985,n35901,G60157);
  nand U38307(G14571,n35989,n35990,n35991);
  nand U38308(n35991,n35900,G60080);
  nand U38309(n35990,n35946,n35701);
  nand U38310(n35701,n35992,n35993);
  nand U38311(n35993,G17,n35621);
  nand U38312(n35992,n34805,G58854);
  nor U38313(n35946,n35994,n35900);
  nand U38314(n35989,n35901,G60158);
  nand U38315(n35995,n34876,n34934,n35996);
  nand U38316(n35782,n35410,n34899);
  nor U38317(n35410,n35997,n34959,n35998);
  nand U38318(G14570,n35999,n36000,n36001,n36002);
  nor U38319(n36002,n36003,n36004);
  nor U38320(n36004,n35026,n36005);
  nor U38321(n36003,n35399,n36006);
  nand U38322(n36001,n36007,n35035);
  nand U38323(n36000,n36008,G60238);
  nand U38324(n35999,n36009,n35029);
  nand U38325(G14569,n36010,n36011,n36012,n36013);
  nor U38326(n36013,n36014,n36015);
  nor U38327(n36015,n35044,n36005);
  nor U38328(n36014,n36016,n36006);
  nand U38329(n36012,n36007,n35049);
  nand U38330(n36011,n36008,G60237);
  nand U38331(n36010,n36009,n35426);
  nand U38332(G14568,n36017,n36018,n36019,n36020);
  nor U38333(n36020,n36021,n36022);
  nor U38334(n36022,n35057,n36005);
  nor U38335(n36021,n36023,n36006);
  nand U38336(n36019,n36007,n35061);
  nand U38337(n36018,n36008,G60236);
  nand U38338(n36017,n36009,n35430);
  nand U38339(G14567,n36024,n36025,n36026,n36027);
  nor U38340(n36027,n36028,n36029);
  nor U38341(n36029,n35069,n36005);
  nor U38342(n36028,n36030,n36006);
  nand U38343(n36026,n36007,n35073);
  nand U38344(n36025,n36008,G60235);
  nand U38345(n36024,n36009,n35434);
  nand U38346(G14566,n36031,n36032,n36033,n36034);
  nor U38347(n36034,n36035,n36036);
  nor U38348(n36036,n35081,n36005);
  and U38349(n36035,n35084,n36037);
  nand U38350(n36033,n36007,n35085);
  nand U38351(n36032,n36008,G60234);
  nand U38352(n36031,n36009,n35438);
  nand U38353(G14565,n36038,n36039,n36040,n36041);
  nor U38354(n36041,n36042,n36043);
  nor U38355(n36043,n35093,n36005);
  nor U38356(n36042,n36044,n36006);
  nand U38357(n36040,n36007,n35097);
  nand U38358(n36039,n36008,G60233);
  nand U38359(n36038,n36009,n35442);
  nand U38360(G14564,n36045,n36046,n36047,n36048);
  nor U38361(n36048,n36049,n36050);
  nor U38362(n36050,n35105,n36005);
  nor U38363(n36049,n36051,n36006);
  nand U38364(n36047,n36007,n35109);
  nand U38365(n36046,n36008,G60232);
  nand U38366(n36045,n36009,n35106);
  nand U38367(G14563,n36052,n36053,n36054,n36055);
  nor U38368(n36055,n36056,n36057);
  nor U38369(n36057,n35117,n36005);
  nor U38370(n36056,n36058,n36006);
  nand U38371(n36054,n36007,n35121);
  nand U38372(n36053,n36008,G60231);
  nand U38373(n36052,n36009,n35449);
  nand U38374(G14562,n36059,n36060,n36061,n36062);
  nor U38375(n36062,n36063,n36064);
  nor U38376(n36064,n35129,n36005);
  nor U38377(n36063,n35632,n36006);
  nand U38378(n36061,n36007,n35133);
  nand U38379(n36060,n36008,G60230);
  nand U38380(n36059,n36009,n35453);
  nand U38381(G14561,n36065,n36066,n36067,n36068);
  nor U38382(n36068,n36069,n36070);
  nor U38383(n36070,n35141,n36005);
  not U38384(n35141,G60070);
  nor U38385(n36069,n35642,n36006);
  nand U38386(n36067,n36007,n35145);
  nand U38387(n36066,n36008,G60229);
  nand U38388(n36065,n36009,n35142);
  nand U38389(G14560,n36071,n36072,n36073,n36074);
  nor U38390(n36074,n36075,n36076);
  nor U38391(n36076,n35153,n36005);
  not U38392(n35153,G60069);
  nor U38393(n36075,n35651,n36006);
  nand U38394(n36073,n36007,n35157);
  nand U38395(n36072,n36008,G60228);
  nand U38396(n36071,n36009,n35460);
  nand U38397(G14559,n36077,n36078,n36079,n36080);
  nor U38398(n36080,n36081,n36082);
  nor U38399(n36082,n35165,n36005);
  not U38400(n35165,G60068);
  nor U38401(n36081,n35660,n36006);
  nand U38402(n36079,n36007,n35169);
  nand U38403(n36078,n36008,G60227);
  nand U38404(n36077,n36009,n35464);
  nand U38405(G14558,n36083,n36084,n36085,n36086);
  nor U38406(n36086,n36087,n36088);
  and U38407(n36088,G60067,n36089);
  nor U38408(n36087,n35179,n36006);
  nand U38409(n36085,n36007,n35180);
  nand U38410(n36084,n36008,G60226);
  nand U38411(n36083,n36009,n35182);
  nand U38412(G14557,n36090,n36091,n36092,n36093);
  nor U38413(n36093,n36094,n36095);
  and U38414(n36095,G60066,n36089);
  nor U38415(n36094,n35191,n36006);
  nand U38416(n36092,n36007,n35192);
  nand U38417(n36091,n36008,G60225);
  nand U38418(n36090,n36009,n35193);
  nand U38419(G14556,n36096,n36097,n36098,n36099);
  nor U38420(n36099,n36100,n36101);
  and U38421(n36101,G60065,n36089);
  nor U38422(n36100,n35201,n36006);
  nand U38423(n36098,n36007,n35202);
  nand U38424(n36097,n36008,G60224);
  nand U38425(n36096,n36009,n35203);
  nand U38426(G14555,n36102,n36103,n36104,n36105);
  nor U38427(n36105,n36106,n36107);
  and U38428(n36107,G60064,n36089);
  nor U38429(n36106,n35211,n36006);
  nand U38430(n36104,n36007,n35212);
  nand U38431(n36103,n36008,G60223);
  nand U38432(n36102,n36009,n35213);
  nand U38433(G14554,n36108,n36109,n36110,n36111);
  nor U38434(n36111,n36112,n36113);
  and U38435(n36113,G60063,n36089);
  nor U38436(n36112,n35221,n36006);
  nand U38437(n36110,n36007,n35222);
  nand U38438(n36109,n36008,G60222);
  nand U38439(n36108,n36009,n35223);
  nand U38440(G14553,n36114,n36115,n36116,n36117);
  nor U38441(n36117,n36118,n36119);
  and U38442(n36119,G60062,n36089);
  nor U38443(n36118,n35231,n36006);
  nand U38444(n36116,n36007,n35232);
  nand U38445(n36115,n36008,G60221);
  nand U38446(n36114,n36009,n35233);
  nand U38447(G14552,n36120,n36121,n36122,n36123);
  nor U38448(n36123,n36124,n36125);
  and U38449(n36125,G60061,n36089);
  nor U38450(n36124,n35241,n36006);
  nand U38451(n36122,n36007,n35242);
  nand U38452(n36121,n36008,G60220);
  nand U38453(n36120,n36009,n35243);
  nand U38454(G14551,n36126,n36127,n36128,n36129);
  nor U38455(n36129,n36130,n36131);
  and U38456(n36131,G60060,n36089);
  nor U38457(n36130,n35251,n36006);
  nand U38458(n36128,n36007,n35252);
  nand U38459(n36127,n36008,G60219);
  nand U38460(n36126,n36009,n35253);
  nand U38461(G14550,n36132,n36133,n36134,n36135);
  nor U38462(n36135,n36136,n36137);
  and U38463(n36137,G60059,n36089);
  nor U38464(n36136,n35261,n36006);
  nand U38465(n36134,n36007,n35262);
  nand U38466(n36133,n36008,G60218);
  nand U38467(n36132,n36009,n35263);
  nand U38468(G14549,n36138,n36139,n36140);
  nor U38469(n36140,n36141,n36142,n36143);
  nor U38470(n36143,n36144,n36145);
  nor U38471(n36142,n36146,n36147);
  and U38472(n36141,n35727,n36007);
  nand U38473(n36139,n36037,n35504);
  nand U38474(n36138,n36089,G60058);
  nand U38475(G14548,n36148,n36149,n36150,n36151);
  nor U38476(n36151,n36152,n36153);
  and U38477(n36153,G60057,n36089);
  nor U38478(n36152,n35284,n36006);
  nand U38479(n36150,n36007,n35285);
  nand U38480(n36149,n36008,G60216);
  nand U38481(n36148,n36009,n35286);
  nand U38482(G14547,n36154,n36155,n36156,n36157);
  nor U38483(n36157,n36158,n36159);
  and U38484(n36159,G60056,n36089);
  nor U38485(n36158,n35294,n36006);
  not U38486(n35294,n35512);
  nand U38487(n36156,n36007,n35295);
  nand U38488(n36155,n36008,G60215);
  nand U38489(n36154,n36009,n35296);
  nand U38490(G14546,n36160,n36161,n36162,n36163);
  nor U38491(n36163,n36164,n36165);
  and U38492(n36165,G60055,n36089);
  nor U38493(n36164,n35304,n36006);
  nand U38494(n36162,n36007,n35305);
  nand U38495(n36161,n36008,G60214);
  nand U38496(n36160,n36009,n35306);
  nand U38497(G14545,n36166,n36167,n36168,n36169);
  nor U38498(n36169,n36170,n36171);
  nor U38499(n36171,n36172,n36005);
  nor U38500(n36170,n35314,n36006);
  nand U38501(n36168,n36007,n35748);
  nand U38502(n36167,n36008,G60213);
  nand U38503(n36166,n36009,n35317);
  nand U38504(G14544,n36173,n36174,n36175,n36176);
  nor U38505(n36176,n36177,n36178);
  nor U38506(n36178,n36179,n36005);
  nor U38507(n36177,n35325,n36006);
  nand U38508(n36175,n36007,n35328);
  nand U38509(n36174,n36008,G60212);
  nand U38510(n36173,n36009,n35329);
  nand U38511(G14543,n36180,n36181,n36182,n36183);
  nor U38512(n36183,n36184,n36185);
  nor U38513(n36185,n36186,n36005);
  nor U38514(n36184,n35338,n36006);
  nand U38515(n36182,n36007,n35340);
  nand U38516(n36181,n36008,G60211);
  nand U38517(n36180,n36009,n34840);
  nand U38518(G14542,n36187,n36188,n36189,n36190);
  nor U38519(n36190,n36191,n36192);
  nor U38520(n36192,n35348,n36005);
  nor U38521(n36191,n36193,n36006);
  nand U38522(n36189,n36007,n35353);
  nand U38523(n36188,n36008,G60210);
  nand U38524(n36187,n36009,n34850);
  nand U38525(G14541,n36194,n36195,n36196,n36197);
  nor U38526(n36197,n36198,n36199);
  nor U38527(n36199,n35361,n36005);
  nor U38528(n36198,n36200,n36006);
  nand U38529(n36196,n36007,n35365);
  nand U38530(n36195,n36008,G60209);
  nand U38531(n36194,n36009,n34860);
  nand U38532(G14540,n36201,n36202,n36203,n36204);
  nor U38533(n36204,n36205,n36206);
  nor U38534(n36206,n35373,n36005);
  nor U38535(n36205,n36207,n36006);
  not U38536(n36006,n36037);
  nand U38537(n36203,n36007,n35376);
  nand U38538(n36202,n36008,G60208);
  nand U38539(n36201,n36009,n34869);
  nand U38540(G14539,n36208,n36209,n36210,n36211);
  nand U38541(n36211,n36007,n35400);
  nor U38542(n36210,n36212,n36213);
  nor U38543(n36213,n35386,n36145);
  not U38544(n36145,n36009);
  nor U38545(n36212,n34982,n36147);
  not U38546(n36147,n36008);
  nand U38547(n36209,n36037,n34938);
  nor U38548(n36037,n36215,n36089);
  nand U38549(n36208,n36089,G60048);
  not U38550(n36089,n36005);
  nand U38551(n36005,n34970,n34896);
  nand U38552(n34896,n34897,n35385,n36216);
  or U38553(n34970,n34960,n34959);
  nand U38554(n34960,n36217,G59875,n36218);
  nand U38555(G14538,n36219,n36220,n36221,n36222);
  nor U38556(n36222,n36223,n36224,n36225);
  nor U38557(n36225,G60047,n36226,n36227);
  nor U38558(n36224,n36228,n36229);
  nor U38559(n36228,n36230,n36231);
  nor U38560(n36230,n36232,n36226);
  nor U38561(n36223,n35030,n36233);
  nand U38562(n36221,n36234,n35032);
  nand U38563(n36220,n36235,n35035);
  nand U38564(n35035,n36236,n36237);
  nand U38565(n36237,n36238,n36239);
  nand U38566(n36239,n36240,n36241);
  nand U38567(n36240,n36242,n36243,n36244);
  nand U38568(n36236,n36245,n36241,n36246);
  nand U38569(n36241,n36247,n36248,n36249);
  nand U38570(n36247,n36250,n36246);
  nand U38571(n36245,n36244,n36250);
  not U38572(n36244,n36248);
  nand U38573(n36248,n36251,n36252,n36253,n36254);
  nand U38574(n36254,n35029,n36255);
  nand U38575(n36253,n36238,n35032);
  not U38576(n35032,n35399);
  xor U38577(n35399,n36256,n36257);
  nand U38578(n36256,n36258,n36259);
  nand U38579(n36259,n36260,n34962);
  nand U38580(n36258,n36261,n35998);
  nand U38581(n36261,n36262,n36263,n36260);
  and U38582(n36260,n36264,n36265);
  nand U38583(n36265,G60206,n36266);
  nand U38584(n36264,G60079,n36267);
  nand U38585(n36263,G60047,n36268);
  nand U38586(n36262,G60174,n36269);
  nand U38587(n36252,G60047,n36270);
  nand U38588(n36251,n36271,G60238);
  nand U38589(n36219,n36272,n35029);
  xor U38590(n35029,n36273,n36274);
  nor U38591(n36274,n36275,n36276,n36277);
  nor U38592(n36277,n36214,n35026);
  not U38593(n35026,G60079);
  nor U38594(n36276,n36278,n36229);
  nor U38595(n36275,n35998,n35030);
  not U38596(n35030,G60238);
  nand U38597(G14537,n36279,n36280,n36281,n36282);
  nor U38598(n36282,n36283,n36284,n36285);
  nor U38599(n36285,n35047,n36233);
  nor U38600(n36284,n36286,n36226);
  nor U38601(n36283,n36287,n36288);
  nand U38602(n36281,n36234,n35048);
  nand U38603(n36280,n36235,n35049);
  nand U38604(n35049,n36289,n36290);
  nand U38605(n36290,n36238,n36291);
  nand U38606(n36291,n36250,n36249);
  nand U38607(n36249,n36242,n36243);
  not U38608(n36242,n36292);
  nand U38609(n36250,n36292,n36293);
  nand U38610(n36289,n36294,n36246);
  xnor U38611(n36294,n36292,n36243);
  not U38612(n36243,n36293);
  nand U38613(n36293,n36295,n36296,n36297,n36298);
  nor U38614(n36298,n36299,n36300);
  nor U38615(n36300,n35047,n36301);
  nor U38616(n36299,n36302,n36287);
  nand U38617(n36297,n36238,n35048);
  nand U38618(n36296,n36303,n36304,n36305);
  nand U38619(n36304,n35426,n36306);
  nand U38620(n36303,n36307,n35046);
  nand U38621(n36307,n36308,n36306);
  nor U38622(n36306,n35058,n35070);
  nand U38623(n36295,n35426,n36309);
  nand U38624(n36292,n36310,n36311);
  nand U38625(n36311,n36238,n36312);
  nand U38626(n36312,n36313,n36314);
  or U38627(n36310,n36314,n36313);
  nand U38628(n36279,n36272,n35426);
  not U38629(n35426,n35046);
  nand U38630(n35046,n36315,n36273);
  nand U38631(n36273,n36316,n36317,n36318);
  xnor U38632(n36318,n36319,n36215);
  nand U38633(n36315,n36320,n36321);
  nand U38634(n36321,n36317,n36316);
  xnor U38635(n36320,n36267,n36319);
  nand U38636(n36319,n36322,n36323,n36324,n36325);
  nor U38637(n36325,n36326,n36327);
  nor U38638(n36327,n36214,n35044);
  not U38639(n35044,G60078);
  nor U38640(n36326,n35998,n35047);
  not U38641(n35047,G60237);
  nand U38642(n36324,G60046,n36328);
  nand U38643(n36323,n35048,n36329);
  not U38644(n35048,n36016);
  nand U38645(n36016,n36257,n36330);
  nand U38646(n36330,n36331,n36332);
  or U38647(n36257,n36332,n36331);
  xor U38648(n36331,n36333,n35998);
  nand U38649(n36333,n36334,n36335,n36336,n36337);
  nor U38650(n36337,n36338,n36339);
  and U38651(n36339,n36266,G60205);
  and U38652(n36338,n36269,G60173);
  nand U38653(n36336,G60078,n36267);
  or U38654(n36335,n36286,n34968);
  nand U38655(n36286,n36227,n36340);
  nand U38656(n36340,n36341,n36342);
  not U38657(n36227,n36232);
  nor U38658(n36232,n36342,n36341);
  nand U38659(n36341,n36343,n36344);
  nand U38660(n36344,n34912,n36287);
  not U38661(n36287,G60046);
  nand U38662(n36343,n36345,n36346,n36347,n35692);
  nor U38663(n36347,n36348,n36349);
  nand U38664(n36349,n36350,n36351,n36352,n36353);
  nand U38665(n36353,n36354,G59998);
  nand U38666(n36352,n36355,G59990);
  nand U38667(n36351,n36356,G59982);
  nand U38668(n36350,n36357,G59974);
  nand U38669(n36348,n36358,n36359,n36360,n36361);
  nand U38670(n36361,n36362,G59966);
  nand U38671(n36360,n36363,G59958);
  nand U38672(n36359,n36364,G59950);
  nand U38673(n36358,n36365,G59942);
  nor U38674(n36346,n36366,n36367,n36368,n36369);
  nor U38675(n36369,n36370,n36371);
  nor U38676(n36368,n36372,n36373);
  nor U38677(n36367,n36374,n36375);
  nor U38678(n36366,n36376,n36377);
  nor U38679(n36345,n36378,n36379,n36380,n36381);
  nor U38680(n36381,n36382,n36383);
  nor U38681(n36380,n36384,n36385);
  nor U38682(n36379,n36386,n36387);
  nor U38683(n36378,n36388,n36389);
  nand U38684(n36334,G60046,n36268);
  nand U38685(n36322,n36390,n36391);
  nand U38686(G14536,n36392,n36393,n36394,n36395);
  nor U38687(n36395,n36396,n36397,n36398);
  nor U38688(n36398,n35059,n36233);
  nor U38689(n36397,n36399,n36226);
  nor U38690(n36396,n36400,n36288);
  nand U38691(n36394,n36234,n35060);
  nand U38692(n36393,n36235,n35061);
  xnor U38693(n35061,n36313,n36401);
  xnor U38694(n36401,n36238,n36314);
  nand U38695(n36314,n36402,n36403);
  nand U38696(n36403,n36404,n36246);
  nand U38697(n36404,n36405,n36406);
  or U38698(n36402,n36405,n36406);
  and U38699(n36313,n36407,n36408,n36409,n36410);
  nor U38700(n36410,n36411,n36412);
  nor U38701(n36412,n35059,n36301);
  nor U38702(n36411,n36302,n36400);
  not U38703(n36400,G60045);
  nand U38704(n36409,n36238,n35060);
  nand U38705(n36408,n36413,n36414,n36305);
  nand U38706(n36414,n35070,n35058);
  nand U38707(n36413,n35434,n36415);
  nand U38708(n36415,n36308,n35058);
  nand U38709(n36407,n35430,n36309);
  nand U38710(n36392,n36272,n35430);
  not U38711(n35430,n35058);
  xnor U38712(n35058,n36316,n36317);
  nor U38713(n36317,n36416,n36417);
  xnor U38714(n36316,n36418,n36215);
  nand U38715(n36418,n36419,n36420,n36421,n36422);
  nor U38716(n36422,n36423,n36424);
  nor U38717(n36424,n36214,n35057);
  nor U38718(n36423,n35998,n35059);
  not U38719(n35059,G60236);
  nand U38720(n36421,G60045,n36328);
  nand U38721(n36420,n35060,n36329);
  not U38722(n35060,n36023);
  nand U38723(n36023,n36332,n36425);
  nand U38724(n36425,n36426,n36427);
  or U38725(n36332,n36427,n36426);
  xor U38726(n36426,n34962,n36428);
  nor U38727(n36428,n36429,n36430,n36431,n36432);
  and U38728(n36432,n36266,G60204);
  nor U38729(n36431,n34968,n36399);
  nand U38730(n36399,n36433,n36342);
  nand U38731(n36342,n36434,n36435);
  or U38732(n36433,n36435,n36434);
  nand U38733(n36435,n36436,n36437);
  nand U38734(n36437,G60045,n34912);
  nand U38735(n36436,n36438,n35692);
  nand U38736(n36438,n36439,n36440,n36441,n36442);
  nor U38737(n36442,n36443,n36444,n36445,n36446);
  nor U38738(n36446,n36447,n36371);
  nor U38739(n36445,n36448,n36373);
  nor U38740(n36444,n36449,n36375);
  nor U38741(n36443,n36450,n36377);
  nor U38742(n36441,n36451,n36452,n36453,n36454);
  nor U38743(n36454,n36455,n36383);
  nor U38744(n36453,n36456,n36385);
  nor U38745(n36452,n36457,n36387);
  nor U38746(n36451,n36458,n36389);
  nor U38747(n36440,n36459,n36460,n36461,n36462);
  nor U38748(n36462,n36463,n36464);
  nor U38749(n36461,n36465,n36466);
  nor U38750(n36460,n36467,n36468);
  nor U38751(n36459,n36469,n36470);
  nor U38752(n36439,n36471,n36472,n36473,n36474);
  nor U38753(n36474,n36475,n36476);
  nor U38754(n36473,n36477,n36478);
  nor U38755(n36472,n36479,n36480);
  nor U38756(n36471,n36481,n36482);
  nor U38757(n36430,n36215,n35057);
  not U38758(n35057,G60077);
  nand U38759(n36429,n36483,n36484);
  nand U38760(n36484,G60045,n36268);
  nand U38761(n36483,G60172,n36269);
  nand U38762(n36419,n36390,n36485);
  nand U38763(G14535,n36486,n36487,n36488,n36489);
  nor U38764(n36489,n36490,n36491,n36492);
  nor U38765(n36492,n35071,n36233);
  nor U38766(n36491,n36493,n36226);
  nor U38767(n36490,n36494,n36288);
  nand U38768(n36488,n36234,n35072);
  nand U38769(n36487,n36235,n35073);
  xor U38770(n35073,n36495,n36406);
  nand U38771(n36406,n36496,n36497,n36498,n36499);
  nor U38772(n36499,n36500,n36501);
  nor U38773(n36501,n36302,n36494);
  nor U38774(n36500,n36030,n36246);
  nand U38775(n36498,n36271,G60235);
  nand U38776(n36497,n35434,n36309);
  nand U38777(n36496,n36308,n36305,n35070);
  xnor U38778(n36495,n36246,n36405);
  nand U38779(n36405,n36502,n36503);
  nand U38780(n36503,n36238,n36504);
  or U38781(n36504,n36505,n36506);
  nand U38782(n36502,n36506,n36505);
  nand U38783(n36486,n36272,n35434);
  not U38784(n35434,n35070);
  xnor U38785(n35070,n36416,n36417);
  xor U38786(n36417,n36507,n36215);
  nand U38787(n36507,n36508,n36509,n36510,n36511);
  nor U38788(n36511,n36512,n36513);
  nor U38789(n36513,n36214,n35069);
  not U38790(n35069,G60076);
  nor U38791(n36512,n35998,n35071);
  not U38792(n35071,G60235);
  nand U38793(n36510,G60044,n36328);
  nand U38794(n36509,n35072,n36329);
  not U38795(n35072,n36030);
  nand U38796(n36030,n36427,n36514);
  nand U38797(n36514,n36515,n36516);
  nand U38798(n36516,n36517,n36518);
  nand U38799(n36427,n36518,n36517,n36519);
  not U38800(n36519,n36515);
  xor U38801(n36515,n36520,n35998);
  nand U38802(n36520,n36521,n36522,n36523,n36524);
  nor U38803(n36524,n36525,n36526);
  and U38804(n36526,n36269,G60171);
  nor U38805(n36525,n36527,n36494);
  nand U38806(n36523,G60076,n36267);
  or U38807(n36522,n36493,n34968);
  nand U38808(n36493,n36528,n36529);
  nand U38809(n36529,n36530,n36531);
  not U38810(n36528,n36434);
  nor U38811(n36434,n36531,n36530);
  nand U38812(n36530,n36532,n36533);
  nand U38813(n36533,n34912,n36494);
  not U38814(n36494,G60044);
  nand U38815(n36532,n36534,n36535,n36536,n35692);
  nor U38816(n36536,n36537,n36538);
  nand U38817(n36538,n36539,n36540,n36541,n36542);
  nand U38818(n36542,n36354,G60000);
  nand U38819(n36541,n36355,G59992);
  nand U38820(n36540,n36356,G59984);
  nand U38821(n36539,n36357,G59976);
  nand U38822(n36537,n36543,n36544,n36545,n36546);
  nand U38823(n36546,n36362,G59968);
  nand U38824(n36545,n36363,G59960);
  nand U38825(n36544,n36364,G59952);
  nand U38826(n36543,n36365,G59944);
  nor U38827(n36535,n36547,n36548,n36549,n36550);
  nor U38828(n36550,n36551,n36371);
  nor U38829(n36549,n36552,n36373);
  nor U38830(n36548,n36553,n36375);
  nor U38831(n36547,n36554,n36377);
  nor U38832(n36534,n36555,n36556,n36557,n36558);
  nor U38833(n36558,n36559,n36383);
  nor U38834(n36557,n36560,n36385);
  nor U38835(n36556,n36561,n36387);
  nor U38836(n36555,n36562,n36389);
  nand U38837(n36521,G60203,n36266);
  nand U38838(n36508,n36390,n36563);
  nand U38839(G14534,n36564,n36565,n36566,n36567);
  nor U38840(n36567,n36568,n36569,n36570);
  nor U38841(n36570,n35083,n36233);
  nor U38842(n36569,n36571,n36226);
  nor U38843(n36568,n36572,n36288);
  nand U38844(n36566,n36234,n35084);
  nand U38845(n36565,n36235,n35085);
  xor U38846(n35085,n36573,n36506);
  nand U38847(n36506,n36574,n36575,n36576,n36577);
  nor U38848(n36577,n36578,n36579);
  nor U38849(n36579,n35083,n36301);
  nor U38850(n36578,n36302,n36572);
  nand U38851(n36576,n36238,n35084);
  nand U38852(n36575,n35442,n36580,n36305,n36581);
  nand U38853(n36574,n35438,n36309);
  nand U38854(n36309,n36582,n36583);
  nand U38855(n36583,n36305,n36581);
  not U38856(n36581,n36308);
  nor U38857(n36308,n35094,n36584,n35082);
  xnor U38858(n36573,n36246,n36505);
  nand U38859(n36505,n36585,n36586);
  nand U38860(n36586,n36238,n36587);
  or U38861(n36587,n36588,n36589);
  nand U38862(n36585,n36589,n36588);
  nand U38863(n36564,n36272,n35438);
  not U38864(n35438,n35082);
  nand U38865(n35082,n36590,n36416);
  or U38866(n36416,n36591,n36592);
  nand U38867(n36590,n36592,n36591);
  or U38868(n36591,n36593,n36594,n36595);
  xor U38869(n36592,n36596,n36215);
  nand U38870(n36596,n36597,n36598,n36599,n36600);
  nor U38871(n36600,n36601,n36602);
  nor U38872(n36602,n36214,n35081);
  nor U38873(n36601,n35998,n35083);
  not U38874(n35083,G60234);
  nand U38875(n36599,G60043,n36328);
  nand U38876(n36598,n35084,n36329);
  xor U38877(n35084,n36517,n36518);
  xnor U38878(n36518,n34962,n36603);
  nor U38879(n36603,n36604,n36605,n36606,n36607);
  and U38880(n36607,n36266,G60202);
  nor U38881(n36606,n34968,n36571);
  nand U38882(n36571,n36531,n36608);
  nand U38883(n36608,n36609,n36610);
  or U38884(n36531,n36610,n36609);
  nand U38885(n36609,n36611,n36612);
  nand U38886(n36612,n34912,n36572);
  not U38887(n36572,G60043);
  nand U38888(n36611,n36613,n36614,n36615,n35692);
  nor U38889(n36615,n36616,n36617);
  nand U38890(n36617,n36618,n36619,n36620,n36621);
  nand U38891(n36621,n36354,G60001);
  nand U38892(n36620,n36355,G59993);
  nand U38893(n36619,n36356,G59985);
  nand U38894(n36618,n36357,G59977);
  nand U38895(n36616,n36622,n36623,n36624,n36625);
  nand U38896(n36625,n36362,G59969);
  nand U38897(n36624,n36363,G59961);
  nand U38898(n36623,n36364,G59953);
  nand U38899(n36622,n36365,G59945);
  nor U38900(n36614,n36626,n36627,n36628,n36629);
  nor U38901(n36629,n36630,n36371);
  nor U38902(n36628,n36631,n36373);
  nor U38903(n36627,n36632,n36375);
  nor U38904(n36626,n36633,n36377);
  nor U38905(n36613,n36634,n36635,n36636,n36637);
  nor U38906(n36637,n36638,n36383);
  nor U38907(n36636,n36639,n36385);
  nor U38908(n36635,n36640,n36387);
  nor U38909(n36634,n36641,n36389);
  nor U38910(n36605,n36215,n35081);
  not U38911(n35081,G60075);
  nand U38912(n36604,n36642,n36643);
  nand U38913(n36643,G60043,n36268);
  nand U38914(n36642,G60170,n36269);
  and U38915(n36517,n36644,n36645);
  nand U38916(n36597,n36390,n36646);
  nand U38917(G14533,n36647,n36648,n36649,n36650);
  nor U38918(n36650,n36651,n36652,n36653);
  nor U38919(n36653,n35095,n36233);
  nor U38920(n36652,n36654,n36226);
  nor U38921(n36651,n36655,n36288);
  nand U38922(n36649,n36234,n35096);
  nand U38923(n36648,n36235,n35097);
  xor U38924(n35097,n36656,n36589);
  nand U38925(n36589,n36657,n36658,n36659,n36660);
  nor U38926(n36660,n36661,n36662);
  nor U38927(n36662,n36302,n36655);
  nor U38928(n36661,n36044,n36246);
  nand U38929(n36659,n36271,G60233);
  nand U38930(n36658,n35442,n36663);
  nand U38931(n36657,n36580,n36305,n35094);
  not U38932(n36580,n36584);
  xnor U38933(n36656,n36246,n36588);
  nand U38934(n36588,n36664,n36665);
  nand U38935(n36665,n36238,n36666);
  or U38936(n36666,n36667,n36668);
  nand U38937(n36664,n36668,n36667);
  nand U38938(n36647,n36272,n35442);
  not U38939(n35442,n35094);
  xor U38940(n35094,n36594,n36669);
  nor U38941(n36669,n36593,n36595);
  xnor U38942(n36594,n36670,n36267);
  nand U38943(n36670,n36671,n36672,n36673,n36674);
  nor U38944(n36674,n36675,n36676);
  nor U38945(n36676,n36214,n35093);
  not U38946(n35093,G60074);
  nor U38947(n36675,n35998,n35095);
  not U38948(n35095,G60233);
  nand U38949(n36673,G60042,n36328);
  nand U38950(n36672,n35096,n36329);
  not U38951(n35096,n36044);
  xnor U38952(n36044,n36645,n36644);
  xnor U38953(n36645,n36677,n35998);
  nand U38954(n36677,n36678,n36679,n36680,n36681);
  nor U38955(n36681,n36682,n36683);
  and U38956(n36683,n36269,G60169);
  nor U38957(n36682,n36527,n36655);
  nand U38958(n36680,G60074,n36267);
  or U38959(n36679,n36654,n34968);
  nand U38960(n36654,n36610,n36684);
  nand U38961(n36684,n36685,n36686);
  or U38962(n36610,n36686,n36685);
  nand U38963(n36685,n36687,n36688);
  nand U38964(n36688,n34912,n36655);
  not U38965(n36655,G60042);
  nand U38966(n36687,n36689,n36690,n36691,n35692);
  nor U38967(n36691,n36692,n36693);
  nand U38968(n36693,n36694,n36695,n36696,n36697);
  nand U38969(n36697,n36354,G60002);
  not U38970(n36354,n36482);
  nand U38971(n36696,n36355,G59994);
  not U38972(n36355,n36480);
  nand U38973(n36695,n36356,G59986);
  not U38974(n36356,n36478);
  nand U38975(n36694,n36357,G59978);
  not U38976(n36357,n36476);
  nand U38977(n36692,n36698,n36699,n36700,n36701);
  nand U38978(n36701,n36362,G59970);
  not U38979(n36362,n36470);
  nand U38980(n36700,n36363,G59962);
  not U38981(n36363,n36468);
  nand U38982(n36699,n36364,G59954);
  not U38983(n36364,n36466);
  nand U38984(n36698,n36365,G59946);
  not U38985(n36365,n36464);
  nor U38986(n36690,n36702,n36703,n36704,n36705);
  nor U38987(n36705,n36706,n36371);
  nor U38988(n36704,n36707,n36373);
  nor U38989(n36703,n36708,n36375);
  nor U38990(n36702,n36709,n36377);
  nor U38991(n36689,n36710,n36711,n36712,n36713);
  nor U38992(n36713,n36714,n36383);
  nor U38993(n36712,n36715,n36385);
  nor U38994(n36711,n36716,n36387);
  nor U38995(n36710,n36717,n36389);
  nand U38996(n36678,G60201,n36266);
  nand U38997(n36671,n36390,n36718);
  nand U38998(G14532,n36719,n36720,n36721,n36722);
  nor U38999(n36722,n36723,n36724,n36725);
  nor U39000(n36725,n35107,n36233);
  nor U39001(n36724,n36051,n36726);
  not U39002(n36051,n35108);
  nor U39003(n36723,n36727,n36288);
  nand U39004(n36721,n36272,n35106);
  nand U39005(n36720,n36728,n36686,n36729);
  nand U39006(n36719,n36235,n35109);
  xor U39007(n35109,n36730,n36668);
  nand U39008(n36668,n36731,n36732,n36733,n36734);
  nor U39009(n36734,n36735,n36736);
  nor U39010(n36736,n35107,n36301);
  nor U39011(n36735,n36302,n36727);
  nand U39012(n36733,n36238,n35108);
  nand U39013(n36732,n35449,n36584,n36737);
  nand U39014(n36731,n35106,n36663);
  nand U39015(n36663,n36582,n36738);
  nand U39016(n36738,n36305,n36584);
  nand U39017(n36584,n36739,n35449,n35106,n35453);
  xor U39018(n35106,n36595,n36593);
  xor U39019(n36593,n36740,n36215);
  nand U39020(n36740,n36741,n36742,n36743,n36744);
  nor U39021(n36744,n36745,n36746);
  nor U39022(n36746,n36214,n35105);
  not U39023(n35105,G60073);
  nor U39024(n36745,n35998,n35107);
  not U39025(n35107,G60232);
  nand U39026(n36743,G60041,n36328);
  nand U39027(n36742,n35108,n36329);
  nor U39028(n35108,n36747,n36644);
  nor U39029(n36644,n36748,n36749);
  and U39030(n36747,n36749,n36748);
  nand U39031(n36748,n36750,n36751,n36752);
  xor U39032(n36749,n36753,n35998);
  nand U39033(n36753,n36754,n36755,n36756,n36757);
  nor U39034(n36757,n36758,n36759);
  and U39035(n36759,n36269,G60168);
  nor U39036(n36758,n36527,n36727);
  nand U39037(n36756,G60073,n36267);
  nand U39038(n36755,n36728,n36686,n35545);
  nand U39039(n36686,n36760,n36761,n36762);
  nand U39040(n36761,n34912,n36727);
  not U39041(n36727,G60041);
  or U39042(n36760,n36763,n34912);
  nand U39043(n36728,n36764,n36765,n36766);
  nand U39044(n36765,G60041,n34912);
  nand U39045(n36764,n36763,n35692);
  nand U39046(n36763,n36767,n36768,n36769,n36770);
  nor U39047(n36770,n36771,n36772,n36773,n36774);
  nor U39048(n36774,n36775,n36371);
  nor U39049(n36773,n36776,n36373);
  nor U39050(n36772,n36777,n36375);
  nor U39051(n36771,n36778,n36377);
  nor U39052(n36769,n36779,n36780,n36781,n36782);
  nor U39053(n36782,n36783,n36383);
  nor U39054(n36781,n36784,n36385);
  nor U39055(n36780,n36785,n36387);
  nor U39056(n36779,n36786,n36389);
  nor U39057(n36768,n36787,n36788,n36789,n36790);
  nor U39058(n36790,n36791,n36464);
  nor U39059(n36789,n36792,n36466);
  nor U39060(n36788,n36793,n36468);
  nor U39061(n36787,n36794,n36470);
  nor U39062(n36767,n36795,n36796,n36797,n36798);
  nor U39063(n36798,n36799,n36476);
  nor U39064(n36797,n36800,n36478);
  nor U39065(n36796,n36801,n36480);
  nor U39066(n36795,n36802,n36482);
  nand U39067(n36754,G60200,n36266);
  nand U39068(n36741,n36390,n36803);
  xnor U39069(n36730,n36246,n36667);
  nand U39070(n36667,n36804,n36805);
  nand U39071(n36805,n36238,n36806);
  or U39072(n36806,n36807,n36808);
  nand U39073(n36804,n36808,n36807);
  nand U39074(G14531,n36809,n36810,n36811,n36812);
  nor U39075(n36812,n36813,n36814,n36815);
  nor U39076(n36815,n35119,n36233);
  nor U39077(n36814,n36816,n36226);
  nor U39078(n36813,n36817,n36288);
  nand U39079(n36811,n36234,n35120);
  nand U39080(n36810,n36235,n35121);
  xor U39081(n35121,n36818,n36808);
  nand U39082(n36808,n36819,n36820,n36821,n36822);
  nor U39083(n36822,n36823,n36824);
  nor U39084(n36824,n36302,n36817);
  nor U39085(n36823,n36058,n36246);
  not U39086(n36058,n35120);
  nand U39087(n36821,n36271,G60231);
  nand U39088(n36820,n36737,n35118);
  nor U39089(n36737,n35130,n35781,n36825);
  nand U39090(n36819,n35449,n36826);
  nand U39091(n36826,n36827,n36828);
  nand U39092(n36828,n36305,n35130);
  not U39093(n36827,n36829);
  xnor U39094(n36818,n36246,n36807);
  nand U39095(n36807,n36830,n36831);
  nand U39096(n36831,n36238,n36832);
  or U39097(n36832,n36833,n36834);
  nand U39098(n36830,n36834,n36833);
  nand U39099(n36809,n36272,n35449);
  not U39100(n35449,n35118);
  nand U39101(n35118,n36595,n36835);
  nand U39102(n36835,n36836,n36837);
  or U39103(n36595,n36837,n36836);
  and U39104(n36836,n36838,n36839);
  nand U39105(n36838,n36840,n36841);
  xor U39106(n36837,n36842,n36215);
  nand U39107(n36842,n36843,n36844,n36845,n36846);
  nor U39108(n36846,n36847,n36848);
  nor U39109(n36848,n36214,n35117);
  not U39110(n35117,G60072);
  nor U39111(n36847,n35998,n35119);
  not U39112(n35119,G60231);
  nand U39113(n36845,G60040,n36328);
  nand U39114(n36844,n35120,n36329);
  xnor U39115(n35120,n36849,n36752);
  xor U39116(n36752,n36850,n34962);
  nand U39117(n36850,n36851,n36852,n36853,n36854);
  nor U39118(n36854,n36855,n36856);
  and U39119(n36856,n36269,G60167);
  nor U39120(n36855,n36527,n36817);
  not U39121(n36817,G60040);
  nand U39122(n36853,G60072,n36267);
  or U39123(n36852,n36816,n34968);
  nand U39124(n36816,n36766,n36857);
  nand U39125(n36857,n36858,n36859);
  not U39126(n36766,n36762);
  nor U39127(n36762,n36859,n36858);
  and U39128(n36858,n36860,n36861);
  nand U39129(n36861,G60040,n34912);
  nand U39130(n36860,n36862,n35692);
  nand U39131(n36862,n36863,n36864,n36865,n36866);
  nor U39132(n36866,n36867,n36868,n36869,n36870);
  nor U39133(n36870,n36871,n36371);
  nor U39134(n36869,n36872,n36373);
  nor U39135(n36868,n36873,n36375);
  nor U39136(n36867,n36874,n36377);
  nor U39137(n36865,n36875,n36876,n36877,n36878);
  nor U39138(n36878,n36879,n36383);
  nor U39139(n36877,n36880,n36385);
  nor U39140(n36876,n36881,n36387);
  nor U39141(n36875,n36882,n36389);
  nor U39142(n36864,n36883,n36884,n36885,n36886);
  nor U39143(n36886,n36887,n36464);
  nor U39144(n36885,n36888,n36466);
  nor U39145(n36884,n36889,n36468);
  nor U39146(n36883,n36890,n36470);
  nor U39147(n36863,n36891,n36892,n36893,n36894);
  nor U39148(n36894,n36895,n36476);
  nor U39149(n36893,n36896,n36478);
  nor U39150(n36892,n36897,n36480);
  nor U39151(n36891,n36898,n36482);
  nand U39152(n36859,n36899,n36900);
  nand U39153(n36851,G60199,n36266);
  nand U39154(n36849,n36751,n36750);
  nand U39155(n36843,n36390,n36901);
  nand U39156(G14530,n36902,n36903,n36904,n36905);
  nor U39157(n36905,n36906,n36907,n36908);
  nor U39158(n36908,n35131,n36233);
  nor U39159(n36907,n35632,n36726);
  nor U39160(n36906,n36909,n36288);
  nand U39161(n36904,n36272,n35453);
  nand U39162(n36903,n36729,n36910);
  nand U39163(n36902,n36235,n35133);
  xor U39164(n35133,n36911,n36834);
  nand U39165(n36834,n36912,n36913,n36914,n36915);
  nor U39166(n36915,n36916,n36917);
  nor U39167(n36917,n36302,n36909);
  nor U39168(n36916,n35632,n36246);
  not U39169(n35632,n35132);
  nand U39170(n36914,n36271,G60230);
  nand U39171(n36913,n35453,n36829);
  not U39172(n35453,n35130);
  nand U39173(n36912,n36739,n36305,n35130);
  xnor U39174(n35130,n36840,n36918);
  and U39175(n36918,n36839,n36841);
  nand U39176(n36841,n36919,n36920,n36921);
  nand U39177(n36921,n36390,n36922);
  nand U39178(n36839,n36923,n36922,n36390);
  nand U39179(n36923,n36919,n36920);
  or U39180(n36920,n36924,n36215);
  nand U39181(n36919,n36215,n36924);
  nand U39182(n36924,n36925,n36926,n36927,n36928);
  nor U39183(n36928,n36929,n36930);
  nor U39184(n36930,n36214,n35129);
  not U39185(n35129,G60071);
  nor U39186(n36929,n35998,n35131);
  not U39187(n35131,G60230);
  nand U39188(n36927,G60039,n36328);
  nand U39189(n36926,n35132,n36329);
  xor U39190(n35132,n36750,n36751);
  xnor U39191(n36750,n36931,n35998);
  nand U39192(n36931,n36932,n36933,n36934,n36935);
  nor U39193(n36935,n36936,n36937);
  and U39194(n36937,n36269,G60166);
  nor U39195(n36936,n36527,n36909);
  not U39196(n36909,G60039);
  nand U39197(n36934,G60071,n36267);
  nand U39198(n36933,n35545,n36910);
  xor U39199(n36910,n36899,n36900);
  nand U39200(n36900,n36938,n36939);
  nand U39201(n36939,G60039,n34912);
  nand U39202(n36938,n36940,n35692);
  nand U39203(n36940,n36941,n36942,n36943,n36944);
  nor U39204(n36944,n36945,n36946,n36947,n36948);
  nor U39205(n36948,n36949,n36371);
  nand U39206(n36371,n36950,n36951);
  nor U39207(n36947,n36952,n36373);
  nand U39208(n36373,n36953,n36951);
  nor U39209(n36946,n36954,n36375);
  nand U39210(n36375,n36955,n36951);
  nor U39211(n36945,n36956,n36377);
  nand U39212(n36377,n36957,n36951);
  and U39213(n36951,n36958,n36959);
  nor U39214(n36943,n36960,n36961,n36962,n36963);
  nor U39215(n36963,n36964,n36383);
  nand U39216(n36383,n36965,n36950);
  nor U39217(n36962,n36966,n36385);
  nand U39218(n36385,n36965,n36953);
  nor U39219(n36961,n36967,n36387);
  nand U39220(n36387,n36965,n36955);
  nor U39221(n36960,n36968,n36389);
  nand U39222(n36389,n36965,n36957);
  and U39223(n36965,n36969,n36959);
  nor U39224(n36942,n36970,n36971,n36972,n36973);
  nor U39225(n36973,n36974,n36464);
  nand U39226(n36464,n36975,n36950);
  nor U39227(n36972,n36976,n36466);
  nand U39228(n36466,n36975,n36953);
  nor U39229(n36971,n36977,n36468);
  nand U39230(n36468,n36975,n36955);
  nor U39231(n36970,n36978,n36470);
  nand U39232(n36470,n36975,n36957);
  nor U39233(n36975,n36959,n36969);
  not U39234(n36969,n36958);
  nor U39235(n36941,n36979,n36980,n36981,n36982);
  nor U39236(n36982,n36983,n36476);
  nand U39237(n36476,n36984,n36950);
  nor U39238(n36950,n36985,n36986);
  nor U39239(n36981,n36987,n36478);
  nand U39240(n36478,n36984,n36953);
  nor U39241(n36953,G60010,n36986);
  nor U39242(n36980,n36988,n36480);
  nand U39243(n36480,n36984,n36955);
  nor U39244(n36955,n36989,n36985);
  nor U39245(n36979,n36990,n36482);
  nand U39246(n36482,n36984,n36957);
  nor U39247(n36957,n36989,G60010);
  nor U39248(n36984,n36959,n36958);
  nand U39249(n36899,n36991,n36992);
  nand U39250(n36992,n36993,G60038);
  nand U39251(n36991,n36391,n35692);
  nand U39252(n36391,n36994,n36995,n36996,n36997);
  nor U39253(n36997,n36998,n36999,n37000,n37001);
  nor U39254(n37001,n37002,n37003);
  nor U39255(n37000,n37004,n37005);
  nor U39256(n36999,n37006,n37007);
  nor U39257(n36998,n37008,n37009);
  nor U39258(n36996,n37010,n37011,n37012,n37013);
  nor U39259(n37013,n37014,n37015);
  nor U39260(n37012,n37016,n37017);
  nor U39261(n37011,n37018,n37019);
  nor U39262(n37010,n37020,n37021);
  nor U39263(n36995,n37022,n37023,n37024,n37025);
  nor U39264(n37025,n36382,n37026);
  nor U39265(n37024,n36384,n37027);
  nor U39266(n37023,n36386,n37028);
  nor U39267(n37022,n36388,n37029);
  nor U39268(n36994,n37030,n37031,n37032,n37033);
  nor U39269(n37033,n36370,n37034);
  nor U39270(n37032,n36372,n37035);
  nor U39271(n37031,n36374,n37036);
  nor U39272(n37030,n36376,n37037);
  nand U39273(n36932,G60198,n36266);
  nand U39274(n36925,n36390,n37038);
  nand U39275(n36840,n37039,n37040);
  nand U39276(n37040,n37041,n37042);
  not U39277(n36739,n36825);
  xnor U39278(n36911,n36246,n36833);
  nand U39279(n36833,n37043,n37044);
  nand U39280(n37044,n36238,n37045);
  or U39281(n37045,n37046,n37047);
  nand U39282(n37043,n37047,n37046);
  nand U39283(G14529,n37048,n37049,n37050,n37051);
  nor U39284(n37051,n37052,n37053,n37054);
  nor U39285(n37054,n35143,n36233);
  and U39286(n37053,n37055,n36729);
  nor U39287(n37052,n37056,n36288);
  nand U39288(n37050,n36234,n35144);
  nand U39289(n37049,n36235,n35145);
  xor U39290(n35145,n37057,n37047);
  nand U39291(n37047,n37058,n37059,n37060,n37061);
  nor U39292(n37061,n37062,n37063);
  nor U39293(n37063,n35143,n36301);
  not U39294(n35143,G60229);
  nor U39295(n37062,n36302,n37056);
  nand U39296(n37060,n36238,n35144);
  nand U39297(n37059,n35460,n36825,n37064);
  nand U39298(n37058,n35142,n36829);
  nand U39299(n36829,n36582,n37065);
  nand U39300(n37065,n36305,n36825);
  nand U39301(n36825,n35142,n37066,n35460,n35464);
  xnor U39302(n37057,n36246,n37046);
  nand U39303(n37046,n37067,n37068);
  nand U39304(n37068,n36238,n37069);
  or U39305(n37069,n37070,n37071);
  nand U39306(n37067,n37071,n37070);
  nand U39307(n37048,n36272,n35142);
  xor U39308(n35142,n37042,n37072);
  and U39309(n37072,n37039,n37041);
  nand U39310(n37041,n37073,n37074,n37075);
  nand U39311(n37075,n36390,n37076);
  nand U39312(n37039,n37077,n37076,n36390);
  nand U39313(n37077,n37073,n37074);
  nand U39314(n37074,n36267,n35642,n37078);
  not U39315(n35642,n35144);
  nand U39316(n37073,n37079,n36215);
  nand U39317(n37079,n37078,n37080);
  nand U39318(n37080,n35144,n36329);
  nor U39319(n35144,n37081,n36751);
  nor U39320(n36751,n37082,n37083,n37084);
  and U39321(n37081,n37082,n37085);
  or U39322(n37085,n37084,n37083);
  xor U39323(n37082,n34962,n37086);
  nor U39324(n37086,n37087,n37088,n37089);
  and U39325(n37089,n36269,G60165);
  nor U39326(n37088,n36527,n37056);
  nand U39327(n37087,n37090,n37091,n37092);
  nand U39328(n37092,G60070,n36267);
  nand U39329(n37091,n35545,n37055);
  nand U39330(n37055,n37093,n37094,n37095);
  nand U39331(n37095,n36993,n37056);
  or U39332(n37094,n37056,n36993,n35692);
  nor U39333(n36993,n37096,n37097);
  not U39334(n37056,G60038);
  nand U39335(n37093,n36485,n35692);
  nand U39336(n36485,n37098,n37099,n37100,n37101);
  nor U39337(n37101,n37102,n37103,n37104,n37105);
  nor U39338(n37105,n36475,n37003);
  nor U39339(n37104,n36477,n37005);
  nor U39340(n37103,n36479,n37007);
  nor U39341(n37102,n36481,n37009);
  nor U39342(n37100,n37106,n37107,n37108,n37109);
  nor U39343(n37109,n36463,n37015);
  nor U39344(n37108,n36465,n37017);
  nor U39345(n37107,n36467,n37019);
  nor U39346(n37106,n36469,n37021);
  nor U39347(n37099,n37110,n37111,n37112,n37113);
  nor U39348(n37113,n36455,n37026);
  nor U39349(n37112,n36456,n37027);
  nor U39350(n37111,n36457,n37028);
  nor U39351(n37110,n36458,n37029);
  nor U39352(n37098,n37114,n37115,n37116,n37117);
  nor U39353(n37117,n36447,n37034);
  nor U39354(n37116,n36448,n37035);
  nor U39355(n37115,n36449,n37036);
  nor U39356(n37114,n36450,n37037);
  nand U39357(n37090,G60197,n36266);
  and U39358(n37078,n37118,n37119,n37120);
  nand U39359(n37120,G60070,n37121);
  nand U39360(n37119,G60038,n36328);
  nand U39361(n37118,G60229,n34962);
  nand U39362(n37042,n37122,n37123);
  nand U39363(n37123,n37124,n37125);
  nand U39364(G14528,n37126,n37127,n37128,n37129);
  nor U39365(n37129,n37130,n37131,n37132);
  nor U39366(n37132,n35155,n36233);
  not U39367(n35155,G60228);
  and U39368(n37131,n37133,n36729);
  nor U39369(n37130,n37096,n36288);
  nand U39370(n37128,n36234,n35156);
  nand U39371(n37127,n36235,n35157);
  xor U39372(n35157,n37134,n37071);
  nand U39373(n37071,n37135,n37136,n37137,n37138);
  nor U39374(n37138,n37139,n37140);
  nor U39375(n37140,n36302,n37096);
  nor U39376(n37139,n35651,n36246);
  nand U39377(n37137,n36271,G60228);
  nand U39378(n37136,n35154,n37064);
  nor U39379(n37064,n35166,n35781,n37141);
  nand U39380(n37135,n35460,n37142);
  nand U39381(n37142,n37143,n37144);
  nand U39382(n37144,n36305,n35166);
  not U39383(n37143,n37145);
  xnor U39384(n37134,n36246,n37070);
  nand U39385(n37070,n37146,n37147);
  nand U39386(n37147,n36238,n37148);
  or U39387(n37148,n37149,n37150);
  nand U39388(n37146,n37150,n37149);
  nand U39389(n37126,n36272,n35460);
  not U39390(n35460,n35154);
  xnor U39391(n35154,n37125,n37151);
  and U39392(n37151,n37122,n37124);
  nand U39393(n37124,n37152,n37153,n37154);
  nand U39394(n37154,n36390,n37155);
  nand U39395(n37122,n37156,n37155,n36390);
  nand U39396(n37156,n37152,n37153);
  nand U39397(n37153,n36267,n35651,n37157);
  nand U39398(n37152,n37158,n36215);
  nand U39399(n37158,n37157,n37159);
  nand U39400(n37159,n35156,n36329);
  not U39401(n35156,n35651);
  xnor U39402(n35651,n37084,n37083);
  xor U39403(n37083,n34962,n37160);
  nor U39404(n37160,n37161,n37162,n37163);
  and U39405(n37163,n36269,G60164);
  nor U39406(n37162,n36527,n37096);
  not U39407(n37096,G60037);
  nand U39408(n37161,n37164,n37165,n37166);
  nand U39409(n37166,G60069,n36267);
  nand U39410(n37165,n35545,n37133);
  nand U39411(n37133,n37167,n37168);
  nand U39412(n37168,n36563,n35692);
  nand U39413(n36563,n37169,n37170,n37171,n37172);
  nor U39414(n37172,n37173,n37174,n37175,n37176);
  nor U39415(n37176,n37177,n37003);
  nor U39416(n37175,n37178,n37005);
  nor U39417(n37174,n37179,n37007);
  nor U39418(n37173,n37180,n37009);
  nor U39419(n37171,n37181,n37182,n37183,n37184);
  nor U39420(n37184,n37185,n37015);
  nor U39421(n37183,n37186,n37017);
  nor U39422(n37182,n37187,n37019);
  nor U39423(n37181,n37188,n37021);
  nor U39424(n37170,n37189,n37190,n37191,n37192);
  nor U39425(n37192,n36559,n37026);
  nor U39426(n37191,n36560,n37027);
  nor U39427(n37190,n36561,n37028);
  nor U39428(n37189,n36562,n37029);
  nor U39429(n37169,n37193,n37194,n37195,n37196);
  nor U39430(n37196,n36551,n37034);
  nor U39431(n37195,n36552,n37035);
  nor U39432(n37194,n36553,n37036);
  nor U39433(n37193,n36554,n37037);
  nand U39434(n37167,n37197,n34912);
  xnor U39435(n37197,G60037,n37097);
  nand U39436(n37097,n37198,G60036);
  nand U39437(n37164,G60196,n36266);
  and U39438(n37157,n37199,n37200,n37201);
  nand U39439(n37201,G60069,n37121);
  nand U39440(n37200,G60037,n36328);
  nand U39441(n37199,G60228,n34962);
  nand U39442(n37125,n37202,n37203);
  nand U39443(n37203,n37204,n37205);
  nand U39444(G14527,n37206,n37207,n37208,n37209);
  nor U39445(n37209,n37210,n37211,n37212);
  nor U39446(n37212,n35167,n36233);
  not U39447(n35167,G60227);
  and U39448(n37211,n37213,n36729);
  nor U39449(n37210,n37214,n36288);
  nand U39450(n37208,n36234,n35168);
  nand U39451(n37207,n36235,n35169);
  xor U39452(n35169,n37215,n37150);
  nand U39453(n37150,n37216,n37217,n37218,n37219);
  nor U39454(n37219,n37220,n37221);
  nor U39455(n37221,n36302,n37214);
  nor U39456(n37220,n35660,n36246);
  nand U39457(n37218,n36271,G60227);
  nand U39458(n37217,n35464,n37145);
  nand U39459(n37216,n37066,n36305,n35166);
  not U39460(n37066,n37141);
  xnor U39461(n37215,n36246,n37149);
  nand U39462(n37149,n37222,n37223);
  nand U39463(n37223,n36238,n37224);
  or U39464(n37224,n37225,n37226);
  nand U39465(n37222,n37226,n37225);
  nand U39466(n37206,n36272,n35464);
  not U39467(n35464,n35166);
  xnor U39468(n35166,n37205,n37227);
  and U39469(n37227,n37202,n37204);
  nand U39470(n37204,n37228,n37229,n37230);
  nand U39471(n37202,n37232,n37231,n36390);
  nand U39472(n37232,n37228,n37229);
  nand U39473(n37229,n36267,n35660,n37233);
  nand U39474(n37228,n37234,n36215);
  nand U39475(n37234,n37233,n37235);
  nand U39476(n37235,n35168,n36329);
  not U39477(n35168,n35660);
  nand U39478(n35660,n37084,n37236);
  nand U39479(n37236,n37237,n37238);
  or U39480(n37084,n37238,n37237);
  xor U39481(n37237,n34962,n37239);
  nor U39482(n37239,n37240,n37241,n37242);
  and U39483(n37242,n36269,G60163);
  nor U39484(n37241,n36527,n37214);
  nand U39485(n37240,n37243,n37244,n37245);
  nand U39486(n37245,G60068,n36267);
  nand U39487(n37244,n35545,n37213);
  nand U39488(n37213,n37246,n37247,n37248);
  nand U39489(n37248,n37198,n37214);
  or U39490(n37247,n37214,n37198,n35692);
  nor U39491(n37198,n37249,n37250);
  not U39492(n37214,G60036);
  nand U39493(n37246,n36646,n35692);
  nand U39494(n36646,n37251,n37252,n37253,n37254);
  nor U39495(n37254,n37255,n37256,n37257,n37258);
  nor U39496(n37258,n37259,n37003);
  nor U39497(n37257,n37260,n37005);
  nor U39498(n37256,n37261,n37007);
  nor U39499(n37255,n37262,n37009);
  nor U39500(n37253,n37263,n37264,n37265,n37266);
  nor U39501(n37266,n37267,n37015);
  nor U39502(n37265,n37268,n37017);
  nor U39503(n37264,n37269,n37019);
  nor U39504(n37263,n37270,n37021);
  nor U39505(n37252,n37271,n37272,n37273,n37274);
  nor U39506(n37274,n36638,n37026);
  nor U39507(n37273,n36639,n37027);
  nor U39508(n37272,n36640,n37028);
  nor U39509(n37271,n36641,n37029);
  nor U39510(n37251,n37275,n37276,n37277,n37278);
  nor U39511(n37278,n36630,n37034);
  nor U39512(n37277,n36631,n37035);
  nor U39513(n37276,n36632,n37036);
  nor U39514(n37275,n36633,n37037);
  nand U39515(n37243,G60195,n36266);
  and U39516(n37233,n37279,n37280,n37281);
  nand U39517(n37281,G60068,n37121);
  nand U39518(n37280,G60036,n36328);
  nand U39519(n37279,G60227,n34962);
  nand U39520(n37205,n37282,n37283);
  nand U39521(n37283,n37284,n37285);
  nand U39522(G14526,n37286,n37287,n37288,n37289);
  nor U39523(n37289,n37290,n37291,n37292);
  nor U39524(n37292,n37293,n36233);
  and U39525(n37291,n37294,n36729);
  nor U39526(n37290,n37250,n36288);
  nand U39527(n37288,n36234,n35468);
  nand U39528(n37287,n36235,n35180);
  xor U39529(n35180,n37295,n37226);
  nand U39530(n37226,n37296,n37297,n37298,n37299);
  nor U39531(n37299,n37300,n37301);
  nor U39532(n37301,n37293,n36301);
  not U39533(n37293,G60226);
  nor U39534(n37300,n36302,n37250);
  nand U39535(n37298,n36238,n35468);
  nand U39536(n37297,n35203,n37302,n35193,n37141);
  nand U39537(n37296,n35182,n37145);
  nand U39538(n37145,n36582,n37303);
  nand U39539(n37303,n36305,n37141);
  nand U39540(n37141,n35213,n37304,n35193,n37305);
  and U39541(n37305,n35182,n35203);
  xnor U39542(n37295,n36246,n37225);
  nand U39543(n37225,n37306,n37307);
  nand U39544(n37307,n36238,n37308);
  or U39545(n37308,n37309,n37310);
  nand U39546(n37306,n37310,n37309);
  nand U39547(n37286,n36272,n35182);
  xor U39548(n35182,n37285,n37311);
  and U39549(n37311,n37282,n37284);
  nand U39550(n37284,n37312,n37313,n37314);
  nand U39551(n37282,n37316,n37315,n36390);
  nand U39552(n37316,n37312,n37313);
  nand U39553(n37313,n36267,n35179,n37317);
  nand U39554(n37312,n37318,n36215);
  nand U39555(n37318,n37317,n37319);
  nand U39556(n37319,n35468,n36329);
  not U39557(n35468,n35179);
  nand U39558(n35179,n37320,n37238);
  or U39559(n37238,n37321,n37322,n37323);
  nand U39560(n37320,n37321,n37324);
  or U39561(n37324,n37323,n37322);
  xor U39562(n37321,n34962,n37325);
  nor U39563(n37325,n37326,n37327,n37328);
  and U39564(n37328,n36269,G60162);
  nor U39565(n37327,n36527,n37250);
  not U39566(n37250,G60035);
  nand U39567(n37326,n37329,n37330,n37331);
  nand U39568(n37331,G60067,n36267);
  nand U39569(n37330,n35545,n37294);
  nand U39570(n37294,n37332,n37333);
  nand U39571(n37333,n36718,n35692);
  nand U39572(n36718,n37334,n37335,n37336,n37337);
  nor U39573(n37337,n37338,n37339,n37340,n37341);
  nor U39574(n37341,n37342,n37003);
  nor U39575(n37340,n37343,n37005);
  nor U39576(n37339,n37344,n37007);
  nor U39577(n37338,n37345,n37009);
  nor U39578(n37336,n37346,n37347,n37348,n37349);
  nor U39579(n37349,n37350,n37015);
  nor U39580(n37348,n37351,n37017);
  nor U39581(n37347,n37352,n37019);
  nor U39582(n37346,n37353,n37021);
  nor U39583(n37335,n37354,n37355,n37356,n37357);
  nor U39584(n37357,n36714,n37026);
  nor U39585(n37356,n36715,n37027);
  nor U39586(n37355,n36716,n37028);
  nor U39587(n37354,n36717,n37029);
  nor U39588(n37334,n37358,n37359,n37360,n37361);
  nor U39589(n37361,n36706,n37034);
  nor U39590(n37360,n36707,n37035);
  nor U39591(n37359,n36708,n37036);
  nor U39592(n37358,n36709,n37037);
  nand U39593(n37332,n37362,n34912);
  xnor U39594(n37362,G60035,n37249);
  or U39595(n37249,n37363,n37364);
  nand U39596(n37329,G60194,n36266);
  and U39597(n37317,n37365,n37366,n37367);
  nand U39598(n37367,G60067,n37121);
  nand U39599(n37366,G60035,n36328);
  nand U39600(n37365,G60226,n34962);
  nand U39601(n37285,n37368,n37369);
  nand U39602(n37369,n37370,n37371);
  nand U39603(G14525,n37372,n37373,n37374,n37375);
  nor U39604(n37375,n37376,n37377,n37378);
  nor U39605(n37378,n37379,n36233);
  not U39606(n37379,G60225);
  and U39607(n37377,n37380,n36729);
  nor U39608(n37376,n37363,n36288);
  nand U39609(n37374,n36234,n35472);
  nand U39610(n37373,n36235,n35192);
  xor U39611(n35192,n37381,n37310);
  nand U39612(n37310,n37382,n37383,n37384,n37385);
  nor U39613(n37385,n37386,n37387);
  nor U39614(n37387,n36302,n37363);
  nor U39615(n37386,n35191,n36246);
  nand U39616(n37384,n36271,G60225);
  nand U39617(n37383,n35193,n37388);
  nand U39618(n37388,n37389,n37390);
  nand U39619(n37390,n36305,n37391);
  nand U39620(n37382,n37302,n35203,n37392);
  xnor U39621(n37381,n36246,n37309);
  nand U39622(n37309,n37393,n37394);
  nand U39623(n37394,n36238,n37395);
  or U39624(n37395,n37396,n37397);
  nand U39625(n37393,n37397,n37396);
  nand U39626(n37372,n36272,n35193);
  not U39627(n35193,n37392);
  xnor U39628(n37392,n37370,n37398);
  and U39629(n37398,n37371,n37368);
  nand U39630(n37368,n37399,n37400,n36390);
  nand U39631(n37399,n37401,n37402);
  nand U39632(n37371,n37401,n37402,n37403);
  nand U39633(n37402,n36267,n35191,n37404);
  nand U39634(n37401,n37405,n36215);
  nand U39635(n37405,n37404,n37406);
  nand U39636(n37406,n35472,n36329);
  not U39637(n35472,n35191);
  xnor U39638(n35191,n37323,n37322);
  xor U39639(n37322,n34962,n37407);
  nor U39640(n37407,n37408,n37409,n37410);
  and U39641(n37410,n36269,G60161);
  nor U39642(n37409,n36527,n37363);
  not U39643(n37363,G60034);
  nand U39644(n37408,n37411,n37412,n37413);
  nand U39645(n37413,G60066,n36267);
  nand U39646(n37412,n35545,n37380);
  nand U39647(n37380,n37414,n37415,n37416);
  or U39648(n37416,n37364,G60034);
  nand U39649(n37415,G60034,n37364,n34912);
  nand U39650(n37364,n37417,n37418);
  nand U39651(n37414,n36803,n35692);
  nand U39652(n36803,n37419,n37420,n37421,n37422);
  nor U39653(n37422,n37423,n37424,n37425,n37426);
  nor U39654(n37426,n36799,n37003);
  nor U39655(n37425,n36800,n37005);
  nor U39656(n37424,n36801,n37007);
  nor U39657(n37423,n36802,n37009);
  nor U39658(n37421,n37427,n37428,n37429,n37430);
  nor U39659(n37430,n36791,n37015);
  nor U39660(n37429,n36792,n37017);
  nor U39661(n37428,n36793,n37019);
  nor U39662(n37427,n36794,n37021);
  nor U39663(n37420,n37431,n37432,n37433,n37434);
  nor U39664(n37434,n36783,n37026);
  nor U39665(n37433,n36784,n37027);
  nor U39666(n37432,n36785,n37028);
  nor U39667(n37431,n36786,n37029);
  nor U39668(n37419,n37435,n37436,n37437,n37438);
  nor U39669(n37438,n36775,n37034);
  nor U39670(n37437,n36776,n37035);
  nor U39671(n37436,n36777,n37036);
  nor U39672(n37435,n36778,n37037);
  nand U39673(n37411,G60193,n36266);
  and U39674(n37404,n37439,n37440,n37441);
  nand U39675(n37441,G60066,n37121);
  nand U39676(n37440,G60034,n36328);
  nand U39677(n37439,G60225,n34962);
  nand U39678(n37370,n37442,n37443);
  nand U39679(n37443,n37444,n37445);
  nand U39680(G14524,n37446,n37447,n37448,n37449);
  nor U39681(n37449,n37450,n37451,n37452);
  nor U39682(n37452,n37453,n36233);
  not U39683(n37453,G60224);
  and U39684(n37451,n37454,n36729);
  nor U39685(n37450,n37455,n36288);
  nand U39686(n37448,n36234,n35476);
  nand U39687(n37447,n36235,n35202);
  xor U39688(n35202,n37456,n37397);
  nand U39689(n37397,n37457,n37458,n37459,n37460);
  nor U39690(n37460,n37461,n37462);
  nor U39691(n37462,n36302,n37455);
  nor U39692(n37461,n35201,n36246);
  nand U39693(n37459,n36271,G60224);
  nand U39694(n37458,n37302,n37391);
  nor U39695(n37302,n37463,n37464,n35781);
  or U39696(n37457,n37391,n37389);
  nor U39697(n37389,n37465,n37466);
  nor U39698(n37466,n35213,n35781);
  xnor U39699(n37456,n36246,n37396);
  nand U39700(n37396,n37467,n37468);
  nand U39701(n37468,n36238,n37469);
  or U39702(n37469,n37470,n37471);
  nand U39703(n37467,n37471,n37470);
  nand U39704(n37446,n36272,n35203);
  not U39705(n35203,n37391);
  xnor U39706(n37391,n37444,n37472);
  and U39707(n37472,n37445,n37442);
  nand U39708(n37442,n37473,n37474,n36390);
  nand U39709(n37473,n37475,n37476);
  nand U39710(n37445,n37475,n37476,n37477);
  nand U39711(n37476,n36267,n35201,n37478);
  nand U39712(n37475,n37479,n36215);
  nand U39713(n37479,n37478,n37480);
  nand U39714(n37480,n35476,n36329);
  not U39715(n35476,n35201);
  nand U39716(n35201,n37323,n37481);
  nand U39717(n37481,n37482,n37483);
  or U39718(n37323,n37483,n37482);
  xor U39719(n37482,n34962,n37484);
  nor U39720(n37484,n37485,n37486,n37487);
  and U39721(n37487,n36269,G60160);
  nor U39722(n37486,n36527,n37455);
  nand U39723(n37485,n37488,n37489,n37490);
  nand U39724(n37490,G60065,n36267);
  nand U39725(n37489,n35545,n37454);
  nand U39726(n37454,n37491,n37492);
  nand U39727(n37492,n36901,n35692);
  nand U39728(n36901,n37493,n37494,n37495,n37496);
  nor U39729(n37496,n37497,n37498,n37499,n37500);
  nor U39730(n37500,n36895,n37003);
  nor U39731(n37499,n36896,n37005);
  nor U39732(n37498,n36897,n37007);
  nor U39733(n37497,n36898,n37009);
  nor U39734(n37495,n37501,n37502,n37503,n37504);
  nor U39735(n37504,n36887,n37015);
  nor U39736(n37503,n36888,n37017);
  nor U39737(n37502,n36889,n37019);
  nor U39738(n37501,n36890,n37021);
  nor U39739(n37494,n37505,n37506,n37507,n37508);
  nor U39740(n37508,n36879,n37026);
  nor U39741(n37507,n36880,n37027);
  nor U39742(n37506,n36881,n37028);
  nor U39743(n37505,n36882,n37029);
  nor U39744(n37493,n37509,n37510,n37511,n37512);
  nor U39745(n37512,n36871,n37034);
  nor U39746(n37511,n36872,n37035);
  nor U39747(n37510,n36873,n37036);
  nor U39748(n37509,n36874,n37037);
  xnor U39749(n37491,n37417,n37418);
  nor U39750(n37418,n37455,n35692);
  not U39751(n37455,G60033);
  nor U39752(n37417,n37513,n37514);
  nand U39753(n37488,G60192,n36266);
  and U39754(n37478,n37515,n37516,n37517);
  nand U39755(n37517,G60065,n37121);
  nand U39756(n37516,G60033,n36328);
  nand U39757(n37515,G60224,n34962);
  nand U39758(n37444,n37518,n37519);
  nand U39759(n37519,n37520,n37521);
  not U39760(n37520,n37522);
  nand U39761(G14523,n37523,n37524,n37525,n37526);
  nor U39762(n37526,n37527,n37528,n37529);
  nor U39763(n37529,n37530,n36233);
  not U39764(n37530,G60223);
  and U39765(n37528,n37531,n36729);
  nor U39766(n37527,n37514,n36288);
  nand U39767(n37525,n36234,n35480);
  nand U39768(n37524,n36235,n35212);
  xor U39769(n35212,n37532,n37471);
  nand U39770(n37471,n37533,n37534);
  nand U39771(n37534,n36238,n37535);
  or U39772(n37535,n37536,n37537);
  nand U39773(n37533,n37537,n37536);
  xnor U39774(n37532,n37470,n36246);
  nand U39775(n37470,n37538,n37539,n37540,n37541);
  nor U39776(n37541,n37542,n37543);
  nor U39777(n37543,n36302,n37514);
  nor U39778(n37542,n35211,n36246);
  nand U39779(n37540,n36271,G60223);
  nand U39780(n37539,n35213,n37465);
  nand U39781(n37465,n36582,n37544);
  nand U39782(n37544,n37464,n36305);
  not U39783(n37464,n37304);
  nand U39784(n37538,n36305,n37304,n37463);
  not U39785(n37463,n35213);
  nand U39786(n37304,n37545,n37546);
  nand U39787(n37546,n37547,n37548);
  or U39788(n37547,n37549,n35223);
  nand U39789(n37545,n35223,n37549);
  nand U39790(n37523,n36272,n35213);
  xor U39791(n35213,n37550,n37522);
  nand U39792(n37550,n37518,n37521);
  nand U39793(n37521,n37551,n37552,n37553);
  nand U39794(n37518,n37555,n37554,n36390);
  nand U39795(n37555,n37551,n37552);
  nand U39796(n37552,n36267,n35211,n37556);
  nand U39797(n37551,n37557,n36215);
  nand U39798(n37557,n37556,n37558);
  nand U39799(n37558,n35480,n36329);
  not U39800(n35480,n35211);
  nand U39801(n35211,n37483,n37559);
  nand U39802(n37559,n37560,n37561);
  or U39803(n37483,n37561,n37560);
  and U39804(n37560,n37562,n37563);
  nand U39805(n37563,n37564,n37565);
  xor U39806(n37561,n34962,n37566);
  nor U39807(n37566,n37567,n37568,n37569);
  and U39808(n37569,n36269,G60159);
  nor U39809(n37568,n36527,n37514);
  nand U39810(n37567,n37570,n37571,n37572);
  nand U39811(n37572,G60064,n36267);
  nand U39812(n37571,n35545,n37531);
  nand U39813(n37531,n37573,n37574,n37575);
  nand U39814(n37575,n37576,n37514);
  not U39815(n37514,G60032);
  nand U39816(n37574,G60032,n37513,n34912);
  not U39817(n37513,n37576);
  nor U39818(n37576,n37577,n37578,n37579);
  nand U39819(n37573,n37038,n35692);
  nand U39820(n37038,n37580,n37581,n37582,n37583);
  nor U39821(n37583,n37584,n37585,n37586,n37587);
  nor U39822(n37587,n36983,n37003);
  nor U39823(n37586,n36987,n37005);
  nor U39824(n37585,n36988,n37007);
  nor U39825(n37584,n36990,n37009);
  nor U39826(n37582,n37588,n37589,n37590,n37591);
  nor U39827(n37591,n36974,n37015);
  nor U39828(n37590,n36976,n37017);
  nor U39829(n37589,n36977,n37019);
  nor U39830(n37588,n36978,n37021);
  nor U39831(n37581,n37592,n37593,n37594,n37595);
  nor U39832(n37595,n36964,n37026);
  nor U39833(n37594,n36966,n37027);
  nor U39834(n37593,n36967,n37028);
  nor U39835(n37592,n36968,n37029);
  nor U39836(n37580,n37596,n37597,n37598,n37599);
  nor U39837(n37599,n36949,n37034);
  nor U39838(n37598,n36952,n37035);
  nor U39839(n37597,n36954,n37036);
  nor U39840(n37596,n36956,n37037);
  nand U39841(n37570,G60191,n36266);
  and U39842(n37556,n37600,n37601,n37602);
  nand U39843(n37602,G60064,n37121);
  nand U39844(n37601,G60032,n36328);
  nand U39845(n37600,G60223,n34962);
  nand U39846(G14522,n37603,n37604,n37605,n37606);
  nor U39847(n37606,n37607,n37608,n37609);
  nor U39848(n37609,G60031,n36226,n37610,n37579);
  nor U39849(n37608,n37611,n37578);
  nor U39850(n37611,n37612,n36231);
  nor U39851(n37612,n37613,n36226);
  nor U39852(n37613,n37610,n37579);
  nor U39853(n37607,n37614,n36233);
  nand U39854(n37605,n36234,n35484);
  nand U39855(n37604,n36235,n35222);
  xor U39856(n35222,n37615,n37537);
  nand U39857(n37537,n37616,n37617,n37618,n37619);
  nor U39858(n37619,n37620,n37621);
  nor U39859(n37621,n37614,n36301);
  not U39860(n37614,G60222);
  nor U39861(n37620,n36302,n37578);
  not U39862(n37578,G60031);
  nand U39863(n37618,n36238,n35484);
  nand U39864(n37617,n36305,n37622);
  xor U39865(n37622,n37549,n37623);
  xor U39866(n37623,n35223,n37548);
  nand U39867(n37549,n37624,n37625);
  nand U39868(n37625,n37626,n37627);
  nand U39869(n37626,n37628,n37629);
  or U39870(n37624,n37628,n37629);
  nand U39871(n37616,n35223,n36255);
  xnor U39872(n37615,n36246,n37536);
  nand U39873(n37536,n37630,n37631);
  nand U39874(n37631,n36238,n37632);
  or U39875(n37632,n37633,n37634);
  nand U39876(n37630,n37634,n37633);
  nand U39877(n37603,n36272,n35223);
  and U39878(n35223,n37522,n37635);
  nand U39879(n37635,n37636,n37637);
  xnor U39880(n37636,n36267,n37638);
  nand U39881(n37522,n37639,n37640);
  xnor U39882(n37639,n37638,n36215);
  nand U39883(n37638,n37641,n37642,n37643,n37644);
  nand U39884(n37644,n35484,n36329);
  not U39885(n35484,n35221);
  xor U39886(n35221,n37645,n37564);
  nand U39887(n37564,n37646,n37647);
  nand U39888(n37647,n37648,n37649);
  nand U39889(n37645,n37565,n37562);
  nand U39890(n37562,n37650,n37548,n35545);
  nand U39891(n37565,n37651,n37652,n37653);
  nand U39892(n37653,n35545,n37548);
  nand U39893(n37548,n37654,n37655,n37656,n37657);
  nor U39894(n37657,n37658,n37659,n37660,n37661);
  nor U39895(n37661,n37006,n37662);
  nor U39896(n37660,n37004,n37663);
  nor U39897(n37659,n37002,n37664);
  nor U39898(n37658,n37018,n37665);
  nor U39899(n37656,n37666,n37667,n37668,n37669);
  nor U39900(n37669,n37016,n37670);
  nor U39901(n37668,n37014,n37671);
  nor U39902(n37667,n36386,n37672);
  nor U39903(n37666,n36384,n37673);
  nor U39904(n37655,n37674,n37675,n37676,n37677);
  nor U39905(n37677,n36382,n37678);
  nor U39906(n37676,n36374,n37679);
  nor U39907(n37675,n36372,n37680);
  nor U39908(n37674,n36370,n37681);
  nor U39909(n37654,n37682,n37683,n37684,n37685);
  nor U39910(n37685,n37008,n37686);
  nor U39911(n37684,n37020,n37687);
  nor U39912(n37683,n36388,n37688);
  nor U39913(n37682,n36376,n37689);
  nand U39914(n37652,n37690,n34962);
  nand U39915(n37651,n37650,n35998);
  nand U39916(n37650,n37691,n37692,n37690);
  and U39917(n37690,n37693,n37694);
  nand U39918(n37694,G60190,n36266);
  nand U39919(n37693,G60063,n36267);
  nand U39920(n37692,G60031,n36268);
  nand U39921(n37691,G60158,n36269);
  nand U39922(n37643,G60031,n36328);
  nand U39923(n37642,G60222,n34962);
  nand U39924(n37641,G60063,n37121);
  nand U39925(G14521,n37695,n37696,n37697,n37698);
  nor U39926(n37698,n37699,n37700,n37701);
  nor U39927(n37701,n35231,n36726);
  nor U39928(n37700,n37628,n37702);
  nor U39929(n37699,n37703,n36233);
  nand U39930(n37697,n36235,n35232);
  xor U39931(n35232,n37704,n37634);
  nand U39932(n37634,n37705,n37706,n37707,n37708);
  nor U39933(n37708,n37709,n37710);
  nor U39934(n37710,n37703,n36301);
  not U39935(n37703,G60221);
  nor U39936(n37709,n36302,n37610);
  not U39937(n37610,G60030);
  nand U39938(n37707,n36238,n35488);
  nand U39939(n37706,n37711,n36305);
  xor U39940(n37711,n37629,n37712);
  xnor U39941(n37712,n37627,n35233);
  nand U39942(n37629,n37713,n37714);
  nand U39943(n37714,n37715,n37716);
  or U39944(n37716,n37717,n37718);
  nand U39945(n37713,n37718,n37717);
  nand U39946(n37705,n35233,n36255);
  not U39947(n35233,n37628);
  nand U39948(n37628,n37637,n37719);
  nand U39949(n37719,n37720,n37721);
  not U39950(n37637,n37640);
  nor U39951(n37640,n37721,n37720);
  xor U39952(n37720,n37722,n36215);
  nand U39953(n37722,n37723,n37724,n37725,n37726);
  nand U39954(n37726,n35488,n36329);
  not U39955(n35488,n35231);
  xor U39956(n35231,n37727,n37649);
  nand U39957(n37649,n37728,n37729);
  nand U39958(n37729,n37730,n37731);
  nand U39959(n37727,n37646,n37648);
  nand U39960(n37648,n37732,n37733);
  nand U39961(n37733,n35545,n37627);
  xnor U39962(n37732,n34962,n37734);
  nand U39963(n37646,n37734,n37627,n35545);
  nand U39964(n37627,n37735,n37736,n37737,n37738);
  nor U39965(n37738,n37739,n37740,n37741,n37742);
  nor U39966(n37742,n36479,n37662);
  nor U39967(n37741,n36477,n37663);
  nor U39968(n37740,n36475,n37664);
  nor U39969(n37739,n36467,n37665);
  nor U39970(n37737,n37743,n37744,n37745,n37746);
  nor U39971(n37746,n36465,n37670);
  nor U39972(n37745,n36463,n37671);
  nor U39973(n37744,n36457,n37672);
  nor U39974(n37743,n36456,n37673);
  nor U39975(n37736,n37747,n37748,n37749,n37750);
  nor U39976(n37750,n36455,n37678);
  nor U39977(n37749,n36449,n37679);
  nor U39978(n37748,n36448,n37680);
  nor U39979(n37747,n36447,n37681);
  nor U39980(n37735,n37751,n37752,n37753,n37754);
  nor U39981(n37754,n36481,n37686);
  nor U39982(n37753,n36469,n37687);
  nor U39983(n37752,n36458,n37688);
  nor U39984(n37751,n36450,n37689);
  nand U39985(n37734,n37755,n37756,n37757,n37758);
  nand U39986(n37758,G60189,n36266);
  nand U39987(n37757,G60062,n36267);
  nand U39988(n37756,G60030,n36268);
  nand U39989(n37755,G60157,n36269);
  nand U39990(n37725,G60030,n36328);
  nand U39991(n37724,G60221,n34962);
  nand U39992(n37723,G60062,n37121);
  xnor U39993(n37704,n36246,n37633);
  nand U39994(n37633,n37759,n37760);
  nand U39995(n37760,n36238,n37761);
  nand U39996(n37761,n37762,n37763);
  or U39997(n37759,n37763,n37762);
  nand U39998(n37696,n37764,n37577,n36729);
  nand U39999(n37577,G60030,n34912);
  nand U40000(n37695,G60030,n37765);
  nand U40001(n37765,n36288,n37766);
  nand U40002(n37766,n36729,n37579);
  not U40003(n37579,n37764);
  nor U40004(n37764,n37767,n37768,n37769);
  nand U40005(G14520,n37770,n37771,n37772,n37773);
  nor U40006(n37773,n37774,n37775,n37776);
  nor U40007(n37776,G60029,n36226,n37777,n37769);
  nor U40008(n37775,n37778,n37768);
  nor U40009(n37778,n37779,n37780);
  nor U40010(n37779,G60028,n36226);
  nor U40011(n37774,n37781,n36233);
  nand U40012(n37772,n36234,n35492);
  nand U40013(n37771,n36235,n35242);
  xnor U40014(n35242,n37762,n37782);
  xnor U40015(n37782,n36238,n37763);
  nand U40016(n37763,n37783,n37784);
  nand U40017(n37784,n37785,n36246);
  nand U40018(n37785,n37786,n37787);
  or U40019(n37783,n37786,n37787);
  and U40020(n37762,n37788,n37789,n37790,n37791);
  nor U40021(n37791,n37792,n37793);
  nor U40022(n37793,n37781,n36301);
  not U40023(n37781,G60220);
  nor U40024(n37792,n36302,n37768);
  not U40025(n37768,G60029);
  nand U40026(n37790,n36238,n35492);
  nand U40027(n37789,n37794,n36305);
  xor U40028(n37794,n37718,n37795);
  xnor U40029(n37795,n37715,n37717);
  not U40030(n37715,n37796);
  nand U40031(n37718,n37797,n37798);
  nand U40032(n37798,n37799,n37800);
  or U40033(n37800,n37801,n37802);
  not U40034(n37799,n37803);
  nand U40035(n37797,n37802,n37801);
  nand U40036(n37788,n35243,n36255);
  nand U40037(n37770,n36272,n35243);
  not U40038(n35243,n37717);
  nand U40039(n37717,n37721,n37804);
  nand U40040(n37804,n37805,n37806);
  or U40041(n37721,n37806,n37805);
  xor U40042(n37805,n37807,n36215);
  nand U40043(n37807,n37808,n37809,n37810,n37811);
  nand U40044(n37811,n35492,n36329);
  not U40045(n35492,n35241);
  xor U40046(n35241,n37812,n37730);
  or U40047(n37730,n37813,n37814);
  nor U40048(n37814,n37815,n37816);
  nand U40049(n37812,n37731,n37728);
  nand U40050(n37728,n37817,n37796,n35545);
  nand U40051(n37731,n37818,n37819,n37820);
  nand U40052(n37820,n35545,n37796);
  nand U40053(n37796,n37821,n37822,n37823,n37824);
  nor U40054(n37824,n37825,n37826,n37827,n37828);
  nor U40055(n37828,n37179,n37662);
  nor U40056(n37827,n37178,n37663);
  nor U40057(n37826,n37177,n37664);
  nor U40058(n37825,n37187,n37665);
  nor U40059(n37823,n37829,n37830,n37831,n37832);
  nor U40060(n37832,n37186,n37670);
  nor U40061(n37831,n37185,n37671);
  nor U40062(n37830,n36561,n37672);
  nor U40063(n37829,n36560,n37673);
  nor U40064(n37822,n37833,n37834,n37835,n37836);
  nor U40065(n37836,n36559,n37678);
  nor U40066(n37835,n36553,n37679);
  nor U40067(n37834,n36552,n37680);
  nor U40068(n37833,n36551,n37681);
  nor U40069(n37821,n37837,n37838,n37839,n37840);
  nor U40070(n37840,n37180,n37686);
  nor U40071(n37839,n37188,n37687);
  nor U40072(n37838,n36562,n37688);
  nor U40073(n37837,n36554,n37689);
  nand U40074(n37819,n37841,n34962);
  nand U40075(n37818,n37817,n35998);
  nand U40076(n37817,n37842,n37843,n37841);
  and U40077(n37841,n37844,n37845);
  nand U40078(n37845,G60188,n36266);
  nand U40079(n37844,G60061,n36267);
  nand U40080(n37843,G60029,n36268);
  nand U40081(n37842,G60156,n36269);
  nand U40082(n37810,G60029,n36328);
  nand U40083(n37809,G60220,n34962);
  nand U40084(n37808,G60061,n37121);
  nand U40085(n37806,n37846,n37847);
  nand U40086(G14519,n37848,n37849,n37850,n37851);
  nor U40087(n37851,n37852,n37853,n37854);
  nor U40088(n37854,n35251,n36726);
  not U40089(n35251,n35496);
  nor U40090(n37853,n37802,n37702);
  nor U40091(n37852,n37855,n36233);
  nand U40092(n37850,n36235,n35252);
  xnor U40093(n35252,n37787,n37856);
  xnor U40094(n37856,n36238,n37786);
  nand U40095(n37786,n37857,n37858,n37859,n37860);
  nor U40096(n37860,n37861,n37862);
  nor U40097(n37862,n37855,n36301);
  not U40098(n37855,G60219);
  nor U40099(n37861,n36302,n37777);
  not U40100(n37777,G60028);
  nand U40101(n37859,n36238,n35496);
  nand U40102(n37858,n36305,n37863);
  xnor U40103(n37863,n37802,n37864);
  xnor U40104(n37864,n37801,n37803);
  nand U40105(n37801,n37865,n37866);
  nand U40106(n37866,n37867,n37868);
  or U40107(n37868,n37869,n37870);
  not U40108(n37867,n37871);
  nand U40109(n37865,n37870,n37869);
  nand U40110(n37857,n35253,n36255);
  not U40111(n35253,n37802);
  xnor U40112(n37802,n37847,n37846);
  xnor U40113(n37847,n37872,n36215);
  nand U40114(n37872,n37873,n37874,n37875,n37876);
  nand U40115(n37876,n35496,n36329);
  xnor U40116(n35496,n37815,n37877);
  nor U40117(n37877,n37813,n37816);
  and U40118(n37816,n37878,n37879,n37880);
  nand U40119(n37880,n37881,n34962);
  nor U40120(n37813,n37879,n37878);
  nand U40121(n37878,n35545,n37803);
  nand U40122(n37803,n37882,n37883,n37884,n37885);
  nor U40123(n37885,n37886,n37887,n37888,n37889);
  nor U40124(n37889,n36631,n37680);
  nor U40125(n37888,n36632,n37679);
  nor U40126(n37887,n36640,n37672);
  nor U40127(n37886,n37269,n37665);
  nor U40128(n37884,n37890,n37891,n37892,n37893);
  nor U40129(n37893,n36639,n37673);
  nor U40130(n37892,n36641,n37688);
  nor U40131(n37891,n37262,n37686);
  nor U40132(n37890,n36630,n37681);
  nor U40133(n37883,n37894,n37895,n37896,n37897);
  nor U40134(n37897,n37268,n37670);
  nor U40135(n37896,n37270,n37687);
  nor U40136(n37895,n37259,n37664);
  nor U40137(n37894,n36638,n37678);
  nor U40138(n37882,n37898,n37899,n37900,n37901);
  nor U40139(n37901,n37260,n37663);
  nor U40140(n37900,n37267,n37671);
  nor U40141(n37899,n36633,n37689);
  nor U40142(n37898,n37261,n37662);
  nand U40143(n37879,n37902,n35998);
  nand U40144(n37902,n37903,n37904,n37881);
  and U40145(n37881,n37905,n37906);
  nand U40146(n37906,G60187,n36266);
  nand U40147(n37905,G60060,n36267);
  nand U40148(n37904,G60028,n36268);
  nand U40149(n37903,G60155,n36269);
  nand U40150(n37815,n37907,n37908);
  nand U40151(n37908,n37909,n37910,n37911);
  nand U40152(n37875,G60028,n36328);
  nand U40153(n37874,G60219,n34962);
  nand U40154(n37873,G60060,n37121);
  nand U40155(n37787,n37912,n37913,n37914);
  or U40156(n37914,n36246,n37915);
  nor U40157(n37915,n37916,n37917,n37918);
  nand U40158(n37912,n37918,n37919,n37917);
  nand U40159(n37849,n37920,n37767,n36729);
  nand U40160(n37767,G60028,n34912);
  not U40161(n37920,n37769);
  nand U40162(n37848,G60028,n37780);
  nand U40163(n37780,n36288,n37921);
  nand U40164(n37921,n36729,n37769);
  nand U40165(n37769,n37922,G60027);
  nand U40166(G14518,n37923,n37924,n37925,n37926);
  nor U40167(n37926,n37927,n37928,n37929);
  and U40168(n37929,n37930,n37922,n36729);
  nor U40169(n37928,n37931,n37930);
  nor U40170(n37931,n37932,n36231);
  nor U40171(n37932,n37922,n36226);
  nor U40172(n37922,n37933,n37934,n37935);
  nor U40173(n37927,n37936,n36233);
  nand U40174(n37925,n36234,n35500);
  nand U40175(n37924,n36235,n35262);
  xnor U40176(n35262,n37937,n37938);
  nor U40177(n37938,n37916,n37939);
  not U40178(n37916,n37940);
  xnor U40179(n37937,n37918,n36246);
  nand U40180(n37918,n37941,n37942,n37943,n37944);
  nor U40181(n37944,n37945,n37946);
  nor U40182(n37946,n37936,n36301);
  not U40183(n37936,G60218);
  nor U40184(n37945,n36302,n37930);
  not U40185(n37930,G60027);
  nand U40186(n37943,n36238,n35500);
  nand U40187(n37942,n37947,n36305);
  xnor U40188(n37947,n37948,n37870);
  not U40189(n37870,n35263);
  xnor U40190(n37948,n37869,n37871);
  nand U40191(n37869,n37949,n37950);
  nand U40192(n37950,n37951,n37952);
  nand U40193(n37952,n35276,n37953);
  nand U40194(n37949,n37954,n36144);
  nand U40195(n37941,n35263,n36255);
  nand U40196(n37923,n36272,n35263);
  nor U40197(n35263,n37846,n37955);
  and U40198(n37955,n37956,n37957);
  nor U40199(n37846,n37957,n37956);
  xor U40200(n37956,n37958,n36215);
  nand U40201(n37958,n37959,n37960,n37961,n37962);
  nand U40202(n37962,n35500,n36329);
  not U40203(n35500,n35261);
  xnor U40204(n35261,n37963,n37964);
  and U40205(n37964,n37911,n37907);
  nand U40206(n37907,n37965,n37966,n37967);
  nand U40207(n37967,n35545,n37871);
  nand U40208(n37966,n37968,n35998);
  nand U40209(n37965,n37969,n34962);
  nand U40210(n37911,n37968,n37871,n35545);
  nand U40211(n37871,n37970,n37971,n37972,n37973);
  nor U40212(n37973,n37974,n37975,n37976,n37977);
  nor U40213(n37977,n36707,n37680);
  nor U40214(n37976,n36708,n37679);
  nor U40215(n37975,n36716,n37672);
  nor U40216(n37974,n37352,n37665);
  nor U40217(n37972,n37978,n37979,n37980,n37981);
  nor U40218(n37981,n36715,n37673);
  nor U40219(n37980,n36717,n37688);
  nor U40220(n37979,n37345,n37686);
  nor U40221(n37978,n36706,n37681);
  nor U40222(n37971,n37982,n37983,n37984,n37985);
  nor U40223(n37985,n37351,n37670);
  nor U40224(n37984,n37353,n37687);
  nor U40225(n37983,n37342,n37664);
  nor U40226(n37982,n36714,n37678);
  nor U40227(n37970,n37986,n37987,n37988,n37989);
  nor U40228(n37989,n37343,n37663);
  nor U40229(n37988,n37350,n37671);
  nor U40230(n37987,n36709,n37689);
  nor U40231(n37986,n37344,n37662);
  nand U40232(n37968,n37990,n37991,n37969);
  and U40233(n37969,n37992,n37993);
  nand U40234(n37993,G60186,n36266);
  nand U40235(n37992,G60059,n36267);
  nand U40236(n37991,G60027,n36268);
  nand U40237(n37990,G60154,n36269);
  nand U40238(n37963,n37910,n37909);
  nand U40239(n37961,G60027,n36328);
  nand U40240(n37960,G60218,n34962);
  nand U40241(n37959,G60059,n37121);
  nand U40242(G14517,n37994,n37995,n37996,n37997);
  nor U40243(n37997,n37998,n37999,n38000);
  nor U40244(n38000,G60026,n36226,n37933,n37935);
  nor U40245(n37999,n38001,n37934);
  nor U40246(n38001,n38002,n38003);
  nor U40247(n38002,G60025,n36226);
  nor U40248(n37998,n36146,n36233);
  nand U40249(n37996,n36234,n35504);
  nand U40250(n37995,n36235,n35727);
  not U40251(n35727,n35275);
  nand U40252(n35275,n38004,n38005);
  nand U40253(n38005,n38006,n37913,n38007);
  nand U40254(n38007,n38008,n37940);
  nand U40255(n38004,n37940,n37939);
  nand U40256(n37939,n37913,n38009);
  nand U40257(n38009,n37917,n38008);
  or U40258(n38008,n37919,n36238);
  not U40259(n37917,n38006);
  nand U40260(n38006,n38010,n38011);
  nand U40261(n38011,n38012,n36246);
  nand U40262(n37940,n36238,n37919);
  nand U40263(n37919,n38013,n38014,n38015,n38016);
  nor U40264(n38016,n38017,n38018);
  nor U40265(n38018,n36146,n36301);
  not U40266(n36146,G60217);
  nor U40267(n38017,n36302,n37934);
  nand U40268(n38015,n36238,n35504);
  nand U40269(n38014,n36305,n38019);
  xnor U40270(n38019,n35276,n38020);
  xnor U40271(n38020,n37951,n37954);
  and U40272(n37951,n38021,n38022);
  nand U40273(n38022,n38023,n38024,n35296);
  nand U40274(n38013,n35276,n36255);
  nand U40275(n37994,n36272,n35276);
  not U40276(n35276,n36144);
  nand U40277(n36144,n38025,n37957);
  nand U40278(n37957,n38026,n38027,n38028);
  xnor U40279(n38028,n38029,n36215);
  nand U40280(n38025,n38030,n38031);
  nand U40281(n38031,n38027,n38026);
  xnor U40282(n38030,n36267,n38029);
  nand U40283(n38029,n38032,n38033,n38034,n38035);
  nand U40284(n38035,n35504,n36329);
  not U40285(n35504,n35271);
  nand U40286(n35271,n38036,n38037);
  or U40287(n38037,n37909,n38038);
  nand U40288(n37909,n38039,n38040);
  nand U40289(n38040,n38041,n38042);
  nand U40290(n38036,n38043,n38042,n38041);
  nand U40291(n38041,n38044,n38045);
  nand U40292(n38043,n38039,n37910);
  not U40293(n37910,n38038);
  nor U40294(n38038,n34968,n37954,n38046);
  not U40295(n37954,n37953);
  nand U40296(n38039,n38046,n38047);
  nand U40297(n38047,n35545,n37953);
  nand U40298(n37953,n38048,n38049,n38050,n38051);
  nor U40299(n38051,n38052,n38053,n38054,n38055);
  nor U40300(n38055,n36801,n37662);
  nor U40301(n38054,n36800,n37663);
  nor U40302(n38053,n36799,n37664);
  nor U40303(n38052,n36793,n37665);
  nor U40304(n38050,n38056,n38057,n38058,n38059);
  nor U40305(n38059,n36792,n37670);
  nor U40306(n38058,n36791,n37671);
  nor U40307(n38057,n36785,n37672);
  nor U40308(n38056,n36784,n37673);
  nor U40309(n38049,n38060,n38061,n38062,n38063);
  nor U40310(n38063,n36783,n37678);
  nor U40311(n38062,n36777,n37679);
  nor U40312(n38061,n36776,n37680);
  nor U40313(n38060,n36775,n37681);
  nor U40314(n38048,n38064,n38065,n38066,n38067);
  nor U40315(n38067,n36802,n37686);
  nor U40316(n38066,n36794,n37687);
  nor U40317(n38065,n36786,n37688);
  nor U40318(n38064,n36778,n37689);
  xor U40319(n38046,n34962,n38068);
  nor U40320(n38068,n38069,n38070,n38071,n38072);
  and U40321(n38072,n36269,G60153);
  nor U40322(n38071,n36527,n37934);
  not U40323(n37934,G60026);
  and U40324(n38070,n36267,G60058);
  nor U40325(n38069,n38073,n35272);
  not U40326(n35272,G60185);
  nand U40327(n38034,G60026,n36328);
  nand U40328(n38033,G60217,n34962);
  nand U40329(n38032,G60058,n37121);
  nand U40330(G14516,n38074,n38075,n38076,n38077);
  nor U40331(n38077,n38078,n38079,n38080);
  nor U40332(n38080,G60025,n37935,n36226);
  and U40333(n38079,n38003,G60025);
  nand U40334(n38003,n36288,n38081);
  nand U40335(n38081,n36729,n37935);
  nand U40336(n37935,G60024,G60023,n38082);
  nor U40337(n38078,n38083,n36233);
  nand U40338(n38076,n36234,n35508);
  nand U40339(n38075,n36235,n35285);
  nand U40340(n35285,n38084,n38085,n38086);
  or U40341(n38086,n37913,n38087);
  nand U40342(n37913,n36238,n38088);
  nand U40343(n38085,n38087,n38012,n36238);
  not U40344(n38012,n38088);
  nand U40345(n38084,n38089,n36246);
  xnor U40346(n38089,n38088,n38087);
  not U40347(n38087,n38010);
  nand U40348(n38010,n38090,n38091);
  nand U40349(n38091,n36238,n38092);
  or U40350(n38092,n38093,n38094);
  nand U40351(n38090,n38094,n38093);
  nand U40352(n38088,n38095,n38096,n38097,n38098);
  nor U40353(n38098,n38099,n38100);
  nor U40354(n38100,n38083,n36301);
  not U40355(n38083,G60216);
  nor U40356(n38099,n36302,n37933);
  not U40357(n37933,G60025);
  nand U40358(n38097,n36238,n35508);
  nand U40359(n38096,n36305,n38101);
  xor U40360(n38101,n38102,n38103);
  nand U40361(n38103,n35296,n38024);
  nand U40362(n38102,n38023,n38021);
  nand U40363(n38021,n35286,n38104);
  or U40364(n38023,n38104,n35286);
  nand U40365(n38095,n35286,n36255);
  nand U40366(n38074,n36272,n35286);
  xor U40367(n35286,n38027,n38026);
  xor U40368(n38026,n38105,n36267);
  nand U40369(n38105,n38106,n38107,n38108,n38109);
  nand U40370(n38109,n35508,n36329);
  not U40371(n35508,n35284);
  xnor U40372(n35284,n38045,n38110);
  and U40373(n38110,n38044,n38042);
  nand U40374(n38042,n38111,n38104,n35545);
  nand U40375(n38044,n38112,n38113,n38114);
  nand U40376(n38114,n35545,n38104);
  nand U40377(n38104,n38115,n38116,n38117,n38118);
  nor U40378(n38118,n38119,n38120,n38121,n38122);
  nor U40379(n38122,n36897,n37662);
  nor U40380(n38121,n36896,n37663);
  nor U40381(n38120,n36895,n37664);
  nor U40382(n38119,n36889,n37665);
  nor U40383(n38117,n38123,n38124,n38125,n38126);
  nor U40384(n38126,n36888,n37670);
  nor U40385(n38125,n36887,n37671);
  nor U40386(n38124,n36881,n37672);
  nor U40387(n38123,n36880,n37673);
  nor U40388(n38116,n38127,n38128,n38129,n38130);
  nor U40389(n38130,n36879,n37678);
  nor U40390(n38129,n36873,n37679);
  nor U40391(n38128,n36872,n37680);
  nor U40392(n38127,n36871,n37681);
  nor U40393(n38115,n38131,n38132,n38133,n38134);
  nor U40394(n38134,n36898,n37686);
  nor U40395(n38133,n36890,n37687);
  nor U40396(n38132,n36882,n37688);
  nor U40397(n38131,n36874,n37689);
  nand U40398(n38113,n38111,n35998);
  nand U40399(n38111,n38135,n38136,n38137);
  nand U40400(n38136,G60025,n36268);
  nand U40401(n38135,G60152,n36269);
  nand U40402(n38112,n38137,n34962);
  and U40403(n38137,n38138,n38139);
  nand U40404(n38139,G60184,n36266);
  nand U40405(n38138,G60057,n36267);
  nand U40406(n38045,n38140,n38141);
  nand U40407(n38141,n38142,n38143);
  not U40408(n38142,n38144);
  nand U40409(n38108,G60025,n36328);
  nand U40410(n38107,G60216,n34962);
  nand U40411(n38106,G60057,n37121);
  nand U40412(G14515,n38145,n38146,n38147,n38148);
  nor U40413(n38148,n38149,n38150,n38151);
  and U40414(n38151,n38152,n36729,G60023,n38082);
  nor U40415(n38150,n38153,n38152);
  nor U40416(n38153,n38154,n38155);
  nor U40417(n38154,G60023,n36226);
  nor U40418(n38149,n38156,n36233);
  nand U40419(n38147,n36234,n35512);
  nand U40420(n38146,n36235,n35295);
  xnor U40421(n35295,n38157,n38093);
  nand U40422(n38093,n38158,n38159,n38160,n38161);
  nor U40423(n38161,n38162,n38163);
  nor U40424(n38163,n38156,n36301);
  not U40425(n38156,G60215);
  nor U40426(n38162,n36302,n38152);
  not U40427(n38152,G60024);
  nand U40428(n38160,n36238,n35512);
  nand U40429(n38159,n38164,n36305);
  xor U40430(n38164,n35296,n38024);
  nand U40431(n38158,n35296,n36255);
  xnor U40432(n38157,n36238,n38094);
  nor U40433(n38094,n38165,n38166);
  nor U40434(n38165,n38167,n38168);
  nand U40435(n38145,n36272,n35296);
  nor U40436(n35296,n38027,n38169);
  and U40437(n38169,n38170,n38171);
  nor U40438(n38027,n38171,n38170);
  xor U40439(n38170,n38172,n36215);
  nand U40440(n38172,n38173,n38174,n38175,n38176);
  nand U40441(n38176,n35512,n36329);
  xor U40442(n35512,n38177,n38144);
  nand U40443(n38177,n38140,n38143);
  nand U40444(n38143,n38178,n38179,n38180);
  nand U40445(n38180,n35545,n38024);
  nand U40446(n38179,n38181,n34962);
  nand U40447(n38178,n38182,n35998);
  nand U40448(n38140,n38182,n38024,n35545);
  nand U40449(n38024,n38183,n38184,n38185,n38186);
  nor U40450(n38186,n38187,n38188,n38189,n38190);
  nor U40451(n38190,n36954,n37679);
  nand U40452(n37679,n38191,n38192);
  nor U40453(n38189,n36956,n37689);
  nand U40454(n37689,n38191,n38193);
  nor U40455(n38188,n36968,n37688);
  nand U40456(n37688,n38194,n38193);
  nor U40457(n38187,n36978,n37687);
  nand U40458(n37687,n38195,n38193);
  nor U40459(n38185,n38196,n38197,n38198,n38199);
  nor U40460(n38199,n36967,n37672);
  nand U40461(n37672,n38194,n38192);
  nor U40462(n38198,n36974,n37671);
  nand U40463(n37671,n38195,n38200);
  nor U40464(n38197,n36949,n37681);
  nand U40465(n37681,n38191,n38200);
  nor U40466(n38196,n36952,n37680);
  nand U40467(n37680,n38191,n38201);
  nor U40468(n38191,n38202,n38203);
  nor U40469(n38184,n38204,n38205,n38206,n38207);
  nor U40470(n38207,n36977,n37665);
  nand U40471(n37665,n38195,n38192);
  nor U40472(n38206,n36983,n37664);
  nand U40473(n37664,n38208,n38200);
  nor U40474(n38205,n36987,n37663);
  nand U40475(n37663,n38208,n38201);
  nor U40476(n38204,n36966,n37673);
  nand U40477(n37673,n38194,n38201);
  nor U40478(n38183,n38209,n38210,n38211,n38212);
  nor U40479(n38212,n36990,n37686);
  nand U40480(n37686,n38208,n38193);
  nor U40481(n38211,n36988,n37662);
  nand U40482(n37662,n38208,n38192);
  nor U40483(n38208,n38213,n38214);
  nor U40484(n38210,n36976,n37670);
  nand U40485(n37670,n38195,n38201);
  nor U40486(n38195,n38214,n38202);
  not U40487(n38202,n38213);
  nor U40488(n38209,n36964,n37678);
  nand U40489(n37678,n38194,n38200);
  nor U40490(n38194,n38213,n38203);
  not U40491(n38203,n38214);
  nand U40492(n38214,n38215,n38216,n38217);
  not U40493(n38217,n38218);
  nand U40494(n38216,G60007,n38219);
  nand U40495(n38215,n38220,G60009);
  xnor U40496(n38213,G60008,n38219);
  nand U40497(n38182,n38221,n38222,n38181);
  and U40498(n38181,n38223,n38224);
  nand U40499(n38224,G60183,n36266);
  nand U40500(n38223,G60056,n36267);
  nand U40501(n38222,G60024,n36268);
  nand U40502(n38221,G60151,n36269);
  nand U40503(n38175,G60024,n36328);
  nand U40504(n38174,G60215,n34962);
  nand U40505(n38173,G60056,n37121);
  or U40506(n38171,n38225,n38226);
  nand U40507(G14514,n38227,n38228,n38229,n38230);
  nor U40508(n38230,n38231,n38232,n38233);
  nor U40509(n38233,G60023,n38234,n36226);
  and U40510(n38232,n38155,G60023);
  nand U40511(n38155,n36288,n38235);
  nand U40512(n38235,n36729,n38234);
  not U40513(n38234,n38082);
  nor U40514(n38082,n38236,n38237);
  nor U40515(n38231,n38238,n36233);
  not U40516(n38238,G60214);
  nand U40517(n38229,n36234,n35516);
  nand U40518(n38228,n36235,n35305);
  xor U40519(n35305,n38167,n38239);
  nor U40520(n38239,n38168,n38166);
  nor U40521(n38166,n38240,n38241);
  and U40522(n38168,n38241,n38240);
  nand U40523(n38240,n38242,n38243,n38244,n38245);
  nand U40524(n38245,n38246,n35306);
  nand U40525(n38244,n35516,n36238);
  nand U40526(n38243,G60023,n36270);
  nand U40527(n38242,n36271,G60214);
  xnor U40528(n38241,n36246,n38247);
  nand U40529(n38247,n38248,n38249,n38250,n38251);
  nand U40530(n38251,n38252,n38253,n38254,n38255);
  nor U40531(n38255,n38256,n38257,n38258,n38259);
  nor U40532(n38259,n36388,n38260);
  nor U40533(n38258,n37020,n38261);
  nor U40534(n38257,n36376,n38262);
  nand U40535(n38256,n38263,n38264);
  nand U40536(n38264,n38265,G59894);
  nand U40537(n38263,n38266,G59886);
  nor U40538(n38254,n38267,n38268,n38269,n38270);
  nor U40539(n38270,n36386,n38271);
  nor U40540(n38269,n37014,n38272);
  nor U40541(n38268,n37008,n38273);
  nor U40542(n38267,n36370,n38274);
  nor U40543(n38253,n38275,n38276,n38277,n38278);
  nor U40544(n38278,n37018,n38279);
  nor U40545(n38277,n37016,n38280);
  nor U40546(n38276,n36382,n38281);
  nor U40547(n38275,n36384,n38282);
  nor U40548(n38252,n38283,n38284,n38285,n36246);
  nor U40549(n38285,n37004,n38286);
  nor U40550(n38284,n37006,n38287);
  nor U40551(n38283,n37002,n38288);
  nand U40552(n38250,n38289,n36922);
  nand U40553(n36922,n38290,n38291,n38292,n38293);
  nor U40554(n38293,n38294,n38295,n38296,n38297);
  nor U40555(n38297,n37006,n38298);
  nor U40556(n38296,n37004,n38299);
  nor U40557(n38295,n37002,n38300);
  nor U40558(n38294,n37018,n38301);
  nor U40559(n38292,n38302,n38303,n38304,n38305);
  nor U40560(n38305,n37016,n38306);
  nor U40561(n38304,n37014,n38307);
  nor U40562(n38303,n36386,n38308);
  nor U40563(n38302,n36384,n38309);
  nor U40564(n38291,n38310,n38311,n38312,n38313);
  nor U40565(n38313,n36382,n38314);
  nor U40566(n38312,n36374,n38315);
  nor U40567(n38311,n36372,n38316);
  nor U40568(n38310,n36370,n38317);
  nor U40569(n38290,n38318,n38319,n38320,n38321);
  nor U40570(n38321,n37008,n38322);
  nor U40571(n38320,n37020,n38323);
  nor U40572(n38319,n36388,n38324);
  nor U40573(n38318,n36376,n38325);
  nand U40574(n38249,n36305,n38326);
  nand U40575(n38326,n38327,n38328,n38329,n38330);
  nor U40576(n38330,n38331,n38332,n38333,n38334);
  nor U40577(n38334,n37008,n38335);
  nor U40578(n38333,n37006,n38336);
  nor U40579(n38332,n37004,n38337);
  nor U40580(n38331,n37002,n38338);
  nor U40581(n38329,n38339,n38340,n38341,n38342);
  nor U40582(n38342,n37020,n38343);
  nor U40583(n38341,n37018,n38344);
  nor U40584(n38340,n37016,n38345);
  nor U40585(n38339,n37014,n38346);
  nor U40586(n38328,n38347,n38348,n38349,n38350);
  nor U40587(n38350,n36388,n38351);
  nor U40588(n38349,n36386,n38352);
  nor U40589(n38348,n36384,n38353);
  nor U40590(n38347,n36382,n38354);
  nor U40591(n38327,n38355,n38356,n38357,n38358);
  nor U40592(n38358,n36376,n38359);
  nor U40593(n38357,n36374,n38360);
  nor U40594(n38356,n36372,n38361);
  nor U40595(n38355,n36370,n38362);
  nand U40596(n38248,n38363,n38364);
  nand U40597(n38167,n38365,n38366);
  nand U40598(n38227,n36272,n35306);
  nand U40599(n35306,n38367,n38368);
  nand U40600(n38368,n38369,n38370);
  or U40601(n38369,n38226,n38371);
  not U40602(n38226,n38372);
  nand U40603(n38367,n38225,n38372);
  nand U40604(n38372,n38373,n38374);
  nand U40605(n38374,n35545,G59998);
  nor U40606(n38225,n38370,n38371);
  nor U40607(n38371,n37008,n38373,n34968);
  nor U40608(n38373,n38375,n38376);
  and U40609(n38376,n38377,n36215);
  nor U40610(n38375,n38377,n35516,n36215);
  not U40611(n35516,n35304);
  nand U40612(n35304,n38144,n38378);
  nand U40613(n38378,n38379,n38380);
  xnor U40614(n38379,n35998,n38381);
  nand U40615(n38144,n38382,n38383);
  xnor U40616(n38382,n34962,n38381);
  and U40617(n38381,n38384,n38385,n38386,n38387);
  nand U40618(n38387,G60182,n36266);
  nand U40619(n38386,G60055,n36267);
  nand U40620(n38385,G60023,n36268);
  nand U40621(n38384,G60150,n36269);
  nand U40622(n38377,n38388,n38389,n38390);
  nand U40623(n38390,G60055,n37121);
  nand U40624(n38389,G60023,n36328);
  nand U40625(n38388,G60214,n34962);
  or U40626(n38370,n38391,n38392);
  and U40627(n38392,n38393,n38394);
  nand U40628(G14513,n38395,n38396,n38397,n38398);
  nor U40629(n38398,n38399,n38400,n38401);
  nor U40630(n38401,n35314,n36726);
  and U40631(n38400,n35317,n36272);
  nor U40632(n38399,n38402,n36233);
  not U40633(n38402,G60213);
  nand U40634(n38397,n36235,n35748);
  not U40635(n35748,n35316);
  nand U40636(n35316,n38403,n38404);
  nand U40637(n38404,n38405,n38406,n38407);
  nand U40638(n38405,n38408,n38365);
  nand U40639(n38403,n38409,n38365);
  nand U40640(n38365,n38410,n38411);
  xnor U40641(n38410,n38412,n36246);
  not U40642(n38409,n38366);
  nand U40643(n38366,n38408,n38413);
  nand U40644(n38413,n38407,n38406);
  nand U40645(n38407,n38414,n38415);
  nand U40646(n38408,n38416,n38417);
  xnor U40647(n38417,n36238,n38412);
  nand U40648(n38412,n38418,n38419,n38420,n38421);
  nand U40649(n38421,n38422,n38423,n38424,n38425);
  nor U40650(n38425,n38426,n38427,n38428,n38429);
  nor U40651(n38429,n36458,n38260);
  nor U40652(n38428,n36469,n38261);
  nor U40653(n38427,n36450,n38262);
  nand U40654(n38426,n38430,n38431);
  nand U40655(n38431,n38265,G59895);
  nand U40656(n38430,n38266,G59887);
  nor U40657(n38424,n38432,n38433,n38434,n38435);
  nor U40658(n38435,n36457,n38271);
  nor U40659(n38434,n36463,n38272);
  nor U40660(n38433,n36481,n38273);
  nor U40661(n38432,n36447,n38274);
  nor U40662(n38423,n38436,n38437,n38438,n38439);
  nor U40663(n38439,n36467,n38279);
  nor U40664(n38438,n36465,n38280);
  nor U40665(n38437,n36455,n38281);
  nor U40666(n38436,n36456,n38282);
  nor U40667(n38422,n38440,n38441,n38442,n36246);
  nor U40668(n38442,n36477,n38286);
  nor U40669(n38441,n36479,n38287);
  nor U40670(n38440,n36475,n38288);
  nand U40671(n38420,n38289,n37076);
  nand U40672(n37076,n38443,n38444,n38445,n38446);
  nor U40673(n38446,n38447,n38448,n38449,n38450);
  nor U40674(n38450,n36479,n38298);
  nor U40675(n38449,n36477,n38299);
  nor U40676(n38448,n36475,n38300);
  nor U40677(n38447,n36467,n38301);
  nor U40678(n38445,n38451,n38452,n38453,n38454);
  nor U40679(n38454,n36465,n38306);
  nor U40680(n38453,n36463,n38307);
  nor U40681(n38452,n36457,n38308);
  nor U40682(n38451,n36456,n38309);
  nor U40683(n38444,n38455,n38456,n38457,n38458);
  nor U40684(n38458,n36455,n38314);
  nor U40685(n38457,n36449,n38315);
  nor U40686(n38456,n36448,n38316);
  nor U40687(n38455,n36447,n38317);
  nor U40688(n38443,n38459,n38460,n38461,n38462);
  nor U40689(n38462,n36481,n38322);
  nor U40690(n38461,n36469,n38323);
  nor U40691(n38460,n36458,n38324);
  nor U40692(n38459,n36450,n38325);
  nand U40693(n38419,n38363,n38463);
  nand U40694(n38463,n38464,n38465,n38466,n38467);
  nor U40695(n38467,n38468,n38469,n38470,n38471);
  nor U40696(n38471,n36477,n38472);
  nor U40697(n38470,n36475,n38473);
  nor U40698(n38469,n36469,n38474);
  nor U40699(n38468,n36465,n38475);
  nor U40700(n38466,n38476,n38477,n38478,n38479);
  nor U40701(n38479,n36463,n38480);
  nor U40702(n38478,n36458,n38481);
  nor U40703(n38477,n36456,n38482);
  nor U40704(n38476,n36455,n38483);
  nor U40705(n38465,n38484,n38485,n38486,n38487);
  nor U40706(n38487,n36450,n38488);
  nor U40707(n38486,n36448,n38489);
  nor U40708(n38485,n36447,n38490);
  nor U40709(n38484,n36481,n38491);
  nor U40710(n38464,n38492,n38493,n38494,n38495);
  nor U40711(n38495,n36479,n38496);
  nor U40712(n38494,n36467,n38497);
  nor U40713(n38493,n36457,n38498);
  nor U40714(n38492,n36449,n38499);
  nand U40715(n38418,n36305,n38500);
  nand U40716(n38500,n38501,n38502,n38503,n38504);
  nor U40717(n38504,n38505,n38506,n38507,n38508);
  nor U40718(n38508,n36481,n38335);
  nor U40719(n38507,n36479,n38336);
  nor U40720(n38506,n36477,n38337);
  nor U40721(n38505,n36475,n38338);
  nor U40722(n38503,n38509,n38510,n38511,n38512);
  nor U40723(n38512,n36469,n38343);
  nor U40724(n38511,n36467,n38344);
  nor U40725(n38510,n36465,n38345);
  nor U40726(n38509,n36463,n38346);
  nor U40727(n38502,n38513,n38514,n38515,n38516);
  nor U40728(n38516,n36458,n38351);
  nor U40729(n38515,n36457,n38352);
  nor U40730(n38514,n36456,n38353);
  nor U40731(n38513,n36455,n38354);
  nor U40732(n38501,n38517,n38518,n38519,n38520);
  nor U40733(n38520,n36450,n38359);
  nor U40734(n38519,n36449,n38360);
  nor U40735(n38518,n36448,n38361);
  nor U40736(n38517,n36447,n38362);
  not U40737(n38416,n38411);
  nand U40738(n38411,n38521,n38522,n38523,n38524);
  nand U40739(n38524,n35317,n38246);
  xor U40740(n35317,n38394,n38525);
  nor U40741(n38525,n38391,n38526);
  not U40742(n38526,n38393);
  nand U40743(n38393,n38527,n38528);
  nand U40744(n38528,n35545,G59999);
  nor U40745(n38391,n34968,n36481,n38527);
  xor U40746(n38527,n38529,n36215);
  nand U40747(n38529,n38530,n38531,n38532,n38533);
  nand U40748(n38533,n35520,n36329);
  nand U40749(n38532,G60022,n36328);
  nand U40750(n38531,G60213,n34962);
  nand U40751(n38530,G60054,n37121);
  nand U40752(n38394,n38534,n38535);
  nand U40753(n38535,n38536,n38537);
  nand U40754(n38536,n38538,n38539);
  nand U40755(n38539,n35545,G60000);
  not U40756(n38534,n38540);
  nand U40757(n38523,n36238,n35520);
  not U40758(n35520,n35314);
  nand U40759(n35314,n38380,n38541);
  nand U40760(n38541,n38542,n38543);
  not U40761(n38380,n38383);
  nor U40762(n38383,n38543,n38542);
  xor U40763(n38542,n34962,n38544);
  nor U40764(n38544,n38545,n38546,n38547,n38548);
  and U40765(n38548,n36269,G60149);
  and U40766(n38547,n36268,G60022);
  nor U40767(n38546,n36215,n36172);
  not U40768(n36172,G60054);
  nor U40769(n38545,n38073,n35315);
  not U40770(n35315,G60181);
  nand U40771(n38522,G60022,n36270);
  nand U40772(n38521,n36271,G60213);
  nand U40773(n38396,n38549,n38237,n36729);
  nand U40774(n38237,G60022,n34912);
  nand U40775(n38395,G60022,n38550);
  nand U40776(n38550,n36288,n38551);
  nand U40777(n38551,n36729,n38236);
  not U40778(n38236,n38549);
  nor U40779(n38549,n38552,n38553,n38554);
  nand U40780(G14512,n38555,n38556,n38557,n38558);
  nor U40781(n38558,n38559,n38560,n38561);
  nor U40782(n38561,G60021,n36226,n38553,n38554);
  nor U40783(n38560,n38562,n38552);
  nor U40784(n38562,n38563,n36231);
  nor U40785(n38563,n38564,n36226);
  nor U40786(n38564,n38553,n38554);
  nor U40787(n38559,n38565,n36233);
  not U40788(n38565,G60212);
  nand U40789(n38557,n36234,n35524);
  nand U40790(n38556,n36235,n35328);
  xor U40791(n35328,n38415,n38566);
  and U40792(n38566,n38414,n38406);
  nand U40793(n38406,n38567,n38568);
  or U40794(n38414,n38568,n38567);
  xnor U40795(n38567,n38569,n36246);
  nand U40796(n38569,n38570,n38571,n38572,n38573);
  nand U40797(n38573,n38574,n38575,n38576,n38577);
  nor U40798(n38577,n38578,n38579,n38580,n38581);
  nor U40799(n38581,n36562,n38260);
  nor U40800(n38580,n37188,n38261);
  nor U40801(n38579,n36554,n38262);
  nand U40802(n38578,n38582,n38583);
  nand U40803(n38583,n38265,G59896);
  nand U40804(n38582,n38266,G59888);
  nor U40805(n38576,n38584,n38585,n38586,n38587);
  nor U40806(n38587,n36561,n38271);
  nor U40807(n38586,n37185,n38272);
  nor U40808(n38585,n37180,n38273);
  nor U40809(n38584,n36551,n38274);
  nor U40810(n38575,n38588,n38589,n38590,n38591);
  nor U40811(n38591,n37187,n38279);
  nor U40812(n38590,n37186,n38280);
  nor U40813(n38589,n36559,n38281);
  nor U40814(n38588,n36560,n38282);
  nor U40815(n38574,n38592,n38593,n38594,n36246);
  nor U40816(n38594,n37178,n38286);
  nor U40817(n38593,n37179,n38287);
  nor U40818(n38592,n37177,n38288);
  nand U40819(n38572,n38289,n37155);
  nand U40820(n37155,n38595,n38596,n38597,n38598);
  nor U40821(n38598,n38599,n38600,n38601,n38602);
  nor U40822(n38602,n37179,n38298);
  nor U40823(n38601,n37178,n38299);
  nor U40824(n38600,n37177,n38300);
  nor U40825(n38599,n37187,n38301);
  nor U40826(n38597,n38603,n38604,n38605,n38606);
  nor U40827(n38606,n37186,n38306);
  nor U40828(n38605,n37185,n38307);
  nor U40829(n38604,n36561,n38308);
  nor U40830(n38603,n36560,n38309);
  nor U40831(n38596,n38607,n38608,n38609,n38610);
  nor U40832(n38610,n36559,n38314);
  nor U40833(n38609,n36553,n38315);
  nor U40834(n38608,n36552,n38316);
  nor U40835(n38607,n36551,n38317);
  nor U40836(n38595,n38611,n38612,n38613,n38614);
  nor U40837(n38614,n37180,n38322);
  nor U40838(n38613,n37188,n38323);
  nor U40839(n38612,n36562,n38324);
  nor U40840(n38611,n36554,n38325);
  nand U40841(n38571,n38363,n38615);
  nand U40842(n38615,n38616,n38617,n38618,n38619);
  nor U40843(n38619,n38620,n38621,n38622,n38623);
  nor U40844(n38623,n37178,n38472);
  nor U40845(n38622,n37177,n38473);
  nor U40846(n38621,n37188,n38474);
  nor U40847(n38620,n37186,n38475);
  nor U40848(n38618,n38624,n38625,n38626,n38627);
  nor U40849(n38627,n37185,n38480);
  nor U40850(n38626,n36562,n38481);
  nor U40851(n38625,n36560,n38482);
  nor U40852(n38624,n36559,n38483);
  nor U40853(n38617,n38628,n38629,n38630,n38631);
  nor U40854(n38631,n36554,n38488);
  nor U40855(n38630,n36552,n38489);
  nor U40856(n38629,n36551,n38490);
  nor U40857(n38628,n37180,n38491);
  nor U40858(n38616,n38632,n38633,n38634,n38635);
  nor U40859(n38635,n37179,n38496);
  nor U40860(n38634,n37187,n38497);
  nor U40861(n38633,n36561,n38498);
  nor U40862(n38632,n36553,n38499);
  nand U40863(n38570,n36305,n38636);
  nand U40864(n38636,n38637,n38638,n38639,n38640);
  nor U40865(n38640,n38641,n38642,n38643,n38644);
  nor U40866(n38644,n37180,n38335);
  nor U40867(n38643,n37179,n38336);
  nor U40868(n38642,n37178,n38337);
  nor U40869(n38641,n37177,n38338);
  nor U40870(n38639,n38645,n38646,n38647,n38648);
  nor U40871(n38648,n37188,n38343);
  nor U40872(n38647,n37187,n38344);
  nor U40873(n38646,n37186,n38345);
  nor U40874(n38645,n37185,n38346);
  nor U40875(n38638,n38649,n38650,n38651,n38652);
  nor U40876(n38652,n36562,n38351);
  nor U40877(n38651,n36561,n38352);
  nor U40878(n38650,n36560,n38353);
  nor U40879(n38649,n36559,n38354);
  nor U40880(n38637,n38653,n38654,n38655,n38656);
  nor U40881(n38656,n36554,n38359);
  nor U40882(n38655,n36553,n38360);
  nor U40883(n38654,n36552,n38361);
  nor U40884(n38653,n36551,n38362);
  nand U40885(n38568,n38657,n38658,n38659,n38660);
  nand U40886(n38660,n35329,n38246);
  nand U40887(n38659,n35524,n36238);
  nand U40888(n38658,G60021,n36270);
  nand U40889(n38657,n36271,G60212);
  nand U40890(n38415,n38661,n38662);
  nand U40891(n38662,n38663,n38664);
  nand U40892(n38663,n38665,n38666);
  or U40893(n38661,n38666,n38665);
  xor U40894(n35329,n38537,n38667);
  nor U40895(n38667,n38668,n38540);
  nor U40896(n38540,n37180,n38538,n34968);
  nor U40897(n38668,n38669,n38670);
  not U40898(n38670,n38538);
  nor U40899(n38538,n38671,n38672);
  and U40900(n38672,n38673,n36215);
  nor U40901(n38671,n38673,n35524,n36215);
  not U40902(n35524,n35325);
  nand U40903(n35325,n38543,n38674);
  nand U40904(n38674,n38675,n38676);
  or U40905(n38543,n38676,n38675);
  xor U40906(n38675,n34962,n38677);
  nor U40907(n38677,n38678,n38679,n38680,n38681);
  and U40908(n38681,n36269,G60148);
  nor U40909(n38680,n36527,n38552);
  not U40910(n38552,G60021);
  nor U40911(n38679,n36215,n36179);
  not U40912(n36179,G60053);
  nor U40913(n38678,n38073,n35326);
  not U40914(n35326,G60180);
  nand U40915(n38676,n38682,n38683);
  nand U40916(n38673,n38684,n38685,n38686);
  nand U40917(n38686,G60053,n37121);
  nand U40918(n38685,G60021,n36328);
  nand U40919(n38684,G60212,n34962);
  nor U40920(n38669,n37180,n34968);
  nand U40921(n38537,n38687,n38688);
  nand U40922(n38688,n38689,n38690);
  nand U40923(G14511,n38691,n38692,n38693,n38694);
  nor U40924(n38694,n38695,n38696,n38697);
  nor U40925(n38697,G60020,n38554,n36226);
  not U40926(n38554,n38698);
  nor U40927(n38696,n38699,n38553);
  nor U40928(n38699,n38700,n36231);
  nor U40929(n38700,n38698,n36226);
  nor U40930(n38698,n38701,n38702);
  nor U40931(n38695,n38703,n36233);
  nand U40932(n38692,n36235,n35340);
  xor U40933(n35340,n38704,n38666);
  xor U40934(n38666,n38705,n36246);
  nand U40935(n38705,n38706,n38707,n38708,n38709);
  nor U40936(n38709,n38710,n38711);
  nor U40937(n38711,n38712,n38713);
  and U40938(n38710,n37231,n38289);
  nand U40939(n37231,n38714,n38715,n38716,n38717);
  nor U40940(n38717,n38718,n38719,n38720,n38721);
  nor U40941(n38721,n37261,n38298);
  nor U40942(n38720,n37260,n38299);
  nor U40943(n38719,n37259,n38300);
  nor U40944(n38718,n37269,n38301);
  nor U40945(n38716,n38722,n38723,n38724,n38725);
  nor U40946(n38725,n37268,n38306);
  nor U40947(n38724,n37267,n38307);
  nor U40948(n38723,n36640,n38308);
  nor U40949(n38722,n36639,n38309);
  nor U40950(n38715,n38726,n38727,n38728,n38729);
  nor U40951(n38729,n36638,n38314);
  nor U40952(n38728,n36632,n38315);
  nor U40953(n38727,n36631,n38316);
  nor U40954(n38726,n36630,n38317);
  nor U40955(n38714,n38730,n38731,n38732,n38733);
  nor U40956(n38733,n37262,n38322);
  nor U40957(n38732,n37270,n38323);
  nor U40958(n38731,n36641,n38324);
  nor U40959(n38730,n36633,n38325);
  nand U40960(n38708,n36305,n38734);
  nand U40961(n38734,n38735,n38736,n38737,n38738);
  nor U40962(n38738,n38739,n38740,n38741,n38742);
  nor U40963(n38742,n37262,n38335);
  nor U40964(n38741,n37261,n38336);
  nor U40965(n38740,n37260,n38337);
  nor U40966(n38739,n37259,n38338);
  nor U40967(n38737,n38743,n38744,n38745,n38746);
  nor U40968(n38746,n37270,n38343);
  nor U40969(n38745,n37269,n38344);
  nor U40970(n38744,n37268,n38345);
  nor U40971(n38743,n37267,n38346);
  nor U40972(n38736,n38747,n38748,n38749,n38750);
  nor U40973(n38750,n36641,n38351);
  nor U40974(n38749,n36640,n38352);
  nor U40975(n38748,n36639,n38353);
  nor U40976(n38747,n36638,n38354);
  nor U40977(n38735,n38751,n38752,n38753,n38754);
  nor U40978(n38754,n36633,n38359);
  nor U40979(n38753,n36632,n38360);
  nor U40980(n38752,n36631,n38361);
  nor U40981(n38751,n36630,n38362);
  nand U40982(n38707,n38755,n38756,n38757,n38758);
  nor U40983(n38758,n38759,n38760,n38761,n38762);
  nor U40984(n38762,n36641,n38260);
  nor U40985(n38761,n37270,n38261);
  nor U40986(n38760,n36633,n38262);
  nand U40987(n38759,n38763,n38764);
  nand U40988(n38764,n38265,G59897);
  nand U40989(n38763,n38266,G59889);
  nor U40990(n38757,n38765,n38766,n38767,n38768);
  nor U40991(n38768,n36640,n38271);
  nor U40992(n38767,n37267,n38272);
  nor U40993(n38766,n37262,n38273);
  nor U40994(n38765,n36630,n38274);
  nor U40995(n38756,n38769,n38770,n38771,n38772);
  nor U40996(n38772,n37269,n38279);
  nor U40997(n38771,n37268,n38280);
  nor U40998(n38770,n36638,n38281);
  nor U40999(n38769,n36639,n38282);
  nor U41000(n38755,n38773,n38774,n38775,n36246);
  nor U41001(n38775,n37260,n38286);
  nor U41002(n38774,n37261,n38287);
  nor U41003(n38773,n37259,n38288);
  nand U41004(n38706,n38363,n38776);
  nand U41005(n38776,n38777,n38778,n38779,n38780);
  nor U41006(n38780,n38781,n38782,n38783,n38784);
  nor U41007(n38784,n37260,n38472);
  nor U41008(n38783,n37259,n38473);
  nor U41009(n38782,n37270,n38474);
  nor U41010(n38781,n37268,n38475);
  nor U41011(n38779,n38785,n38786,n38787,n38788);
  nor U41012(n38788,n37267,n38480);
  nor U41013(n38787,n36641,n38481);
  nor U41014(n38786,n36639,n38482);
  nor U41015(n38785,n36638,n38483);
  nor U41016(n38778,n38789,n38790,n38791,n38792);
  nor U41017(n38792,n36633,n38488);
  nor U41018(n38791,n36631,n38489);
  nor U41019(n38790,n36630,n38490);
  nor U41020(n38789,n37262,n38491);
  nor U41021(n38777,n38793,n38794,n38795,n38796);
  nor U41022(n38796,n37261,n38496);
  nor U41023(n38795,n37269,n38497);
  nor U41024(n38794,n36640,n38498);
  nor U41025(n38793,n36632,n38499);
  xor U41026(n38704,n38664,n38665);
  and U41027(n38665,n38797,n38798,n38799,n38800);
  nand U41028(n38800,n34840,n38246);
  nand U41029(n38799,G60020,n36270);
  nand U41030(n38798,n36238,n35528);
  nand U41031(n38797,n36271,G60211);
  nand U41032(n38664,n38801,n38802);
  nand U41033(n38802,n38803,n38804);
  nand U41034(n38691,n36234,n35528);
  nand U41035(G14510,n38805,n38806,n38807,n38808);
  nor U41036(n38808,n38809,n38810,n38811);
  nor U41037(n38811,G60019,n38701,n36226);
  nor U41038(n38810,n38812,n38702);
  nor U41039(n38812,n38813,n36231);
  and U41040(n38813,n38701,n36729);
  nand U41041(n38701,n34912,n38814);
  nand U41042(n38814,n38815,n38816);
  nor U41043(n38809,n35351,n36233);
  nand U41044(n38806,n36235,n35353);
  xor U41045(n35353,n38804,n38817);
  and U41046(n38817,n38801,n38803);
  or U41047(n38803,n38818,n38819);
  nand U41048(n38801,n38819,n38818);
  nand U41049(n38818,n38820,n38821,n38822,n38823);
  nand U41050(n38823,n34850,n38246);
  nand U41051(n38822,G60019,n36270);
  nand U41052(n38821,n36238,n35352);
  nand U41053(n38820,n36271,G60210);
  xnor U41054(n38819,n36246,n38824);
  nand U41055(n38824,n38825,n38826,n38827,n38828);
  nor U41056(n38828,n38829,n38830);
  nor U41057(n38830,n38712,n38831);
  nor U41058(n38829,n38832,n35781);
  nor U41059(n38832,n38833,n38834,n38835,n38836);
  nand U41060(n38836,n38837,n38838,n38839,n38840);
  nand U41061(n38840,n38841,G59882);
  nand U41062(n38839,n38842,G59890);
  nand U41063(n38838,n38843,G59898);
  nand U41064(n38837,n38844,G59906);
  nand U41065(n38835,n38845,n38846,n38847,n38848);
  nand U41066(n38848,n38849,G59914);
  nand U41067(n38847,n38850,G59922);
  nand U41068(n38846,n38851,G59930);
  nand U41069(n38845,n38852,G59938);
  nand U41070(n38834,n38853,n38854,n38855,n38856);
  nand U41071(n38856,n38857,G59946);
  nand U41072(n38855,n38858,G59954);
  nand U41073(n38854,n38859,G59962);
  nand U41074(n38853,n38860,G59970);
  nand U41075(n38833,n38861,n38862,n38863,n38864);
  nand U41076(n38864,n38865,G59978);
  nand U41077(n38863,n38866,G59986);
  nand U41078(n38862,n38867,G59994);
  nand U41079(n38861,n38868,G60002);
  nand U41080(n38827,n38289,n37315);
  nand U41081(n37315,n38869,n38870,n38871,n38872);
  nor U41082(n38872,n38873,n38874,n38875,n38876);
  nor U41083(n38876,n37344,n38298);
  nor U41084(n38875,n37343,n38299);
  nor U41085(n38874,n37342,n38300);
  nor U41086(n38873,n37352,n38301);
  nor U41087(n38871,n38877,n38878,n38879,n38880);
  nor U41088(n38880,n37351,n38306);
  nor U41089(n38879,n37350,n38307);
  nor U41090(n38878,n36716,n38308);
  nor U41091(n38877,n36715,n38309);
  nor U41092(n38870,n38881,n38882,n38883,n38884);
  nor U41093(n38884,n36714,n38314);
  nor U41094(n38883,n36708,n38315);
  nor U41095(n38882,n36707,n38316);
  nor U41096(n38881,n36706,n38317);
  nor U41097(n38869,n38885,n38886,n38887,n38888);
  nor U41098(n38888,n37345,n38322);
  nor U41099(n38887,n37353,n38323);
  nor U41100(n38886,n36717,n38324);
  nor U41101(n38885,n36709,n38325);
  nand U41102(n38826,n38889,n38890,n38891,n38892);
  nor U41103(n38892,n38893,n38894,n38895,n38896);
  nor U41104(n38896,n36717,n38260);
  nor U41105(n38895,n37353,n38261);
  nor U41106(n38894,n36709,n38262);
  nand U41107(n38893,n38897,n38898);
  nand U41108(n38898,n38265,G59898);
  nand U41109(n38897,n38266,G59890);
  nor U41110(n38891,n38899,n38900,n38901,n38902);
  nor U41111(n38902,n36716,n38271);
  nor U41112(n38901,n37350,n38272);
  nor U41113(n38900,n37345,n38273);
  nor U41114(n38899,n36706,n38274);
  nor U41115(n38890,n38903,n38904,n38905,n38906);
  nor U41116(n38906,n37352,n38279);
  nor U41117(n38905,n37351,n38280);
  nor U41118(n38904,n36714,n38281);
  nor U41119(n38903,n36715,n38282);
  nor U41120(n38889,n38907,n38908,n38909,n36246);
  nor U41121(n38909,n37343,n38286);
  nor U41122(n38908,n37344,n38287);
  nor U41123(n38907,n37342,n38288);
  nand U41124(n38825,n38363,n38910);
  nand U41125(n38910,n38911,n38912,n38913,n38914);
  nor U41126(n38914,n38915,n38916,n38917,n38918);
  nor U41127(n38918,n37343,n38472);
  nor U41128(n38917,n37342,n38473);
  nor U41129(n38916,n37353,n38474);
  nor U41130(n38915,n37351,n38475);
  nor U41131(n38913,n38919,n38920,n38921,n38922);
  nor U41132(n38922,n37350,n38480);
  nor U41133(n38921,n36717,n38481);
  nor U41134(n38920,n36715,n38482);
  nor U41135(n38919,n36714,n38483);
  nor U41136(n38912,n38923,n38924,n38925,n38926);
  nor U41137(n38926,n36709,n38488);
  nor U41138(n38925,n36707,n38489);
  nor U41139(n38924,n36706,n38490);
  nor U41140(n38923,n37345,n38491);
  nor U41141(n38911,n38927,n38928,n38929,n38930);
  nor U41142(n38930,n37344,n38496);
  nor U41143(n38929,n37352,n38497);
  nor U41144(n38928,n36716,n38498);
  nor U41145(n38927,n36708,n38499);
  nand U41146(n38804,n38931,n38932);
  nand U41147(n38932,n38933,n38934);
  nand U41148(n38805,n36234,n35352);
  nand U41149(G14509,n38935,n38936,n38937,n38938);
  nor U41150(n38938,n38939,n38940,n38941);
  and U41151(n38941,n38815,n38816,n36729);
  not U41152(n36729,n36226);
  nor U41153(n38940,n38942,n38815);
  nor U41154(n38942,n38943,n36231);
  nor U41155(n38943,n36226,n38816);
  nand U41156(n38816,G60016,n34912,G60017);
  nor U41157(n38939,n35363,n36233);
  not U41158(n35363,G60209);
  nand U41159(n38936,n36235,n35365);
  xor U41160(n35365,n38933,n38944);
  and U41161(n38944,n38934,n38931);
  nand U41162(n38931,n38945,n38946);
  nand U41163(n38946,n38947,n38948);
  nand U41164(n38934,n38947,n38948,n38949);
  not U41165(n38949,n38945);
  nand U41166(n38945,n38950,n38951,n38952,n38953);
  nand U41167(n38953,n34860,n38246);
  nand U41168(n38246,n36582,n35781);
  nand U41169(n38952,G60018,n36270);
  not U41170(n36270,n36302);
  nand U41171(n38951,n36238,n35364);
  nand U41172(n38950,n36271,G60209);
  not U41173(n36271,n36301);
  nand U41174(n38948,n36238,n38954,n38955);
  nand U41175(n38954,n38956,n38957,n38958,n38959);
  nor U41176(n38959,n38960,n38961,n38962,n38963);
  nor U41177(n38963,n36777,n38964);
  nor U41178(n38962,n36778,n38262);
  nor U41179(n38961,n36786,n38260);
  nor U41180(n38960,n36794,n38261);
  nor U41181(n38958,n38965,n38966,n38967,n38968);
  nor U41182(n38968,n36791,n38272);
  nor U41183(n38967,n36802,n38273);
  nor U41184(n38966,n36775,n38274);
  nor U41185(n38965,n36776,n38969);
  nor U41186(n38957,n38970,n38971,n38972,n38973);
  nor U41187(n38973,n36792,n38280);
  nor U41188(n38972,n36783,n38281);
  nor U41189(n38971,n36784,n38282);
  nor U41190(n38970,n36785,n38271);
  nor U41191(n38956,n38974,n38975,n38976,n38977);
  nor U41192(n38977,n36800,n38286);
  nor U41193(n38976,n36801,n38287);
  nor U41194(n38975,n36799,n38288);
  nor U41195(n38974,n36793,n38279);
  nand U41196(n38947,n38978,n36246);
  nand U41197(n38978,n38955,n38979,n38980,n38981);
  nand U41198(n38980,n38363,n38982);
  nand U41199(n38982,n38983,n38984,n38985,n38986);
  nor U41200(n38986,n38987,n38988,n38989,n38990);
  nor U41201(n38990,n36800,n38472);
  nor U41202(n38989,n36799,n38473);
  nor U41203(n38988,n36794,n38474);
  nor U41204(n38987,n36792,n38475);
  nor U41205(n38985,n38991,n38992,n38993,n38994);
  nor U41206(n38994,n36791,n38480);
  nor U41207(n38993,n36786,n38481);
  nor U41208(n38992,n36784,n38482);
  nor U41209(n38991,n36783,n38483);
  nor U41210(n38984,n38995,n38996,n38997,n38998);
  nor U41211(n38998,n36778,n38488);
  nor U41212(n38997,n36776,n38489);
  nor U41213(n38996,n36775,n38490);
  nor U41214(n38995,n36802,n38491);
  nor U41215(n38983,n38999,n39000,n39001,n39002);
  nor U41216(n39002,n36801,n38496);
  nor U41217(n39001,n36793,n38497);
  nor U41218(n39000,n36785,n38498);
  nor U41219(n38999,n36777,n38499);
  nand U41220(n38979,n38289,n37400);
  nand U41221(n37400,n39003,n39004,n39005,n39006);
  nor U41222(n39006,n39007,n39008,n39009,n39010);
  nor U41223(n39010,n36801,n38298);
  nor U41224(n39009,n36800,n38299);
  nor U41225(n39008,n36799,n38300);
  nor U41226(n39007,n36793,n38301);
  nor U41227(n39005,n39011,n39012,n39013,n39014);
  nor U41228(n39014,n36792,n38306);
  nor U41229(n39013,n36791,n38307);
  nor U41230(n39012,n36785,n38308);
  nor U41231(n39011,n36784,n38309);
  nor U41232(n39004,n39015,n39016,n39017,n39018);
  nor U41233(n39018,n36783,n38314);
  nor U41234(n39017,n36777,n38315);
  nor U41235(n39016,n36776,n38316);
  nor U41236(n39015,n36775,n38317);
  nor U41237(n39003,n39019,n39020,n39021,n39022);
  nor U41238(n39022,n36802,n38322);
  nor U41239(n39021,n36794,n38323);
  nor U41240(n39020,n36786,n38324);
  nor U41241(n39019,n36778,n38325);
  and U41242(n38955,n39023,n39024);
  nand U41243(n39024,n36305,n39025);
  nand U41244(n39025,n39026,n39027,n39028,n39029);
  nor U41245(n39029,n39030,n39031,n39032,n39033);
  nor U41246(n39033,n36802,n38335);
  nor U41247(n39032,n36801,n38336);
  nor U41248(n39031,n36800,n38337);
  nor U41249(n39030,n36799,n38338);
  nor U41250(n39028,n39034,n39035,n39036,n39037);
  nor U41251(n39037,n36794,n38343);
  nor U41252(n39036,n36793,n38344);
  nor U41253(n39035,n36792,n38345);
  nor U41254(n39034,n36791,n38346);
  nor U41255(n39027,n39038,n39039,n39040,n39041);
  nor U41256(n39041,n36786,n38351);
  nor U41257(n39040,n36785,n38352);
  nor U41258(n39039,n36784,n38353);
  nor U41259(n39038,n36783,n38354);
  nor U41260(n39026,n39042,n39043,n39044,n39045);
  nor U41261(n39045,n36778,n38359);
  nor U41262(n39044,n36777,n38360);
  nor U41263(n39043,n36776,n38361);
  nor U41264(n39042,n36775,n38362);
  nand U41265(n39023,G60008,n35695);
  nand U41266(n38933,n39046,n39047);
  nand U41267(n39047,n39048,n39049);
  nand U41268(n38935,n36234,n35364);
  nand U41269(G14508,n39050,n39051,n39052,n39053);
  nor U41270(n39053,n39054,n39055,n39056);
  nor U41271(n39056,G60017,n39057,n36226);
  nor U41272(n39055,n39058,n39059);
  nor U41273(n39058,n39060,n36231);
  nor U41274(n39054,n34984,n36233);
  nand U41275(n39051,n36235,n35376);
  xor U41276(n35376,n39049,n39061);
  and U41277(n39061,n39048,n39046);
  or U41278(n39046,n39062,n39063);
  nand U41279(n39048,n39063,n39062);
  xor U41280(n39062,n39064,n36246);
  nand U41281(n39064,n39065,n39066,n39067,n39068);
  nor U41282(n39068,n39069,n39070,n39071,n39072);
  nor U41283(n39072,n39073,n35781);
  nor U41284(n39073,n39074,n39075,n39076,n39077);
  nand U41285(n39077,n39078,n39079,n39080,n39081);
  nand U41286(n39081,n38841,G59884);
  nand U41287(n39080,n38842,G59892);
  nand U41288(n39079,n38843,G59900);
  nand U41289(n39078,n38844,G59908);
  nand U41290(n39076,n39082,n39083,n39084,n39085);
  nand U41291(n39085,n38849,G59916);
  nand U41292(n39084,n38850,G59924);
  nand U41293(n39083,n38851,G59932);
  nand U41294(n39082,n38852,G59940);
  nand U41295(n39075,n39086,n39087,n39088,n39089);
  nand U41296(n39089,n38857,G59948);
  nand U41297(n39088,n38858,G59956);
  nand U41298(n39087,n38859,G59964);
  nand U41299(n39086,n38860,G59972);
  nand U41300(n39074,n39090,n39091,n39092,n39093);
  nand U41301(n39093,n38865,G59980);
  nand U41302(n39092,n38866,G59988);
  nand U41303(n39091,n38867,G59996);
  nand U41304(n39090,n38868,G60004);
  nor U41305(n39071,n39094,n39095,n39096,n39097);
  nand U41306(n39097,n36238,n39098,n39099,n39100);
  nand U41307(n39100,n39101,G59972);
  nand U41308(n39099,n39102,G59940);
  nand U41309(n39098,n39103,G59908);
  nand U41310(n39096,n39104,n39105,n39106,n39107);
  nand U41311(n39107,n38265,G59900);
  nand U41312(n39106,n38266,G59892);
  nand U41313(n39105,n39108,G59884);
  nand U41314(n39104,n39109,G60004);
  nand U41315(n39095,n39110,n39111,n39112,n39113);
  nand U41316(n39113,n39114,G59948);
  nand U41317(n39112,n39115,G59932);
  nand U41318(n39111,n39116,G59924);
  nand U41319(n39110,n39117,G59916);
  nand U41320(n39094,n39118,n39119,n39120,n39121);
  nor U41321(n39121,n39122,n39123);
  nor U41322(n39123,n36896,n38286);
  nor U41323(n39122,n36897,n38287);
  nand U41324(n39120,n39124,G59980);
  nand U41325(n39119,n39125,G59956);
  nand U41326(n39118,n39126,G59964);
  nand U41327(n39067,G60009,n35695);
  nand U41328(n39066,n38363,n39127);
  nand U41329(n39127,n39128,n39129,n39130,n39131);
  nor U41330(n39131,n39132,n39133,n39134,n39135);
  nor U41331(n39135,n36896,n38472);
  nor U41332(n39134,n36895,n38473);
  nor U41333(n39133,n36890,n38474);
  nor U41334(n39132,n36888,n38475);
  nor U41335(n39130,n39136,n39137,n39138,n39139);
  nor U41336(n39139,n36887,n38480);
  nor U41337(n39138,n36882,n38481);
  nor U41338(n39137,n36880,n38482);
  nor U41339(n39136,n36879,n38483);
  nor U41340(n39129,n39140,n39141,n39142,n39143);
  nor U41341(n39143,n36874,n38488);
  nor U41342(n39142,n36872,n38489);
  nor U41343(n39141,n36871,n38490);
  nor U41344(n39140,n36898,n38491);
  nor U41345(n39128,n39144,n39145,n39146,n39147);
  nor U41346(n39147,n36897,n38496);
  nor U41347(n39146,n36889,n38497);
  nor U41348(n39145,n36881,n38498);
  nor U41349(n39144,n36873,n38499);
  nand U41350(n39065,n38289,n37474);
  nand U41351(n37474,n39148,n39149,n39150,n39151);
  nor U41352(n39151,n39152,n39153,n39154,n39155);
  nor U41353(n39155,n36897,n38298);
  nor U41354(n39154,n36896,n38299);
  nor U41355(n39153,n36895,n38300);
  nor U41356(n39152,n36889,n38301);
  nor U41357(n39150,n39156,n39157,n39158,n39159);
  nor U41358(n39159,n36888,n38306);
  nor U41359(n39158,n36887,n38307);
  nor U41360(n39157,n36881,n38308);
  nor U41361(n39156,n36880,n38309);
  nor U41362(n39149,n39160,n39161,n39162,n39163);
  nor U41363(n39163,n36879,n38314);
  nor U41364(n39162,n36873,n38315);
  nor U41365(n39161,n36872,n38316);
  nor U41366(n39160,n36871,n38317);
  nor U41367(n39148,n39164,n39165,n39166,n39167);
  nor U41368(n39167,n36898,n38322);
  nor U41369(n39166,n36890,n38323);
  nor U41370(n39165,n36882,n38324);
  nor U41371(n39164,n36874,n38325);
  and U41372(n39063,n39168,n39169,n39170,n39171);
  nand U41373(n39171,n34869,n36305);
  nor U41374(n39170,n39172,n39173);
  nor U41375(n39173,n34984,n36301);
  nor U41376(n39172,n36302,n39059);
  nand U41377(n39169,n36238,n35375);
  nand U41378(n39168,n34869,n36255);
  nand U41379(n39049,n39174,n39175);
  nand U41380(n39175,n36238,n39176);
  nand U41381(n39176,n39177,n39178);
  not U41382(n39177,n39179);
  nand U41383(n39050,n36234,n35375);
  nand U41384(G14507,n39180,n39181,n39182,n39183);
  nor U41385(n39183,n39184,n39060,n39185);
  nor U41386(n39185,n39057,n36288);
  nor U41387(n39060,G60016,n36226);
  nand U41388(n36226,n39186,n39187);
  nor U41389(n39184,n34982,n36233);
  nand U41390(n39182,n36235,n35400);
  xnor U41391(n35400,n36246,n39188);
  nor U41392(n39188,n39189,n39190);
  not U41393(n39190,n39174);
  nand U41394(n39174,n39191,n39179);
  nor U41395(n39189,n39191,n39179);
  nand U41396(n39179,n39192,n39193,n38712,n39194);
  nor U41397(n39194,n39195,n39196,n39197);
  nor U41398(n39197,n34982,n36301);
  nand U41399(n36301,n39198,n35692,n39199);
  nor U41400(n39196,n35386,n35781);
  nor U41401(n39195,n36302,n39057);
  nand U41402(n39193,n36238,n34938);
  nand U41403(n39192,n34884,n36255);
  not U41404(n36255,n36582);
  nor U41405(n36582,n38363,n38289);
  xnor U41406(n39191,n39178,n36246);
  nand U41407(n39178,n39202,n39203,n39204,n39205);
  nor U41408(n39205,n39200,n39201,n39206,n39207);
  nor U41409(n39207,n39208,n35781);
  nor U41410(n39208,n39209,n39210,n39211,n39212);
  nand U41411(n39212,n39213,n39214,n39215,n39216);
  nand U41412(n39216,n38841,G59885);
  not U41413(n38841,n38362);
  nand U41414(n38362,n39217,n39218);
  nand U41415(n39215,n38842,G59893);
  not U41416(n38842,n38361);
  nand U41417(n38361,n39217,n39219);
  nand U41418(n39214,n38843,G59901);
  not U41419(n38843,n38360);
  nand U41420(n38360,n39220,n39218);
  nand U41421(n39213,n38844,G59909);
  not U41422(n38844,n38359);
  nand U41423(n38359,n39220,n39219);
  nand U41424(n39211,n39221,n39222,n39223,n39224);
  nand U41425(n39224,n38849,G59917);
  not U41426(n38849,n38354);
  nand U41427(n38354,n39217,n39225);
  nand U41428(n39223,n38850,G59925);
  not U41429(n38850,n38353);
  nand U41430(n38353,n39217,n39226);
  nor U41431(n39217,n39227,n39228);
  nand U41432(n39222,n38851,G59933);
  not U41433(n38851,n38352);
  nand U41434(n38352,n39220,n39225);
  nand U41435(n39221,n38852,G59941);
  not U41436(n38852,n38351);
  nand U41437(n38351,n39220,n39226);
  nor U41438(n39220,n39229,n39227);
  nand U41439(n39210,n39230,n39231,n39232,n39233);
  nand U41440(n39233,n38857,G59949);
  not U41441(n38857,n38346);
  nand U41442(n38346,n39218,n39234);
  nand U41443(n39232,n38858,G59957);
  not U41444(n38858,n38345);
  nand U41445(n38345,n39219,n39234);
  nand U41446(n39231,n38859,G59965);
  not U41447(n38859,n38344);
  nand U41448(n38344,n39218,n39235);
  nor U41449(n39218,n39236,G60010);
  nand U41450(n39230,n38860,G59973);
  not U41451(n38860,n38343);
  nand U41452(n38343,n39219,n39235);
  nor U41453(n39219,n39236,n36985);
  nand U41454(n39209,n39237,n39238,n39239,n39240);
  nand U41455(n39240,n38865,G59981);
  not U41456(n38865,n38338);
  nand U41457(n38338,n39225,n39234);
  nand U41458(n39239,n38866,G59989);
  not U41459(n38866,n38337);
  nand U41460(n38337,n39226,n39234);
  and U41461(n39234,n39229,n39227);
  not U41462(n39229,n39228);
  nand U41463(n39238,n38867,G59997);
  not U41464(n38867,n38336);
  nand U41465(n38336,n39235,n39225);
  and U41466(n39225,n39236,n36985);
  nand U41467(n39237,n38868,G60005);
  not U41468(n38868,n38335);
  nand U41469(n38335,n39235,n39226);
  and U41470(n39226,G60010,n39236);
  and U41471(n39235,n39228,n39227);
  nor U41472(n39206,n39241,n39242,n39243,n39244);
  nand U41473(n39244,n36238,n39245,n39246,n39247);
  nand U41474(n39247,n39101,G59973);
  not U41475(n39101,n38261);
  nand U41476(n38261,n39248,n39249);
  nand U41477(n39246,n39102,G59941);
  not U41478(n39102,n38260);
  nand U41479(n38260,n39250,n39251);
  nand U41480(n39245,n39103,G59909);
  not U41481(n39103,n38262);
  nand U41482(n38262,n39251,n39249);
  nand U41483(n39243,n39252,n39253,n39254,n39255);
  nand U41484(n39255,n38265,G59901);
  not U41485(n38265,n38964);
  nand U41486(n38964,n39256,n39251);
  nand U41487(n39254,n38266,G59893);
  not U41488(n38266,n38969);
  nand U41489(n38969,n39257,n39249);
  nand U41490(n39253,n39108,G59885);
  not U41491(n39108,n38274);
  nand U41492(n38274,n39257,n39256);
  nand U41493(n39252,n39109,G60005);
  not U41494(n39109,n38273);
  nand U41495(n38273,n39250,n39248);
  nand U41496(n39242,n39258,n39259,n39260,n39261);
  nand U41497(n39261,n39114,G59949);
  not U41498(n39114,n38272);
  nand U41499(n38272,n39262,n39256);
  nand U41500(n39260,n39115,G59933);
  not U41501(n39115,n38271);
  nand U41502(n38271,n39263,n39251);
  nor U41503(n39251,n35350,n34869);
  nand U41504(n39259,n39116,G59925);
  not U41505(n39116,n38282);
  nand U41506(n38282,n39257,n39250);
  nand U41507(n39258,n39117,G59917);
  not U41508(n39117,n38281);
  nand U41509(n38281,n39263,n39257);
  nor U41510(n39257,n35374,n35350);
  not U41511(n35350,n34850);
  nand U41512(n39241,n39264,n39265,n39266,n39267);
  nor U41513(n39267,n39268,n39269);
  nor U41514(n39269,n36987,n38286);
  nand U41515(n38286,n39262,n39250);
  nor U41516(n39250,n34884,n34860);
  nor U41517(n39268,n36988,n38287);
  nand U41518(n38287,n39263,n39248);
  nand U41519(n39266,n39124,G59981);
  not U41520(n39124,n38288);
  nand U41521(n38288,n39263,n39262);
  nor U41522(n39263,n35386,n34860);
  nand U41523(n39265,n39125,G59957);
  not U41524(n39125,n38280);
  nand U41525(n38280,n39262,n39249);
  nor U41526(n39249,n34884,n35362);
  nor U41527(n39262,n35374,n34850);
  nand U41528(n39264,n39126,G59965);
  not U41529(n39126,n38279);
  nand U41530(n38279,n39256,n39248);
  nor U41531(n39248,n34869,n34850);
  nor U41532(n39256,n35362,n35386);
  not U41533(n35386,n34884);
  nand U41534(n39204,G60010,n35695);
  nand U41535(n39203,n38363,n39270);
  nand U41536(n39270,n39271,n39272,n39273,n39274);
  nor U41537(n39274,n39275,n39276,n39277,n39278);
  nor U41538(n39278,n36987,n38472);
  nor U41539(n39277,n36983,n38473);
  nor U41540(n39276,n36978,n38474);
  nor U41541(n39275,n36976,n38475);
  nor U41542(n39273,n39279,n39280,n39281,n39282);
  nor U41543(n39282,n36974,n38480);
  nor U41544(n39281,n36968,n38481);
  nor U41545(n39280,n36966,n38482);
  nor U41546(n39279,n36964,n38483);
  nor U41547(n39272,n39283,n39284,n39285,n39286);
  nor U41548(n39286,n36956,n38488);
  nor U41549(n39285,n36952,n38489);
  nor U41550(n39284,n36949,n38490);
  nor U41551(n39283,n36990,n38491);
  nor U41552(n39271,n39287,n39288,n39289,n39290);
  nor U41553(n39290,n36988,n38496);
  nor U41554(n39289,n36977,n38497);
  nor U41555(n39288,n36967,n38498);
  nor U41556(n39287,n36954,n38499);
  nand U41557(n39202,n38289,n37554);
  nand U41558(n37554,n39291,n39292,n39293,n39294);
  nor U41559(n39294,n39295,n39296,n39297,n39298);
  nor U41560(n39298,n36988,n38298);
  nand U41561(n38298,n39299,n39300);
  nor U41562(n39297,n36987,n38299);
  nand U41563(n38299,n39301,n39299);
  nor U41564(n39296,n36983,n38300);
  nand U41565(n38300,n39299,n39302);
  nor U41566(n39295,n36977,n38301);
  nand U41567(n38301,n39303,n39300);
  nor U41568(n39293,n39304,n39305,n39306,n39307);
  nor U41569(n39307,n36976,n38306);
  nand U41570(n38306,n39301,n39303);
  nor U41571(n39306,n36974,n38307);
  nand U41572(n38307,n39302,n39303);
  nor U41573(n39305,n36967,n38308);
  nand U41574(n38308,n39308,n39300);
  nor U41575(n39304,n36966,n38309);
  nand U41576(n38309,n39308,n39301);
  nor U41577(n39292,n39309,n39310,n39311,n39312);
  nor U41578(n39312,n36964,n38314);
  nand U41579(n38314,n39308,n39302);
  nor U41580(n39311,n36954,n38315);
  nand U41581(n38315,n39313,n39300);
  nor U41582(n39300,n39314,n35375);
  nor U41583(n39310,n36952,n38316);
  nand U41584(n38316,n39313,n39301);
  nor U41585(n39301,n34938,n36207);
  nor U41586(n39309,n36949,n38317);
  nand U41587(n38317,n39313,n39302);
  nor U41588(n39302,n36207,n39314);
  nor U41589(n39291,n39315,n39316,n39317,n39318);
  nor U41590(n39318,n36990,n38322);
  nand U41591(n38322,n39319,n39299);
  nor U41592(n39299,n35364,n35352);
  nor U41593(n39317,n36978,n38323);
  nand U41594(n38323,n39319,n39303);
  nor U41595(n39303,n36200,n35352);
  nor U41596(n39316,n36968,n38324);
  nand U41597(n38324,n39319,n39308);
  nor U41598(n39308,n36193,n35364);
  nor U41599(n39315,n36956,n38325);
  nand U41600(n38325,n39319,n39313);
  nor U41601(n39313,n36200,n36193);
  nor U41602(n39319,n34938,n35375);
  nor U41603(n38289,n34885,n35994,n39320);
  nand U41604(n39321,n39322,n39323,n39324,n39325);
  nand U41605(n39181,n36234,n34938);
  not U41606(n36234,n36726);
  nand U41607(n36726,n39186,n39326);
  nand U41608(n39326,n39327,n39328,n39329,n39330);
  nand U41609(n39180,n36272,n34884);
  not U41610(n36272,n37702);
  nand U41611(n37702,n39186,n39331);
  nand U41612(n39331,n39332,n39333,n39334,n39335);
  nor U41613(n39335,n39336,n39337);
  not U41614(n39333,n39338);
  nor U41615(n39186,n34898,n36231);
  not U41616(n36231,n36288);
  nand U41617(n36288,n35407,n39339);
  nand U41618(n39339,n34876,n39340);
  nand U41619(n39340,n39341,n39342,n39343,n39344);
  nand U41620(n39344,n38712,n35388,n39345);
  nand U41621(n39343,n39346,n34899);
  nand U41622(n39346,n39347,n39348);
  nand U41623(n39348,n39345,n39349,n39350);
  nand U41624(n39347,n39351,n34934);
  nand U41625(n39351,n39352,n39353);
  nand U41626(n39353,n39354,n35695);
  nand U41627(n39354,n34911,n34913);
  nand U41628(n39352,n39199,n34914);
  nand U41629(n39342,n34934,n39355);
  nand U41630(n35407,n34897,n35385,n34929);
  nand U41631(G14506,n39356,n39357,n39358);
  nand U41632(n39358,n34936,G60014);
  nand U41633(n39357,n34937,n35375);
  nand U41634(n39356,n34939,n34868);
  nand U41635(G14505,n39359,n39360,n39361);
  nand U41636(n39361,n34936,G60013);
  nand U41637(n39360,n34937,n35364);
  nand U41638(n39359,n34939,n34859);
  nand U41639(G14504,n39362,n39363,n39364);
  nand U41640(n39364,n34936,G60012);
  nand U41641(n39363,n34937,n35352);
  and U41642(n34937,n39365,n34935);
  nand U41643(n39365,n39366,n39367);
  nand U41644(n39367,n36215,n34898);
  nand U41645(n39362,n34939,n39368);
  nor U41646(n34939,n34936,G59875,n36215);
  not U41647(n34936,n34935);
  nor U41648(G14503,n39369,n34935);
  nand U41649(n34935,n39370,n34874,n39371);
  nand U41650(n34874,G60244,n39372);
  nand U41651(n39370,n34885,n39372);
  nand U41652(G14502,n39373,n39374,n39375,n39376);
  nor U41653(n39376,n39377,n39378,n39379);
  nor U41654(n39379,n35694,n39380);
  nor U41655(n39378,n39381,n39382);
  nor U41656(n39377,n37009,n39383);
  nand U41657(n39375,n39384,G60005);
  nand U41658(n39374,n39385,n39386);
  nand U41659(n39373,n35778,n39387);
  nand U41660(G14501,n39388,n39389,n39390,n39391);
  nor U41661(n39391,n39392,n39393,n39394);
  nor U41662(n39394,n35684,n39380);
  nor U41663(n39393,n39395,n39382);
  nor U41664(n39392,n37009,n39396);
  nand U41665(n39390,n39384,G60004);
  nand U41666(n39389,n39397,n39386);
  nand U41667(n39388,n35773,n39387);
  nand U41668(G14500,n39398,n39399,n39400,n39401);
  nor U41669(n39401,n39402,n39403,n39404);
  nor U41670(n39404,n35676,n39380);
  nor U41671(n39403,n39405,n39382);
  nor U41672(n39402,n37009,n39406);
  nand U41673(n39400,n39384,G60003);
  nand U41674(n39399,n39407,n39386);
  nand U41675(n39398,n35768,n39387);
  nand U41676(G14499,n39408,n39409,n39410,n39411);
  nor U41677(n39411,n39412,n39413,n39414);
  nor U41678(n39414,n35668,n39380);
  nor U41679(n39413,n39415,n39382);
  nor U41680(n39412,n37009,n39416);
  nand U41681(n39410,n39384,G60002);
  nand U41682(n39409,n39417,n39386);
  nand U41683(n39408,n35763,n39387);
  nand U41684(G14498,n39418,n39419,n39420,n39421);
  nor U41685(n39421,n39422,n39423,n39424);
  nor U41686(n39424,n35659,n39380);
  nor U41687(n39423,n39425,n39382);
  nor U41688(n39422,n37009,n39426);
  nand U41689(n39420,n39384,G60001);
  nand U41690(n39419,n39427,n39386);
  nand U41691(n39418,n35758,n39387);
  nand U41692(G14497,n39428,n39429,n39430,n39431);
  nor U41693(n39431,n39432,n39433,n39434);
  nor U41694(n39434,n35650,n39380);
  nor U41695(n39433,n39435,n39382);
  nor U41696(n39432,n37009,n39436);
  nand U41697(n39430,n39384,G60000);
  nand U41698(n39429,n39437,n39386);
  nand U41699(n39428,n35753,n39387);
  nand U41700(G14496,n39438,n39439,n39440,n39441);
  nor U41701(n39441,n39442,n39443,n39444);
  nor U41702(n39444,n35641,n39380);
  nor U41703(n39443,n39445,n39382);
  nor U41704(n39442,n37009,n39446);
  nand U41705(n39440,n39384,G59999);
  nand U41706(n39439,n39447,n39386);
  nand U41707(n39438,n35747,n39387);
  nand U41708(G14495,n39448,n39449,n39450,n39451);
  nor U41709(n39451,n39452,n39453,n39454);
  nor U41710(n39454,n35631,n39380);
  nand U41711(n39380,n39455,n37009,n39456);
  nor U41712(n39453,n39457,n39382);
  nor U41713(n39452,n37009,n39458);
  nand U41714(n39450,n39384,G59998);
  and U41715(n39384,n39459,n39460);
  nand U41716(n39460,n39461,n39462,n39463);
  nand U41717(n39463,G59875,n38491);
  nand U41718(n39461,n39464,n39465);
  nand U41719(n39459,n39466,n39467);
  nand U41720(n39449,n39468,n39386);
  nand U41721(n39386,n39469,n39470);
  or U41722(n39470,n39465,n36215);
  nand U41723(n39469,n39455,G59875);
  not U41724(n39455,n38491);
  nand U41725(n39448,n35742,n39387);
  nand U41726(n39387,n39471,n39472);
  nand U41727(n39472,n39466,n39464);
  nand U41728(n39464,n39473,n39474);
  not U41729(n39466,n39382);
  nand U41730(n39382,n39475,n39476);
  or U41731(n39471,n39474,n39465);
  nand U41732(n39465,n39477,n39478);
  nand U41733(n39474,n37009,n38491,n39456);
  nand U41734(n37009,n39479,n39480);
  nand U41735(G14494,n39481,n39482,n39483,n39484);
  nor U41736(n39484,n39485,n39486,n39487);
  nor U41737(n39487,n39488,n35691);
  nor U41738(n39486,n39489,n39490);
  nor U41739(n39485,n36988,n39491);
  nand U41740(n39483,n39492,n39493);
  nand U41741(n39482,n39494,n39495);
  nand U41742(n39481,n39496,n39497);
  nand U41743(G14493,n39498,n39499,n39500,n39501);
  nor U41744(n39501,n39502,n39503,n39504);
  nor U41745(n39504,n39488,n35683);
  nor U41746(n39503,n39489,n39505);
  nor U41747(n39502,n36897,n39491);
  nand U41748(n39500,n39492,n39506);
  nand U41749(n39499,n39507,n39495);
  nand U41750(n39498,n39496,n39508);
  nand U41751(G14492,n39509,n39510,n39511,n39512);
  nor U41752(n39512,n39513,n39514,n39515);
  nor U41753(n39515,n39488,n35675);
  nor U41754(n39514,n39489,n39516);
  nor U41755(n39513,n36801,n39491);
  nand U41756(n39511,n39492,n39517);
  nand U41757(n39510,n39518,n39495);
  nand U41758(n39509,n39496,n39519);
  nand U41759(G14491,n39520,n39521,n39522,n39523);
  nor U41760(n39523,n39524,n39525,n39526);
  nor U41761(n39526,n39488,n35667);
  nor U41762(n39525,n39489,n39527);
  nor U41763(n39524,n37344,n39491);
  nand U41764(n39522,n39492,n39528);
  nand U41765(n39521,n39529,n39495);
  nand U41766(n39520,n39496,n39530);
  nand U41767(G14490,n39531,n39532,n39533,n39534);
  nor U41768(n39534,n39535,n39536,n39537);
  nor U41769(n39537,n39488,n35658);
  nor U41770(n39536,n39489,n39538);
  nor U41771(n39535,n37261,n39491);
  nand U41772(n39533,n39492,n39539);
  nand U41773(n39532,n39540,n39495);
  nand U41774(n39531,n39496,n39541);
  nand U41775(G14489,n39542,n39543,n39544,n39545);
  nor U41776(n39545,n39546,n39547,n39548);
  nor U41777(n39548,n39488,n35649);
  nor U41778(n39547,n39489,n39549);
  nor U41779(n39546,n37179,n39491);
  nand U41780(n39544,n39492,n39550);
  nand U41781(n39543,n39551,n39495);
  nand U41782(n39542,n39496,n39552);
  nand U41783(G14488,n39553,n39554,n39555,n39556);
  nor U41784(n39556,n39557,n39558,n39559);
  nor U41785(n39559,n39488,n35640);
  nor U41786(n39558,n39489,n39560);
  nor U41787(n39557,n36479,n39491);
  nand U41788(n39555,n39492,n39561);
  nand U41789(n39554,n39562,n39495);
  nand U41790(n39553,n39496,n39563);
  nand U41791(G14487,n39564,n39565,n39566,n39567);
  nor U41792(n39567,n39568,n39569,n39570);
  nor U41793(n39570,n39488,n35630);
  and U41794(n39488,n39571,n39572);
  nand U41795(n39572,n39456,n39573,n37007,n38496);
  nand U41796(n39573,n39574,n39575);
  nand U41797(n39571,n39496,n39576);
  nor U41798(n39569,n39489,n39577);
  and U41799(n39489,n39578,n39579);
  or U41800(n39579,n39575,n36215);
  nand U41801(n39578,n39580,G59875);
  nor U41802(n39568,n37006,n39491);
  nand U41803(n39491,n39581,n39582);
  nand U41804(n39582,n39583,n39462,n39584);
  nand U41805(n39584,n39576,n39575);
  nand U41806(n39583,n39585,n38496);
  nand U41807(n39585,n39586,n34898);
  nand U41808(n39586,n39575,n37007);
  nand U41809(n39575,n39587,n39478);
  nand U41810(n39581,n39496,n39467);
  nand U41811(n39566,n39492,n39588);
  and U41812(n39492,n39456,n39580);
  not U41813(n39580,n38496);
  nand U41814(n39565,n39589,n39495);
  not U41815(n39495,n37007);
  nand U41816(n37007,n39590,n39480);
  nand U41817(n39564,n39496,n39591);
  not U41818(n39496,n39574);
  nand U41819(n39574,n39592,n39476);
  nand U41820(G14486,n39593,n39594,n39595,n39596);
  nor U41821(n39596,n39597,n39598,n39599);
  nor U41822(n39599,n35694,n39600);
  nor U41823(n39598,n39381,n39601);
  nor U41824(n39597,n37005,n39383);
  nand U41825(n39595,n39602,G59989);
  nand U41826(n39594,n39385,n39603);
  nand U41827(n39593,n35778,n39604);
  nand U41828(G14485,n39605,n39606,n39607,n39608);
  nor U41829(n39608,n39609,n39610,n39611);
  nor U41830(n39611,n35684,n39600);
  nor U41831(n39610,n39395,n39601);
  nor U41832(n39609,n37005,n39396);
  nand U41833(n39607,n39602,G59988);
  nand U41834(n39606,n39397,n39603);
  nand U41835(n39605,n35773,n39604);
  nand U41836(G14484,n39612,n39613,n39614,n39615);
  nor U41837(n39615,n39616,n39617,n39618);
  nor U41838(n39618,n35676,n39600);
  nor U41839(n39617,n39405,n39601);
  nor U41840(n39616,n37005,n39406);
  nand U41841(n39614,n39602,G59987);
  nand U41842(n39613,n39407,n39603);
  nand U41843(n39612,n35768,n39604);
  nand U41844(G14483,n39619,n39620,n39621,n39622);
  nor U41845(n39622,n39623,n39624,n39625);
  nor U41846(n39625,n35668,n39600);
  nor U41847(n39624,n39415,n39601);
  nor U41848(n39623,n37005,n39416);
  nand U41849(n39621,n39602,G59986);
  nand U41850(n39620,n39417,n39603);
  nand U41851(n39619,n35763,n39604);
  nand U41852(G14482,n39626,n39627,n39628,n39629);
  nor U41853(n39629,n39630,n39631,n39632);
  nor U41854(n39632,n35659,n39600);
  nor U41855(n39631,n39425,n39601);
  nor U41856(n39630,n37005,n39426);
  nand U41857(n39628,n39602,G59985);
  nand U41858(n39627,n39427,n39603);
  nand U41859(n39626,n35758,n39604);
  nand U41860(G14481,n39633,n39634,n39635,n39636);
  nor U41861(n39636,n39637,n39638,n39639);
  nor U41862(n39639,n35650,n39600);
  nor U41863(n39638,n39435,n39601);
  nor U41864(n39637,n37005,n39436);
  nand U41865(n39635,n39602,G59984);
  nand U41866(n39634,n39437,n39603);
  nand U41867(n39633,n35753,n39604);
  nand U41868(G14480,n39640,n39641,n39642,n39643);
  nor U41869(n39643,n39644,n39645,n39646);
  nor U41870(n39646,n35641,n39600);
  nor U41871(n39645,n39445,n39601);
  nor U41872(n39644,n37005,n39446);
  nand U41873(n39642,n39602,G59983);
  nand U41874(n39641,n39447,n39603);
  nand U41875(n39640,n35747,n39604);
  nand U41876(G14479,n39647,n39648,n39649,n39650);
  nor U41877(n39650,n39651,n39652,n39653);
  nor U41878(n39653,n35631,n39600);
  nand U41879(n39600,n39654,n37005,n39456);
  nor U41880(n39652,n39457,n39601);
  nor U41881(n39651,n37005,n39458);
  nand U41882(n39649,n39602,G59982);
  and U41883(n39602,n39655,n39656);
  nand U41884(n39656,n39657,n39462,n39658);
  nand U41885(n39658,G59875,n38472);
  nand U41886(n39657,n39659,n39660);
  nand U41887(n39655,n39661,n39467);
  nand U41888(n39648,n39468,n39603);
  nand U41889(n39603,n39662,n39663);
  or U41890(n39663,n39660,n36215);
  nand U41891(n39662,n39654,G59875);
  not U41892(n39654,n38472);
  nand U41893(n39647,n35742,n39604);
  nand U41894(n39604,n39664,n39665);
  nand U41895(n39665,n39661,n39659);
  nand U41896(n39659,n39473,n39666);
  not U41897(n39661,n39601);
  nand U41898(n39601,n39667,n39476);
  or U41899(n39664,n39666,n39660);
  nand U41900(n39660,n39668,n39478);
  nand U41901(n39666,n37005,n38472,n39456);
  nand U41902(n37005,n39669,n39479);
  nand U41903(G14478,n39670,n39671,n39672,n39673);
  nor U41904(n39673,n39674,n39675,n39676);
  nor U41905(n39676,n39381,n39677);
  nor U41906(n39675,n37003,n39383);
  nor U41907(n39674,n35694,n39678);
  nand U41908(n39672,n39679,G59981);
  nand U41909(n39671,n39385,n39680);
  nand U41910(n39670,n35778,n39681);
  nand U41911(G14477,n39682,n39683,n39684,n39685);
  nor U41912(n39685,n39686,n39687,n39688);
  nor U41913(n39688,n39395,n39677);
  nor U41914(n39687,n37003,n39396);
  nor U41915(n39686,n35684,n39678);
  nand U41916(n39684,n39679,G59980);
  nand U41917(n39683,n39397,n39680);
  nand U41918(n39682,n35773,n39681);
  nand U41919(G14476,n39689,n39690,n39691,n39692);
  nor U41920(n39692,n39693,n39694,n39695);
  nor U41921(n39695,n39405,n39677);
  nor U41922(n39694,n37003,n39406);
  nor U41923(n39693,n35676,n39678);
  nand U41924(n39691,n39679,G59979);
  nand U41925(n39690,n39407,n39680);
  nand U41926(n39689,n35768,n39681);
  nand U41927(G14475,n39696,n39697,n39698,n39699);
  nor U41928(n39699,n39700,n39701,n39702);
  nor U41929(n39702,n39415,n39677);
  nor U41930(n39701,n37003,n39416);
  nor U41931(n39700,n35668,n39678);
  nand U41932(n39698,n39679,G59978);
  nand U41933(n39697,n39417,n39680);
  nand U41934(n39696,n35763,n39681);
  nand U41935(G14474,n39703,n39704,n39705,n39706);
  nor U41936(n39706,n39707,n39708,n39709);
  nor U41937(n39709,n39425,n39677);
  nor U41938(n39708,n37003,n39426);
  nor U41939(n39707,n35659,n39678);
  nand U41940(n39705,n39679,G59977);
  nand U41941(n39704,n39427,n39680);
  nand U41942(n39703,n35758,n39681);
  nand U41943(G14473,n39710,n39711,n39712,n39713);
  nor U41944(n39713,n39714,n39715,n39716);
  nor U41945(n39716,n39435,n39677);
  nor U41946(n39715,n37003,n39436);
  nor U41947(n39714,n35650,n39678);
  nand U41948(n39712,n39679,G59976);
  nand U41949(n39711,n39437,n39680);
  nand U41950(n39710,n35753,n39681);
  nand U41951(G14472,n39717,n39718,n39719,n39720);
  nor U41952(n39720,n39721,n39722,n39723);
  nor U41953(n39723,n39445,n39677);
  nor U41954(n39722,n37003,n39446);
  nor U41955(n39721,n35641,n39678);
  nand U41956(n39719,n39679,G59975);
  nand U41957(n39718,n39447,n39680);
  nand U41958(n39717,n35747,n39681);
  nand U41959(G14471,n39724,n39725,n39726,n39727);
  nor U41960(n39727,n39728,n39729,n39730);
  nor U41961(n39730,n39457,n39677);
  nor U41962(n39729,n37003,n39458);
  nor U41963(n39728,n35631,n39678);
  nand U41964(n39678,n39456,n39731);
  nand U41965(n39726,n39679,G59974);
  and U41966(n39679,n39732,n39733);
  nand U41967(n39733,n39734,n39462,n39735);
  nand U41968(n39735,G59875,n38473);
  nand U41969(n39734,n39736,n39737);
  nand U41970(n39732,n39738,n39467);
  nand U41971(n39725,n39468,n39680);
  nand U41972(n39680,n39739,n39740);
  nand U41973(n39740,n39741,n36267);
  nand U41974(n39739,n39731,G59875);
  not U41975(n39731,n38473);
  nand U41976(n39724,n35742,n39681);
  nand U41977(n39681,n39742,n39743);
  nand U41978(n39743,n39456,n37003,n39741);
  not U41979(n39741,n39737);
  nand U41980(n39737,n39744,n39478);
  nor U41981(n39478,n39745,n39746);
  nand U41982(n39742,n39738,n39736);
  nand U41983(n39736,n39473,n39747);
  nand U41984(n39747,n37003,n38473,n39456);
  nand U41985(n37003,n39669,n39590);
  not U41986(n39738,n39677);
  nand U41987(n39677,n39476,n39748);
  nor U41988(n39476,G60013,G60012);
  nand U41989(G14470,n39749,n39750,n39751,n39752);
  nor U41990(n39752,n39753,n39754,n39755);
  nor U41991(n39755,n35694,n39756);
  nor U41992(n39754,n39381,n39757);
  nor U41993(n39753,n37021,n39383);
  nand U41994(n39751,n39758,G59973);
  nand U41995(n39750,n39385,n39759);
  nand U41996(n39749,n35778,n39760);
  nand U41997(G14469,n39761,n39762,n39763,n39764);
  nor U41998(n39764,n39765,n39766,n39767);
  nor U41999(n39767,n35684,n39756);
  nor U42000(n39766,n39395,n39757);
  nor U42001(n39765,n37021,n39396);
  nand U42002(n39763,n39758,G59972);
  nand U42003(n39762,n39397,n39759);
  nand U42004(n39761,n35773,n39760);
  nand U42005(G14468,n39768,n39769,n39770,n39771);
  nor U42006(n39771,n39772,n39773,n39774);
  nor U42007(n39774,n35676,n39756);
  nor U42008(n39773,n39405,n39757);
  nor U42009(n39772,n37021,n39406);
  nand U42010(n39770,n39758,G59971);
  nand U42011(n39769,n39407,n39759);
  nand U42012(n39768,n35768,n39760);
  nand U42013(G14467,n39775,n39776,n39777,n39778);
  nor U42014(n39778,n39779,n39780,n39781);
  nor U42015(n39781,n35668,n39756);
  nor U42016(n39780,n39415,n39757);
  nor U42017(n39779,n37021,n39416);
  nand U42018(n39777,n39758,G59970);
  nand U42019(n39776,n39417,n39759);
  nand U42020(n39775,n35763,n39760);
  nand U42021(G14466,n39782,n39783,n39784,n39785);
  nor U42022(n39785,n39786,n39787,n39788);
  nor U42023(n39788,n35659,n39756);
  nor U42024(n39787,n39425,n39757);
  nor U42025(n39786,n37021,n39426);
  nand U42026(n39784,n39758,G59969);
  nand U42027(n39783,n39427,n39759);
  nand U42028(n39782,n35758,n39760);
  nand U42029(G14465,n39789,n39790,n39791,n39792);
  nor U42030(n39792,n39793,n39794,n39795);
  nor U42031(n39795,n35650,n39756);
  nor U42032(n39794,n39435,n39757);
  nor U42033(n39793,n37021,n39436);
  nand U42034(n39791,n39758,G59968);
  nand U42035(n39790,n39437,n39759);
  nand U42036(n39789,n35753,n39760);
  nand U42037(G14464,n39796,n39797,n39798,n39799);
  nor U42038(n39799,n39800,n39801,n39802);
  nor U42039(n39802,n35641,n39756);
  nor U42040(n39801,n39445,n39757);
  nor U42041(n39800,n37021,n39446);
  nand U42042(n39798,n39758,G59967);
  nand U42043(n39797,n39447,n39759);
  nand U42044(n39796,n35747,n39760);
  nand U42045(G14463,n39803,n39804,n39805,n39806);
  nor U42046(n39806,n39807,n39808,n39809);
  nor U42047(n39809,n35631,n39756);
  nand U42048(n39756,n39810,n37021,n39456);
  nor U42049(n39808,n39457,n39757);
  nor U42050(n39807,n37021,n39458);
  nand U42051(n39805,n39758,G59966);
  and U42052(n39758,n39811,n39812);
  nand U42053(n39812,n39813,n39462,n39814);
  nand U42054(n39814,G59875,n38474);
  nand U42055(n39813,n39815,n39816);
  nand U42056(n39811,n39817,n39467);
  nand U42057(n39804,n39468,n39759);
  nand U42058(n39759,n39818,n39819);
  or U42059(n39819,n39816,n36215);
  nand U42060(n39818,n39810,G59875);
  not U42061(n39810,n38474);
  nand U42062(n39803,n35742,n39760);
  nand U42063(n39760,n39820,n39821);
  nand U42064(n39821,n39817,n39815);
  nand U42065(n39815,n39473,n39822);
  not U42066(n39817,n39757);
  nand U42067(n39757,n39475,n39823);
  or U42068(n39820,n39822,n39816);
  nand U42069(n39816,n39824,n39477);
  nand U42070(n39822,n37021,n38474,n39456);
  nand U42071(n37021,n39825,n39480);
  nand U42072(G14462,n39826,n39827,n39828,n39829);
  nor U42073(n39829,n39830,n39831,n39832);
  nor U42074(n39832,n39381,n39833);
  nor U42075(n39831,n37019,n39383);
  nor U42076(n39830,n35694,n39834);
  nand U42077(n39828,n39835,G59965);
  nand U42078(n39827,n39385,n39836);
  nand U42079(n39826,n35778,n39837);
  nand U42080(G14461,n39838,n39839,n39840,n39841);
  nor U42081(n39841,n39842,n39843,n39844);
  nor U42082(n39844,n39395,n39833);
  nor U42083(n39843,n37019,n39396);
  nor U42084(n39842,n35684,n39834);
  nand U42085(n39840,n39835,G59964);
  nand U42086(n39839,n39397,n39836);
  nand U42087(n39838,n35773,n39837);
  nand U42088(G14460,n39845,n39846,n39847,n39848);
  nor U42089(n39848,n39849,n39850,n39851);
  nor U42090(n39851,n39405,n39833);
  nor U42091(n39850,n37019,n39406);
  nor U42092(n39849,n35676,n39834);
  nand U42093(n39847,n39835,G59963);
  nand U42094(n39846,n39407,n39836);
  nand U42095(n39845,n35768,n39837);
  nand U42096(G14459,n39852,n39853,n39854,n39855);
  nor U42097(n39855,n39856,n39857,n39858);
  nor U42098(n39858,n39415,n39833);
  nor U42099(n39857,n37019,n39416);
  nor U42100(n39856,n35668,n39834);
  nand U42101(n39854,n39835,G59962);
  nand U42102(n39853,n39417,n39836);
  nand U42103(n39852,n35763,n39837);
  nand U42104(G14458,n39859,n39860,n39861,n39862);
  nor U42105(n39862,n39863,n39864,n39865);
  nor U42106(n39865,n39425,n39833);
  nor U42107(n39864,n37019,n39426);
  nor U42108(n39863,n35659,n39834);
  nand U42109(n39861,n39835,G59961);
  nand U42110(n39860,n39427,n39836);
  nand U42111(n39859,n35758,n39837);
  nand U42112(G14457,n39866,n39867,n39868,n39869);
  nor U42113(n39869,n39870,n39871,n39872);
  nor U42114(n39872,n39435,n39833);
  nor U42115(n39871,n37019,n39436);
  nor U42116(n39870,n35650,n39834);
  nand U42117(n39868,n39835,G59960);
  nand U42118(n39867,n39437,n39836);
  nand U42119(n39866,n35753,n39837);
  nand U42120(G14456,n39873,n39874,n39875,n39876);
  nor U42121(n39876,n39877,n39878,n39879);
  nor U42122(n39879,n39445,n39833);
  nor U42123(n39878,n37019,n39446);
  nor U42124(n39877,n35641,n39834);
  nand U42125(n39875,n39835,G59959);
  nand U42126(n39874,n39447,n39836);
  nand U42127(n39873,n35747,n39837);
  nand U42128(G14455,n39880,n39881,n39882,n39883);
  nor U42129(n39883,n39884,n39885,n39886);
  nor U42130(n39886,n39457,n39833);
  nor U42131(n39885,n37019,n39458);
  nor U42132(n39884,n35631,n39834);
  nand U42133(n39834,n39456,n39887);
  nand U42134(n39882,n39835,G59958);
  and U42135(n39835,n39888,n39889);
  nand U42136(n39889,n39890,n39462,n39891);
  nand U42137(n39891,G59875,n38497);
  nand U42138(n39890,n39892,n39893);
  nand U42139(n39888,n39894,n39467);
  nand U42140(n39881,n39468,n39836);
  nand U42141(n39836,n39895,n39896);
  nand U42142(n39896,n39897,n36267);
  nand U42143(n39895,n39887,G59875);
  not U42144(n39887,n38497);
  nand U42145(n39880,n35742,n39837);
  nand U42146(n39837,n39898,n39899);
  nand U42147(n39899,n39456,n37019,n39897);
  not U42148(n39897,n39893);
  nand U42149(n39893,n39824,n39587);
  nand U42150(n39898,n39894,n39892);
  nand U42151(n39892,n39473,n39900);
  nand U42152(n39900,n37019,n38497,n39456);
  nand U42153(n37019,n39901,n39480);
  nor U42154(n39480,n39902,n39903);
  not U42155(n39894,n39833);
  nand U42156(n39833,n39592,n39823);
  nand U42157(G14454,n39904,n39905,n39906,n39907);
  nor U42158(n39907,n39908,n39909,n39910);
  nor U42159(n39910,n35694,n39911);
  nor U42160(n39909,n39381,n39912);
  nor U42161(n39908,n37017,n39383);
  nand U42162(n39906,n39913,G59957);
  nand U42163(n39905,n39385,n39914);
  nand U42164(n39904,n35778,n39915);
  nand U42165(G14453,n39916,n39917,n39918,n39919);
  nor U42166(n39919,n39920,n39921,n39922);
  nor U42167(n39922,n35684,n39911);
  nor U42168(n39921,n39395,n39912);
  nor U42169(n39920,n37017,n39396);
  nand U42170(n39918,n39913,G59956);
  nand U42171(n39917,n39397,n39914);
  nand U42172(n39916,n35773,n39915);
  nand U42173(G14452,n39923,n39924,n39925,n39926);
  nor U42174(n39926,n39927,n39928,n39929);
  nor U42175(n39929,n35676,n39911);
  nor U42176(n39928,n39405,n39912);
  nor U42177(n39927,n37017,n39406);
  nand U42178(n39925,n39913,G59955);
  nand U42179(n39924,n39407,n39914);
  nand U42180(n39923,n35768,n39915);
  nand U42181(G14451,n39930,n39931,n39932,n39933);
  nor U42182(n39933,n39934,n39935,n39936);
  nor U42183(n39936,n35668,n39911);
  nor U42184(n39935,n39415,n39912);
  nor U42185(n39934,n37017,n39416);
  nand U42186(n39932,n39913,G59954);
  nand U42187(n39931,n39417,n39914);
  nand U42188(n39930,n35763,n39915);
  nand U42189(G14450,n39937,n39938,n39939,n39940);
  nor U42190(n39940,n39941,n39942,n39943);
  nor U42191(n39943,n35659,n39911);
  nor U42192(n39942,n39425,n39912);
  nor U42193(n39941,n37017,n39426);
  nand U42194(n39939,n39913,G59953);
  nand U42195(n39938,n39427,n39914);
  nand U42196(n39937,n35758,n39915);
  nand U42197(G14449,n39944,n39945,n39946,n39947);
  nor U42198(n39947,n39948,n39949,n39950);
  nor U42199(n39950,n35650,n39911);
  nor U42200(n39949,n39435,n39912);
  nor U42201(n39948,n37017,n39436);
  nand U42202(n39946,n39913,G59952);
  nand U42203(n39945,n39437,n39914);
  nand U42204(n39944,n35753,n39915);
  nand U42205(G14448,n39951,n39952,n39953,n39954);
  nor U42206(n39954,n39955,n39956,n39957);
  nor U42207(n39957,n35641,n39911);
  nor U42208(n39956,n39445,n39912);
  nor U42209(n39955,n37017,n39446);
  nand U42210(n39953,n39913,G59951);
  nand U42211(n39952,n39447,n39914);
  nand U42212(n39951,n35747,n39915);
  nand U42213(G14447,n39958,n39959,n39960,n39961);
  nor U42214(n39961,n39962,n39963,n39964);
  nor U42215(n39964,n35631,n39911);
  nand U42216(n39911,n39965,n37017,n39456);
  nor U42217(n39963,n39457,n39912);
  nor U42218(n39962,n37017,n39458);
  nand U42219(n39960,n39913,G59950);
  and U42220(n39913,n39966,n39967);
  nand U42221(n39967,n39968,n39462,n39969);
  nand U42222(n39969,G59875,n38475);
  nand U42223(n39968,n39970,n39971);
  nand U42224(n39966,n39972,n39467);
  nand U42225(n39959,n39468,n39914);
  nand U42226(n39914,n39973,n39974);
  or U42227(n39974,n39971,n36215);
  nand U42228(n39973,n39965,G59875);
  not U42229(n39965,n38475);
  nand U42230(n39958,n35742,n39915);
  nand U42231(n39915,n39975,n39976);
  nand U42232(n39976,n39972,n39970);
  nand U42233(n39970,n39473,n39977);
  not U42234(n39972,n39912);
  nand U42235(n39912,n39667,n39823);
  or U42236(n39975,n39977,n39971);
  nand U42237(n39971,n39824,n39668);
  nand U42238(n39977,n37017,n38475,n39456);
  nand U42239(n37017,n39825,n39669);
  nand U42240(G14446,n39978,n39979,n39980,n39981);
  nor U42241(n39981,n39982,n39983,n39984);
  nor U42242(n39984,n35694,n39985);
  nor U42243(n39983,n37015,n39383);
  nor U42244(n39982,n39381,n39986);
  nand U42245(n39980,n39987,G59949);
  nand U42246(n39979,n39385,n39988);
  nand U42247(n39978,n35778,n39989);
  nand U42248(G14445,n39990,n39991,n39992,n39993);
  nor U42249(n39993,n39994,n39995,n39996);
  nor U42250(n39996,n35684,n39985);
  nor U42251(n39995,n37015,n39396);
  nor U42252(n39994,n39395,n39986);
  nand U42253(n39992,n39987,G59948);
  nand U42254(n39991,n39397,n39988);
  nand U42255(n39990,n35773,n39989);
  nand U42256(G14444,n39997,n39998,n39999,n40000);
  nor U42257(n40000,n40001,n40002,n40003);
  nor U42258(n40003,n35676,n39985);
  nor U42259(n40002,n37015,n39406);
  nor U42260(n40001,n39405,n39986);
  nand U42261(n39999,n39987,G59947);
  nand U42262(n39998,n39407,n39988);
  nand U42263(n39997,n35768,n39989);
  nand U42264(G14443,n40004,n40005,n40006,n40007);
  nor U42265(n40007,n40008,n40009,n40010);
  nor U42266(n40010,n35668,n39985);
  nor U42267(n40009,n37015,n39416);
  nor U42268(n40008,n39415,n39986);
  nand U42269(n40006,n39987,G59946);
  nand U42270(n40005,n39417,n39988);
  nand U42271(n40004,n35763,n39989);
  nand U42272(G14442,n40011,n40012,n40013,n40014);
  nor U42273(n40014,n40015,n40016,n40017);
  nor U42274(n40017,n35659,n39985);
  nor U42275(n40016,n37015,n39426);
  nor U42276(n40015,n39425,n39986);
  nand U42277(n40013,n39987,G59945);
  nand U42278(n40012,n39427,n39988);
  nand U42279(n40011,n35758,n39989);
  nand U42280(G14441,n40018,n40019,n40020,n40021);
  nor U42281(n40021,n40022,n40023,n40024);
  nor U42282(n40024,n35650,n39985);
  nor U42283(n40023,n37015,n39436);
  nor U42284(n40022,n39435,n39986);
  nand U42285(n40020,n39987,G59944);
  nand U42286(n40019,n39437,n39988);
  nand U42287(n40018,n35753,n39989);
  nand U42288(G14440,n40025,n40026,n40027,n40028);
  nor U42289(n40028,n40029,n40030,n40031);
  nor U42290(n40031,n35641,n39985);
  nor U42291(n40030,n37015,n39446);
  nor U42292(n40029,n39445,n39986);
  nand U42293(n40027,n39987,G59943);
  nand U42294(n40026,n39447,n39988);
  nand U42295(n40025,n35747,n39989);
  nand U42296(G14439,n40032,n40033,n40034,n40035);
  nor U42297(n40035,n40036,n40037,n40038);
  nor U42298(n40038,n35631,n39985);
  nand U42299(n39985,n39456,n40039);
  nor U42300(n40037,n37015,n39458);
  nor U42301(n40036,n39457,n39986);
  nand U42302(n40034,n39987,G59942);
  and U42303(n39987,n40040,n40041);
  nand U42304(n40041,n40042,n39462,n40043);
  nand U42305(n40043,G59875,n38480);
  nand U42306(n40042,n40044,n40045);
  nand U42307(n40040,n40046,n39467);
  nand U42308(n40033,n39468,n39988);
  nand U42309(n39988,n40047,n40048);
  nand U42310(n40048,n40049,n36267);
  nand U42311(n40047,n40039,G59875);
  not U42312(n40039,n38480);
  nand U42313(n40032,n35742,n39989);
  nand U42314(n39989,n40050,n40051);
  nand U42315(n40051,n39456,n37015,n40049);
  not U42316(n40049,n40045);
  nand U42317(n40045,n39824,n39744);
  nor U42318(n39824,n39745,n40052);
  nand U42319(n40050,n40046,n40044);
  nand U42320(n40044,n39473,n40053);
  nand U42321(n40053,n37015,n38480,n39456);
  nand U42322(n37015,n39901,n39669);
  nor U42323(n39669,n39903,n40054);
  nand U42324(G14438,n40055,n40056,n40057,n40058);
  nor U42325(n40058,n40059,n40060,n40061);
  nor U42326(n40061,n35694,n40062);
  nor U42327(n40060,n39381,n40063);
  nor U42328(n40059,n37029,n39383);
  nand U42329(n40057,n40064,G59941);
  nand U42330(n40056,n39385,n40065);
  nand U42331(n40055,n35778,n40066);
  nand U42332(G14437,n40067,n40068,n40069,n40070);
  nor U42333(n40070,n40071,n40072,n40073);
  nor U42334(n40073,n35684,n40062);
  nor U42335(n40072,n39395,n40063);
  nor U42336(n40071,n37029,n39396);
  nand U42337(n40069,n40064,G59940);
  nand U42338(n40068,n39397,n40065);
  nand U42339(n40067,n35773,n40066);
  nand U42340(G14436,n40074,n40075,n40076,n40077);
  nor U42341(n40077,n40078,n40079,n40080);
  nor U42342(n40080,n35676,n40062);
  nor U42343(n40079,n39405,n40063);
  nor U42344(n40078,n37029,n39406);
  nand U42345(n40076,n40064,G59939);
  nand U42346(n40075,n39407,n40065);
  nand U42347(n40074,n35768,n40066);
  nand U42348(G14435,n40081,n40082,n40083,n40084);
  nor U42349(n40084,n40085,n40086,n40087);
  nor U42350(n40087,n35668,n40062);
  nor U42351(n40086,n39415,n40063);
  nor U42352(n40085,n37029,n39416);
  nand U42353(n40083,n40064,G59938);
  nand U42354(n40082,n39417,n40065);
  nand U42355(n40081,n35763,n40066);
  nand U42356(G14434,n40088,n40089,n40090,n40091);
  nor U42357(n40091,n40092,n40093,n40094);
  nor U42358(n40094,n35659,n40062);
  nor U42359(n40093,n39425,n40063);
  nor U42360(n40092,n37029,n39426);
  nand U42361(n40090,n40064,G59937);
  nand U42362(n40089,n39427,n40065);
  nand U42363(n40088,n35758,n40066);
  nand U42364(G14433,n40095,n40096,n40097,n40098);
  nor U42365(n40098,n40099,n40100,n40101);
  nor U42366(n40101,n35650,n40062);
  nor U42367(n40100,n39435,n40063);
  nor U42368(n40099,n37029,n39436);
  nand U42369(n40097,n40064,G59936);
  nand U42370(n40096,n39437,n40065);
  nand U42371(n40095,n35753,n40066);
  nand U42372(G14432,n40102,n40103,n40104,n40105);
  nor U42373(n40105,n40106,n40107,n40108);
  nor U42374(n40108,n35641,n40062);
  nor U42375(n40107,n39445,n40063);
  nor U42376(n40106,n37029,n39446);
  nand U42377(n40104,n40064,G59935);
  nand U42378(n40103,n39447,n40065);
  nand U42379(n40102,n35747,n40066);
  nand U42380(G14431,n40109,n40110,n40111,n40112);
  nor U42381(n40112,n40113,n40114,n40115);
  nor U42382(n40115,n35631,n40062);
  nand U42383(n40062,n40116,n37029,n39456);
  nor U42384(n40114,n39457,n40063);
  nor U42385(n40113,n37029,n39458);
  nand U42386(n40111,n40064,G59934);
  and U42387(n40064,n40117,n40118);
  nand U42388(n40118,n40119,n39462,n40120);
  nand U42389(n40120,G59875,n38481);
  nand U42390(n40119,n40121,n40122);
  nand U42391(n40117,n40123,n39467);
  nand U42392(n40110,n39468,n40065);
  nand U42393(n40065,n40124,n40125);
  or U42394(n40125,n40122,n36215);
  nand U42395(n40124,n40116,G59875);
  not U42396(n40116,n38481);
  nand U42397(n40109,n35742,n40066);
  nand U42398(n40066,n40126,n40127);
  nand U42399(n40127,n40123,n40121);
  nand U42400(n40121,n39473,n40128);
  not U42401(n40123,n40063);
  nand U42402(n40063,n40129,n39475);
  or U42403(n40126,n40128,n40122);
  nand U42404(n40122,n40130,n39477);
  nand U42405(n40128,n37029,n38481,n39456);
  nand U42406(n37029,n40131,n39479);
  nand U42407(G14430,n40132,n40133,n40134,n40135);
  nor U42408(n40135,n40136,n40137,n40138);
  nor U42409(n40138,n40139,n35691);
  nor U42410(n40137,n40140,n39490);
  nor U42411(n40136,n36967,n40141);
  nand U42412(n40134,n40142,n39493);
  nand U42413(n40133,n39494,n40143);
  nand U42414(n40132,n40144,n39497);
  nand U42415(G14429,n40145,n40146,n40147,n40148);
  nor U42416(n40148,n40149,n40150,n40151);
  nor U42417(n40151,n40139,n35683);
  nor U42418(n40150,n40140,n39505);
  nor U42419(n40149,n36881,n40141);
  nand U42420(n40147,n40142,n39506);
  nand U42421(n40146,n39507,n40143);
  nand U42422(n40145,n40144,n39508);
  nand U42423(G14428,n40152,n40153,n40154,n40155);
  nor U42424(n40155,n40156,n40157,n40158);
  nor U42425(n40158,n40139,n35675);
  nor U42426(n40157,n40140,n39516);
  nor U42427(n40156,n36785,n40141);
  nand U42428(n40154,n40142,n39517);
  nand U42429(n40153,n39518,n40143);
  nand U42430(n40152,n40144,n39519);
  nand U42431(G14427,n40159,n40160,n40161,n40162);
  nor U42432(n40162,n40163,n40164,n40165);
  nor U42433(n40165,n40139,n35667);
  nor U42434(n40164,n40140,n39527);
  nor U42435(n40163,n36716,n40141);
  nand U42436(n40161,n40142,n39528);
  nand U42437(n40160,n39529,n40143);
  nand U42438(n40159,n40144,n39530);
  nand U42439(G14426,n40166,n40167,n40168,n40169);
  nor U42440(n40169,n40170,n40171,n40172);
  nor U42441(n40172,n40139,n35658);
  nor U42442(n40171,n40140,n39538);
  nor U42443(n40170,n36640,n40141);
  nand U42444(n40168,n40142,n39539);
  nand U42445(n40167,n39540,n40143);
  nand U42446(n40166,n40144,n39541);
  nand U42447(G14425,n40173,n40174,n40175,n40176);
  nor U42448(n40176,n40177,n40178,n40179);
  nor U42449(n40179,n40139,n35649);
  nor U42450(n40178,n40140,n39549);
  nor U42451(n40177,n36561,n40141);
  nand U42452(n40175,n40142,n39550);
  nand U42453(n40174,n39551,n40143);
  nand U42454(n40173,n40144,n39552);
  nand U42455(G14424,n40180,n40181,n40182,n40183);
  nor U42456(n40183,n40184,n40185,n40186);
  nor U42457(n40186,n40139,n35640);
  nor U42458(n40185,n40140,n39560);
  nor U42459(n40184,n36457,n40141);
  nand U42460(n40182,n40142,n39561);
  nand U42461(n40181,n39562,n40143);
  nand U42462(n40180,n40144,n39563);
  nand U42463(G14423,n40187,n40188,n40189,n40190);
  nor U42464(n40190,n40191,n40192,n40193);
  nor U42465(n40193,n40139,n35630);
  and U42466(n40139,n40194,n40195);
  nand U42467(n40195,n39456,n40196,n37028,n38498);
  nand U42468(n40196,n40197,n40198);
  nand U42469(n40194,n40144,n39576);
  nor U42470(n40192,n40140,n39577);
  and U42471(n40140,n40199,n40200);
  or U42472(n40200,n40198,n36215);
  nand U42473(n40199,n40201,G59875);
  nor U42474(n40191,n36386,n40141);
  nand U42475(n40141,n40202,n40203);
  nand U42476(n40203,n40204,n39462,n40205);
  nand U42477(n40205,n39576,n40198);
  nand U42478(n40204,n40206,n38498);
  nand U42479(n40206,n40207,n34898);
  nand U42480(n40207,n40198,n37028);
  nand U42481(n40198,n40130,n39587);
  nand U42482(n40202,n40144,n39467);
  nand U42483(n40189,n40142,n39588);
  and U42484(n40142,n39456,n40201);
  not U42485(n40201,n38498);
  nand U42486(n40188,n39589,n40143);
  not U42487(n40143,n37028);
  nand U42488(n37028,n40131,n39590);
  nand U42489(n40187,n40144,n39591);
  not U42490(n40144,n40197);
  nand U42491(n40197,n40129,n39592);
  nand U42492(G14422,n40208,n40209,n40210,n40211);
  nor U42493(n40211,n40212,n40213,n40214);
  nor U42494(n40214,n35694,n40215);
  nor U42495(n40213,n39381,n40216);
  nor U42496(n40212,n37027,n39383);
  nand U42497(n40210,n40217,G59925);
  nand U42498(n40209,n39385,n40218);
  nand U42499(n40208,n35778,n40219);
  nand U42500(G14421,n40220,n40221,n40222,n40223);
  nor U42501(n40223,n40224,n40225,n40226);
  nor U42502(n40226,n35684,n40215);
  nor U42503(n40225,n39395,n40216);
  nor U42504(n40224,n37027,n39396);
  nand U42505(n40222,n40217,G59924);
  nand U42506(n40221,n39397,n40218);
  nand U42507(n40220,n35773,n40219);
  nand U42508(G14420,n40227,n40228,n40229,n40230);
  nor U42509(n40230,n40231,n40232,n40233);
  nor U42510(n40233,n35676,n40215);
  nor U42511(n40232,n39405,n40216);
  nor U42512(n40231,n37027,n39406);
  nand U42513(n40229,n40217,G59923);
  nand U42514(n40228,n39407,n40218);
  nand U42515(n40227,n35768,n40219);
  nand U42516(G14419,n40234,n40235,n40236,n40237);
  nor U42517(n40237,n40238,n40239,n40240);
  nor U42518(n40240,n35668,n40215);
  nor U42519(n40239,n39415,n40216);
  nor U42520(n40238,n37027,n39416);
  nand U42521(n40236,n40217,G59922);
  nand U42522(n40235,n39417,n40218);
  nand U42523(n40234,n35763,n40219);
  nand U42524(G14418,n40241,n40242,n40243,n40244);
  nor U42525(n40244,n40245,n40246,n40247);
  nor U42526(n40247,n35659,n40215);
  nor U42527(n40246,n39425,n40216);
  nor U42528(n40245,n37027,n39426);
  nand U42529(n40243,n40217,G59921);
  nand U42530(n40242,n39427,n40218);
  nand U42531(n40241,n35758,n40219);
  nand U42532(G14417,n40248,n40249,n40250,n40251);
  nor U42533(n40251,n40252,n40253,n40254);
  nor U42534(n40254,n35650,n40215);
  nor U42535(n40253,n39435,n40216);
  nor U42536(n40252,n37027,n39436);
  nand U42537(n40250,n40217,G59920);
  nand U42538(n40249,n39437,n40218);
  nand U42539(n40248,n35753,n40219);
  nand U42540(G14416,n40255,n40256,n40257,n40258);
  nor U42541(n40258,n40259,n40260,n40261);
  nor U42542(n40261,n35641,n40215);
  nor U42543(n40260,n39445,n40216);
  nor U42544(n40259,n37027,n39446);
  nand U42545(n40257,n40217,G59919);
  nand U42546(n40256,n39447,n40218);
  nand U42547(n40255,n35747,n40219);
  nand U42548(G14415,n40262,n40263,n40264,n40265);
  nor U42549(n40265,n40266,n40267,n40268);
  nor U42550(n40268,n35631,n40215);
  nand U42551(n40215,n40269,n37027,n39456);
  nor U42552(n40267,n39457,n40216);
  nor U42553(n40266,n37027,n39458);
  nand U42554(n40264,n40217,G59918);
  and U42555(n40217,n40270,n40271);
  nand U42556(n40271,n40272,n39462,n40273);
  nand U42557(n40273,G59875,n38482);
  nand U42558(n40272,n40274,n40275);
  nand U42559(n40270,n40276,n39467);
  nand U42560(n40263,n39468,n40218);
  nand U42561(n40218,n40277,n40278);
  or U42562(n40278,n40275,n36215);
  nand U42563(n40277,n40269,G59875);
  not U42564(n40269,n38482);
  nand U42565(n40262,n35742,n40219);
  nand U42566(n40219,n40279,n40280);
  nand U42567(n40280,n40276,n40274);
  nand U42568(n40274,n39473,n40281);
  not U42569(n40276,n40216);
  nand U42570(n40216,n40129,n39667);
  or U42571(n40279,n40281,n40275);
  nand U42572(n40275,n40130,n39668);
  nand U42573(n40281,n37027,n38482,n39456);
  nand U42574(n37027,n40282,n39479);
  and U42575(n39479,n40283,n40284);
  nand U42576(G14414,n40285,n40286,n40287,n40288);
  nor U42577(n40288,n40289,n40290,n40291);
  nor U42578(n40291,n39381,n40292);
  nor U42579(n40290,n37026,n39383);
  nor U42580(n40289,n35694,n40293);
  nand U42581(n40287,n40294,G59917);
  nand U42582(n40286,n39385,n40295);
  nand U42583(n40285,n35778,n40296);
  nand U42584(G14413,n40297,n40298,n40299,n40300);
  nor U42585(n40300,n40301,n40302,n40303);
  nor U42586(n40303,n39395,n40292);
  nor U42587(n40302,n37026,n39396);
  nor U42588(n40301,n35684,n40293);
  nand U42589(n40299,n40294,G59916);
  nand U42590(n40298,n39397,n40295);
  nand U42591(n40297,n35773,n40296);
  nand U42592(G14412,n40304,n40305,n40306,n40307);
  nor U42593(n40307,n40308,n40309,n40310);
  nor U42594(n40310,n39405,n40292);
  nor U42595(n40309,n37026,n39406);
  nor U42596(n40308,n35676,n40293);
  nand U42597(n40306,n40294,G59915);
  nand U42598(n40305,n39407,n40295);
  nand U42599(n40304,n35768,n40296);
  nand U42600(G14411,n40311,n40312,n40313,n40314);
  nor U42601(n40314,n40315,n40316,n40317);
  nor U42602(n40317,n39415,n40292);
  nor U42603(n40316,n37026,n39416);
  nor U42604(n40315,n35668,n40293);
  nand U42605(n40313,n40294,G59914);
  nand U42606(n40312,n39417,n40295);
  nand U42607(n40311,n35763,n40296);
  nand U42608(G14410,n40318,n40319,n40320,n40321);
  nor U42609(n40321,n40322,n40323,n40324);
  nor U42610(n40324,n39425,n40292);
  nor U42611(n40323,n37026,n39426);
  nor U42612(n40322,n35659,n40293);
  nand U42613(n40320,n40294,G59913);
  nand U42614(n40319,n39427,n40295);
  nand U42615(n40318,n35758,n40296);
  nand U42616(G14409,n40325,n40326,n40327,n40328);
  nor U42617(n40328,n40329,n40330,n40331);
  nor U42618(n40331,n39435,n40292);
  nor U42619(n40330,n37026,n39436);
  nor U42620(n40329,n35650,n40293);
  nand U42621(n40327,n40294,G59912);
  nand U42622(n40326,n39437,n40295);
  nand U42623(n40325,n35753,n40296);
  nand U42624(G14408,n40332,n40333,n40334,n40335);
  nor U42625(n40335,n40336,n40337,n40338);
  nor U42626(n40338,n39445,n40292);
  nor U42627(n40337,n37026,n39446);
  nor U42628(n40336,n35641,n40293);
  nand U42629(n40334,n40294,G59911);
  nand U42630(n40333,n39447,n40295);
  nand U42631(n40332,n35747,n40296);
  nand U42632(G14407,n40339,n40340,n40341,n40342);
  nor U42633(n40342,n40343,n40344,n40345);
  nor U42634(n40345,n39457,n40292);
  nor U42635(n40344,n37026,n39458);
  nor U42636(n40343,n35631,n40293);
  nand U42637(n40293,n39456,n40346);
  nand U42638(n40341,n40294,G59910);
  and U42639(n40294,n40347,n40348);
  nand U42640(n40348,n40349,n39462,n40350);
  nand U42641(n40350,G59875,n38483);
  nand U42642(n40349,n40351,n40352);
  nand U42643(n40347,n40353,n39467);
  nand U42644(n40340,n39468,n40295);
  nand U42645(n40295,n40354,n40355);
  nand U42646(n40355,n40356,n36267);
  nand U42647(n40354,n40346,G59875);
  not U42648(n40346,n38483);
  nand U42649(n40339,n35742,n40296);
  nand U42650(n40296,n40357,n40358);
  nand U42651(n40358,n39456,n37026,n40356);
  not U42652(n40356,n40352);
  nand U42653(n40352,n40130,n39744);
  nor U42654(n40130,n39746,n40359);
  nand U42655(n40357,n40353,n40351);
  nand U42656(n40351,n39473,n40360);
  nand U42657(n40360,n37026,n38483,n39456);
  nand U42658(n37026,n40282,n39590);
  and U42659(n39590,n40361,n40283);
  not U42660(n40353,n40292);
  nand U42661(n40292,n40129,n39748);
  nand U42662(G14406,n40362,n40363,n40364,n40365);
  nor U42663(n40365,n40366,n40367,n40368);
  nor U42664(n40368,n35694,n40369);
  nor U42665(n40367,n39381,n40370);
  nor U42666(n40366,n37037,n39383);
  nand U42667(n40364,n40371,G59909);
  nand U42668(n40363,n39385,n40372);
  nand U42669(n40362,n35778,n40373);
  nand U42670(G14405,n40374,n40375,n40376,n40377);
  nor U42671(n40377,n40378,n40379,n40380);
  nor U42672(n40380,n35684,n40369);
  nor U42673(n40379,n39395,n40370);
  nor U42674(n40378,n37037,n39396);
  nand U42675(n40376,n40371,G59908);
  nand U42676(n40375,n39397,n40372);
  nand U42677(n40374,n35773,n40373);
  nand U42678(G14404,n40381,n40382,n40383,n40384);
  nor U42679(n40384,n40385,n40386,n40387);
  nor U42680(n40387,n35676,n40369);
  nor U42681(n40386,n39405,n40370);
  nor U42682(n40385,n37037,n39406);
  nand U42683(n40383,n40371,G59907);
  nand U42684(n40382,n39407,n40372);
  nand U42685(n40381,n35768,n40373);
  nand U42686(G14403,n40388,n40389,n40390,n40391);
  nor U42687(n40391,n40392,n40393,n40394);
  nor U42688(n40394,n35668,n40369);
  nor U42689(n40393,n39415,n40370);
  nor U42690(n40392,n37037,n39416);
  nand U42691(n40390,n40371,G59906);
  nand U42692(n40389,n39417,n40372);
  nand U42693(n40388,n35763,n40373);
  nand U42694(G14402,n40395,n40396,n40397,n40398);
  nor U42695(n40398,n40399,n40400,n40401);
  nor U42696(n40401,n35659,n40369);
  nor U42697(n40400,n39425,n40370);
  nor U42698(n40399,n37037,n39426);
  nand U42699(n40397,n40371,G59905);
  nand U42700(n40396,n39427,n40372);
  nand U42701(n40395,n35758,n40373);
  nand U42702(G14401,n40402,n40403,n40404,n40405);
  nor U42703(n40405,n40406,n40407,n40408);
  nor U42704(n40408,n35650,n40369);
  nor U42705(n40407,n39435,n40370);
  nor U42706(n40406,n37037,n39436);
  nand U42707(n40404,n40371,G59904);
  nand U42708(n40403,n39437,n40372);
  nand U42709(n40402,n35753,n40373);
  nand U42710(G14400,n40409,n40410,n40411,n40412);
  nor U42711(n40412,n40413,n40414,n40415);
  nor U42712(n40415,n35641,n40369);
  nor U42713(n40414,n39445,n40370);
  nor U42714(n40413,n37037,n39446);
  nand U42715(n40411,n40371,G59903);
  nand U42716(n40410,n39447,n40372);
  nand U42717(n40409,n35747,n40373);
  nand U42718(G14399,n40416,n40417,n40418,n40419);
  nor U42719(n40419,n40420,n40421,n40422);
  nor U42720(n40422,n35631,n40369);
  nand U42721(n40369,n40423,n37037,n39456);
  nor U42722(n40421,n39457,n40370);
  nor U42723(n40420,n37037,n39458);
  nand U42724(n40418,n40371,G59902);
  and U42725(n40371,n40424,n40425);
  nand U42726(n40425,n40426,n39462,n40427);
  nand U42727(n40427,G59875,n38488);
  nand U42728(n40426,n40428,n40429);
  nand U42729(n40424,n40430,n39467);
  nand U42730(n40417,n39468,n40372);
  nand U42731(n40372,n40431,n40432);
  or U42732(n40432,n40429,n36215);
  nand U42733(n40431,n40423,G59875);
  not U42734(n40423,n38488);
  nand U42735(n40416,n35742,n40373);
  nand U42736(n40373,n40433,n40434);
  nand U42737(n40434,n40430,n40428);
  nand U42738(n40428,n39473,n40435);
  not U42739(n40430,n40370);
  nand U42740(n40370,n40436,n39475);
  nor U42741(n39475,G60015,G60014);
  or U42742(n40433,n40435,n40429);
  nand U42743(n40429,n40437,n39477);
  nor U42744(n39477,n40438,n40439);
  nand U42745(n40435,n37037,n38488,n39456);
  nand U42746(n37037,n40131,n39825);
  nand U42747(G14398,n40440,n40441,n40442,n40443);
  nor U42748(n40443,n40444,n40445,n40446);
  nor U42749(n40446,n40447,n35691);
  nor U42750(n40445,n40448,n39490);
  nor U42751(n40444,n36954,n40449);
  nand U42752(n40442,n40450,n39493);
  nand U42753(n40441,n39494,n40451);
  nand U42754(n40440,n40452,n39497);
  nand U42755(G14397,n40453,n40454,n40455,n40456);
  nor U42756(n40456,n40457,n40458,n40459);
  nor U42757(n40459,n40447,n35683);
  nor U42758(n40458,n40448,n39505);
  nor U42759(n40457,n36873,n40449);
  nand U42760(n40455,n40450,n39506);
  nand U42761(n40454,n39507,n40451);
  nand U42762(n40453,n40452,n39508);
  nand U42763(G14396,n40460,n40461,n40462,n40463);
  nor U42764(n40463,n40464,n40465,n40466);
  nor U42765(n40466,n40447,n35675);
  nor U42766(n40465,n40448,n39516);
  nor U42767(n40464,n36777,n40449);
  nand U42768(n40462,n40450,n39517);
  nand U42769(n40461,n39518,n40451);
  nand U42770(n40460,n40452,n39519);
  nand U42771(G14395,n40467,n40468,n40469,n40470);
  nor U42772(n40470,n40471,n40472,n40473);
  nor U42773(n40473,n40447,n35667);
  nor U42774(n40472,n40448,n39527);
  nor U42775(n40471,n36708,n40449);
  nand U42776(n40469,n40450,n39528);
  nand U42777(n40468,n39529,n40451);
  nand U42778(n40467,n40452,n39530);
  nand U42779(G14394,n40474,n40475,n40476,n40477);
  nor U42780(n40477,n40478,n40479,n40480);
  nor U42781(n40480,n40447,n35658);
  nor U42782(n40479,n40448,n39538);
  nor U42783(n40478,n36632,n40449);
  nand U42784(n40476,n40450,n39539);
  nand U42785(n40475,n39540,n40451);
  nand U42786(n40474,n40452,n39541);
  nand U42787(G14393,n40481,n40482,n40483,n40484);
  nor U42788(n40484,n40485,n40486,n40487);
  nor U42789(n40487,n40447,n35649);
  nor U42790(n40486,n40448,n39549);
  nor U42791(n40485,n36553,n40449);
  nand U42792(n40483,n40450,n39550);
  nand U42793(n40482,n39551,n40451);
  nand U42794(n40481,n40452,n39552);
  nand U42795(G14392,n40488,n40489,n40490,n40491);
  nor U42796(n40491,n40492,n40493,n40494);
  nor U42797(n40494,n40447,n35640);
  nor U42798(n40493,n40448,n39560);
  nor U42799(n40492,n36449,n40449);
  nand U42800(n40490,n40450,n39561);
  nand U42801(n40489,n39562,n40451);
  nand U42802(n40488,n40452,n39563);
  nand U42803(G14391,n40495,n40496,n40497,n40498);
  nor U42804(n40498,n40499,n40500,n40501);
  nor U42805(n40501,n40447,n35630);
  and U42806(n40447,n40502,n40503);
  nand U42807(n40503,n39456,n40504,n37036,n38499);
  nand U42808(n40504,n40505,n40506);
  nand U42809(n40502,n40452,n39576);
  nor U42810(n40500,n40448,n39577);
  and U42811(n40448,n40507,n40508);
  or U42812(n40508,n40506,n36215);
  nand U42813(n40507,n40509,G59875);
  nor U42814(n40499,n36374,n40449);
  nand U42815(n40449,n40510,n40511);
  nand U42816(n40511,n40512,n39462,n40513);
  nand U42817(n40513,n39576,n40506);
  nand U42818(n40512,n40514,n38499);
  nand U42819(n40514,n40515,n34898);
  nand U42820(n40515,n40506,n37036);
  nand U42821(n40506,n40437,n39587);
  nor U42822(n39587,n40438,G60015);
  nand U42823(n40510,n40452,n39467);
  nand U42824(n40497,n40450,n39588);
  and U42825(n40450,n39456,n40509);
  not U42826(n40509,n38499);
  nand U42827(n40496,n39589,n40451);
  not U42828(n40451,n37036);
  nand U42829(n37036,n40131,n39901);
  nor U42830(n40131,n39902,n40516);
  not U42831(n39589,n39458);
  nand U42832(n40495,n40452,n39591);
  not U42833(n40452,n40505);
  nand U42834(n40505,n40436,n39592);
  nand U42835(G14390,n40517,n40518,n40519,n40520);
  nor U42836(n40520,n40521,n40522,n40523);
  nor U42837(n40523,n35694,n40524);
  nor U42838(n40522,n39381,n40525);
  nor U42839(n40521,n37035,n39383);
  nand U42840(n40519,n40526,G59893);
  nand U42841(n40518,n39385,n40527);
  nand U42842(n40517,n35778,n40528);
  nand U42843(G14389,n40529,n40530,n40531,n40532);
  nor U42844(n40532,n40533,n40534,n40535);
  nor U42845(n40535,n35684,n40524);
  nor U42846(n40534,n39395,n40525);
  nor U42847(n40533,n37035,n39396);
  nand U42848(n40531,n40526,G59892);
  nand U42849(n40530,n39397,n40527);
  nand U42850(n40529,n35773,n40528);
  nand U42851(G14388,n40536,n40537,n40538,n40539);
  nor U42852(n40539,n40540,n40541,n40542);
  nor U42853(n40542,n35676,n40524);
  nor U42854(n40541,n39405,n40525);
  nor U42855(n40540,n37035,n39406);
  nand U42856(n40538,n40526,G59891);
  nand U42857(n40537,n39407,n40527);
  nand U42858(n40536,n35768,n40528);
  nand U42859(G14387,n40543,n40544,n40545,n40546);
  nor U42860(n40546,n40547,n40548,n40549);
  nor U42861(n40549,n35668,n40524);
  nor U42862(n40548,n39415,n40525);
  nor U42863(n40547,n37035,n39416);
  nand U42864(n40545,n40526,G59890);
  nand U42865(n40544,n39417,n40527);
  nand U42866(n40543,n35763,n40528);
  nand U42867(G14386,n40550,n40551,n40552,n40553);
  nor U42868(n40553,n40554,n40555,n40556);
  nor U42869(n40556,n35659,n40524);
  nor U42870(n40555,n39425,n40525);
  nor U42871(n40554,n37035,n39426);
  nand U42872(n40552,n40526,G59889);
  nand U42873(n40551,n39427,n40527);
  nand U42874(n40550,n35758,n40528);
  nand U42875(G14385,n40557,n40558,n40559,n40560);
  nor U42876(n40560,n40561,n40562,n40563);
  nor U42877(n40563,n35650,n40524);
  nor U42878(n40562,n39435,n40525);
  nor U42879(n40561,n37035,n39436);
  nand U42880(n40559,n40526,G59888);
  nand U42881(n40558,n39437,n40527);
  nand U42882(n40557,n35753,n40528);
  nand U42883(G14384,n40564,n40565,n40566,n40567);
  nor U42884(n40567,n40568,n40569,n40570);
  nor U42885(n40570,n35641,n40524);
  nor U42886(n40569,n39445,n40525);
  nor U42887(n40568,n37035,n39446);
  nand U42888(n40566,n40526,G59887);
  nand U42889(n40565,n39447,n40527);
  nand U42890(n40564,n35747,n40528);
  nand U42891(G14383,n40571,n40572,n40573,n40574);
  nor U42892(n40574,n40575,n40576,n40577);
  nor U42893(n40577,n35631,n40524);
  nand U42894(n40524,n40578,n37035,n39456);
  nor U42895(n40576,n39457,n40525);
  nor U42896(n40575,n37035,n39458);
  nand U42897(n40573,n40526,G59886);
  and U42898(n40526,n40579,n40580);
  nand U42899(n40580,n40581,n39462,n40582);
  nand U42900(n40582,G59875,n38489);
  nand U42901(n40581,n40583,n40584);
  nand U42902(n40579,n40585,n39467);
  nand U42903(n40572,n39468,n40527);
  nand U42904(n40527,n40586,n40587);
  or U42905(n40587,n40584,n36215);
  nand U42906(n40586,n40578,G59875);
  not U42907(n40578,n38489);
  nand U42908(n40571,n35742,n40528);
  nand U42909(n40528,n40588,n40589);
  nand U42910(n40589,n40585,n40583);
  nand U42911(n40583,n39473,n40590);
  not U42912(n40585,n40525);
  nand U42913(n40525,n40436,n39667);
  or U42914(n40588,n40590,n40584);
  nand U42915(n40584,n40437,n39668);
  nor U42916(n39668,n40439,n40591);
  nand U42917(n40590,n37035,n38489,n39456);
  nand U42918(n37035,n40282,n39825);
  nor U42919(n39825,n40283,n40361);
  nand U42920(G14382,n40592,n40593,n40594,n40595);
  nor U42921(n40595,n40596,n40597,n40598);
  nor U42922(n40598,n35694,n40599);
  not U42923(n35694,n39493);
  nor U42924(n39493,n40600,n40601);
  nor U42925(n40601,G16,n34805);
  nor U42926(n40600,G58855,n35621);
  nor U42927(n40597,n39381,n40602);
  not U42928(n39381,n39497);
  nand U42929(n39497,n40603,n40604);
  nand U42930(n40604,n40605,n35692);
  nand U42931(n40603,n39385,G59875);
  nor U42932(n40596,n40606,n39490);
  not U42933(n39490,n39385);
  nor U42934(n39385,n35691,n39371);
  not U42935(n35691,n35778);
  nand U42936(n40594,n40607,G59885);
  nand U42937(n40593,n35778,n40608);
  nand U42938(n35778,n40609,n40610);
  nand U42939(n40610,G32,n35621);
  nand U42940(n40609,G58839,n34805);
  nand U42941(n40592,n39494,n40611);
  not U42942(n39494,n39383);
  nand U42943(n39383,n40612,n40613,n39456);
  nand U42944(n40613,n34805,n21775);
  not U42945(n21775,G58863);
  nand U42946(n40612,n35621,n35622);
  not U42947(n35622,G8);
  nand U42948(G14381,n40614,n40615,n40616,n40617);
  nor U42949(n40617,n40618,n40619,n40620);
  nor U42950(n40620,n35684,n40599);
  not U42951(n35684,n39506);
  nor U42952(n39506,n40621,n40622);
  nor U42953(n40622,G15,n34805);
  nor U42954(n40621,G58856,n35621);
  nor U42955(n40619,n39395,n40602);
  not U42956(n39395,n39508);
  nand U42957(n39508,n40623,n40624);
  nand U42958(n40624,n40605,n34911);
  nand U42959(n40623,n39397,G59875);
  nor U42960(n40618,n40606,n39505);
  not U42961(n39505,n39397);
  nor U42962(n39397,n35683,n39371);
  not U42963(n35683,n35773);
  nand U42964(n40616,n40607,G59884);
  nand U42965(n40615,n35773,n40608);
  nand U42966(n35773,n40625,n40626);
  nand U42967(n40626,G31,n35621);
  nand U42968(n40625,G58840,n34805);
  nand U42969(n40614,n39507,n40611);
  not U42970(n39507,n39396);
  nand U42971(n39396,n40627,n40628,n39456);
  nand U42972(n40628,n34805,n21763);
  not U42973(n21763,G58864);
  nand U42974(n40627,n35621,n35611);
  not U42975(n35611,G7);
  nand U42976(G14380,n40629,n40630,n40631,n40632);
  nor U42977(n40632,n40633,n40634,n40635);
  nor U42978(n40635,n35676,n40599);
  not U42979(n35676,n39517);
  nor U42980(n39517,n40636,n40637);
  nor U42981(n40637,G14,n34805);
  nor U42982(n40636,G58857,n35621);
  nor U42983(n40634,n39405,n40602);
  not U42984(n39405,n39519);
  nand U42985(n39519,n40638,n40639);
  nand U42986(n40639,n40605,n35695);
  nand U42987(n40638,n39407,G59875);
  nor U42988(n40633,n40606,n39516);
  not U42989(n39516,n39407);
  nor U42990(n39407,n35675,n39371);
  not U42991(n35675,n35768);
  nand U42992(n40631,n40607,G59883);
  nand U42993(n40630,n35768,n40608);
  nand U42994(n35768,n40640,n40641);
  nand U42995(n40641,G30,n35621);
  nand U42996(n40640,G58841,n34805);
  nand U42997(n40629,n39518,n40611);
  not U42998(n39518,n39406);
  nand U42999(n39406,n40642,n40643,n39456);
  nand U43000(n40643,n34805,n21753);
  not U43001(n21753,G58865);
  nand U43002(n40642,n35621,n35602);
  not U43003(n35602,G6);
  nand U43004(G14379,n40644,n40645,n40646,n40647);
  nor U43005(n40647,n40648,n40649,n40650);
  nor U43006(n40650,n35668,n40599);
  not U43007(n35668,n39528);
  nor U43008(n39528,n40651,n40652);
  nor U43009(n40652,G13,n34805);
  nor U43010(n40651,G58858,n35621);
  nor U43011(n40649,n39415,n40602);
  not U43012(n39415,n39530);
  nand U43013(n39530,n40653,n40654);
  nand U43014(n40654,n40605,n35541);
  nand U43015(n40653,n39417,G59875);
  nor U43016(n40648,n40606,n39527);
  not U43017(n39527,n39417);
  nor U43018(n39417,n35667,n39371);
  not U43019(n35667,n35763);
  nand U43020(n40646,n40607,G59882);
  nand U43021(n40645,n35763,n40608);
  nand U43022(n35763,n40655,n40656);
  nand U43023(n40656,G29,n35621);
  nand U43024(n40655,G58842,n34805);
  nand U43025(n40644,n39529,n40611);
  not U43026(n39529,n39416);
  nand U43027(n39416,n40657,n40658,n39456);
  nand U43028(n40658,n34805,n21743);
  not U43029(n21743,G58866);
  nand U43030(n40657,n35621,n35593);
  not U43031(n35593,G5);
  nand U43032(G14378,n40659,n40660,n40661,n40662);
  nor U43033(n40662,n40663,n40664,n40665);
  nor U43034(n40665,n35659,n40599);
  not U43035(n35659,n39539);
  nor U43036(n39539,n40666,n40667);
  nor U43037(n40667,G12,n34805);
  nor U43038(n40666,G58859,n35621);
  nor U43039(n40664,n39425,n40602);
  not U43040(n39425,n39541);
  nand U43041(n39541,n40668,n40669);
  nand U43042(n40669,n40605,n39355);
  nand U43043(n40668,n39427,G59875);
  nor U43044(n40663,n40606,n39538);
  not U43045(n39538,n39427);
  nor U43046(n39427,n35658,n39371);
  not U43047(n35658,n35758);
  nand U43048(n40661,n40607,G59881);
  nand U43049(n40660,n35758,n40608);
  nand U43050(n35758,n40670,n40671);
  nand U43051(n40671,G28,n35621);
  nand U43052(n40670,G58843,n34805);
  nand U43053(n40659,n39540,n40611);
  not U43054(n39540,n39426);
  nand U43055(n39426,n40672,n40673,n39456);
  nand U43056(n40673,n34805,n21733);
  not U43057(n21733,G58867);
  nand U43058(n40672,n35621,n35584);
  not U43059(n35584,G4);
  nand U43060(G14377,n40674,n40675,n40676,n40677);
  nor U43061(n40677,n40678,n40679,n40680);
  nor U43062(n40680,n35650,n40599);
  not U43063(n35650,n39550);
  nor U43064(n39550,n40681,n40682);
  nor U43065(n40682,G11,n34805);
  nor U43066(n40681,G58860,n35621);
  nor U43067(n40679,n39435,n40602);
  not U43068(n39435,n39552);
  nand U43069(n39552,n40683,n40684);
  nand U43070(n40684,n40605,n40685);
  nand U43071(n40683,n39437,G59875);
  nor U43072(n40678,n40606,n39549);
  not U43073(n39549,n39437);
  nor U43074(n39437,n35649,n39371);
  not U43075(n35649,n35753);
  nand U43076(n40676,n40607,G59880);
  nand U43077(n40675,n35753,n40608);
  nand U43078(n35753,n40686,n40687);
  nand U43079(n40687,G27,n35621);
  nand U43080(n40686,G58844,n34805);
  nand U43081(n40674,n39551,n40611);
  not U43082(n39551,n39436);
  nand U43083(n39436,n40688,n40689,n39456);
  nand U43084(n40689,n34805,n21723);
  not U43085(n21723,G58868);
  nand U43086(n40688,n35621,n35575);
  not U43087(n35575,G3);
  nand U43088(G14376,n40690,n40691,n40692,n40693);
  nor U43089(n40693,n40694,n40695,n40696);
  nor U43090(n40696,n35641,n40599);
  not U43091(n35641,n39561);
  nor U43092(n39561,n40697,n40698);
  nor U43093(n40698,G10,n34805);
  nor U43094(n40697,G58861,n35621);
  nor U43095(n40695,n39445,n40602);
  not U43096(n39445,n39563);
  nand U43097(n39563,n40699,n40700);
  nand U43098(n40700,n40605,n35388);
  nand U43099(n40699,n39447,G59875);
  nor U43100(n40694,n40606,n39560);
  not U43101(n39560,n39447);
  nor U43102(n39447,n35640,n39371);
  not U43103(n35640,n35747);
  nand U43104(n40692,n40607,G59879);
  nand U43105(n40691,n35747,n40608);
  nand U43106(n35747,n40701,n40702);
  nand U43107(n40702,G26,n35621);
  nand U43108(n40701,G58845,n34805);
  nand U43109(n40690,n39562,n40611);
  not U43110(n40611,n37034);
  not U43111(n39562,n39446);
  nand U43112(n39446,n40703,n40704,n39456);
  nand U43113(n40704,n34805,n21711);
  not U43114(n21711,G58869);
  nand U43115(n40703,n35621,n35564);
  not U43116(n35564,G2);
  nand U43117(G14375,n40705,n40706,n40707,n40708);
  nor U43118(n40708,n40709,n40710,n40711);
  nor U43119(n40711,n39457,n40602);
  not U43120(n39457,n39591);
  nand U43121(n39591,n40712,n40713);
  nand U43122(n40713,n40605,n40714);
  nor U43123(n40605,n34901,n39371);
  nand U43124(n40712,n39468,G59875);
  nor U43125(n40710,n40606,n39577);
  not U43126(n39577,n39468);
  nor U43127(n39468,n35630,n39371);
  not U43128(n35630,n35742);
  and U43129(n40606,n40715,n40716);
  nand U43130(n40716,n40717,n36267);
  nand U43131(n40715,n40718,G59875);
  nor U43132(n40709,n37034,n39458);
  nand U43133(n39458,n40719,n40720,n39456);
  nand U43134(n40720,n34805,n26902);
  not U43135(n26902,G58870);
  or U43136(n40719,n34805,G1);
  or U43137(n40707,n40599,n35631);
  not U43138(n35631,n39588);
  nor U43139(n39588,n40721,n40722);
  nor U43140(n40722,G9,n34805);
  nor U43141(n40721,G58862,n35621);
  nand U43142(n40599,n39456,n40718);
  not U43143(n40718,n38490);
  nand U43144(n40706,n35742,n40608);
  nand U43145(n40608,n40723,n40724);
  nand U43146(n40724,n39456,n37034,n40717);
  not U43147(n40717,n40725);
  nand U43148(n40723,n40726,n40727);
  nand U43149(n35742,n40728,n40729);
  nand U43150(n40729,G25,n35621);
  nand U43151(n40728,G58846,n34805);
  nand U43152(n35621,G59809,n40730);
  nand U43153(n40730,n40731,n40732,n40733,n40734);
  nor U43154(n40734,n40735,n40736);
  or U43155(n40736,G59831,G59832,G59833,G59834);
  or U43156(n40735,G59835,G59836,G59837,G59838);
  nor U43157(n40733,n40737,G59824,G59826,G59825);
  or U43158(n40737,G59827,G59828,G59829,G59830);
  nor U43159(n40732,n40738,G59817,G59819,G59818);
  or U43160(n40738,G59820,G59821,G59822,G59823);
  nor U43161(n40731,n40739,G59810,G59812,G59811);
  or U43162(n40739,G59813,G59814,G59815,G59816);
  nand U43163(n40705,n40607,G59878);
  and U43164(n40607,n40740,n40741);
  nand U43165(n40741,n40742,n39462,n40743);
  nand U43166(n40743,G59875,n38490);
  nor U43167(n39462,n39371,n34929);
  nand U43168(n40742,n40727,n40725);
  nand U43169(n40725,n40437,n39744);
  nor U43170(n39744,G60015,n40591);
  nor U43171(n40437,n40052,n40359);
  not U43172(n40052,n39746);
  nand U43173(n40727,n39473,n40744);
  nand U43174(n40744,n37034,n38490,n39456);
  nand U43175(n37034,n40282,n39901);
  nor U43176(n39901,n40283,n40284);
  nor U43177(n40282,n40516,n40054);
  not U43178(n39473,n39576);
  nor U43179(n39576,n36215,n39371);
  nand U43180(n40740,n40726,n39467);
  nand U43181(n39467,n40746,n40747,n40748);
  or U43182(n40748,n34873,n34885);
  nand U43183(n40747,n34900,n40749);
  nand U43184(n40746,n34898,n35385,G59876);
  not U43185(n40726,n40602);
  nand U43186(n40602,n40436,n39748);
  nor U43187(n40436,n40750,n40751);
  nand U43188(G14374,n35409,n40752,n40753,n40754);
  nand U43189(n40754,n40755,G59877);
  nand U43190(n40753,n40756,n40757);
  nand U43191(n40756,n40758,n40759,n40760);
  nand U43192(n40760,n40761,n34934);
  nand U43193(n40759,n40762,n35385);
  nand U43194(n40762,G59874,n34934,n34929);
  nand U43195(n40758,n34839,n40763);
  nand U43196(n35409,G59874,G59877,n34929);
  nand U43197(G14373,n40764,n35408,n40765);
  nand U43198(n40765,G59876,n40766);
  nand U43199(n40766,n40757,n40752);
  nand U43200(n40752,G59877,n34898,n35790);
  nand U43201(n35408,n34898,n35385,n36267);
  nand U43202(n40764,n40767,n40757);
  nand U43203(n40767,n35417,n40768);
  nand U43204(n40768,n34899,n34897,n36217);
  not U43205(n35417,n34876);
  nor U43206(n34876,n35997,n35385);
  nand U43207(G14372,n35997,n39366,n40769,n40770);
  or U43208(n40770,n40745,G59877);
  nand U43209(n40769,n34899,n34898,G59876,G59877);
  nand U43210(G14371,n40771,n34873,n40772);
  nand U43211(n40772,n40755,G59874);
  not U43212(n40755,n40757);
  nand U43213(n40757,n40773,n40774,n40775);
  nand U43214(n40775,n40776,n35385);
  nand U43215(n40776,n35790,G59876);
  nand U43216(n40774,n35996,n34914,n35392);
  nor U43217(n35392,G60246,n35790);
  nand U43218(n40773,n40777,n39366);
  or U43219(n40777,n40763,n35997);
  not U43220(n35997,n34839);
  nor U43221(n34839,n34898,G59876);
  nand U43222(n40763,n40778,n40779,n40780,n40781);
  nor U43223(n40781,n40782,n40783,n40784,n40785);
  and U43224(n40785,n34840,n34841);
  xnor U43225(n34840,n40786,n38689);
  and U43226(n38689,n40787,n40788);
  nand U43227(n40787,n40789,n40790);
  nand U43228(n40786,n38690,n38687);
  nand U43229(n38687,n40791,n40792);
  or U43230(n38690,n40792,n40791);
  nor U43231(n40791,n34968,n37262);
  xor U43232(n40792,n40793,n36267);
  nand U43233(n40793,n40794,n40795,n40796,n40797);
  nor U43234(n40797,n40798,n40799);
  nor U43235(n40799,n36214,n36186);
  nor U43236(n40798,n35998,n38703);
  not U43237(n38703,G60211);
  nand U43238(n40796,G60020,n36328);
  nand U43239(n40795,G60006,n40800);
  nand U43240(n40800,n35789,n40801);
  nand U43241(n40801,n35894,G59877);
  nand U43242(n40794,n35528,n36329);
  not U43243(n35528,n35338);
  xnor U43244(n35338,n38683,n38682);
  xnor U43245(n38683,n34962,n40802);
  nor U43246(n40802,n40803,n40804,n40805,n40806);
  and U43247(n40806,n36269,G60147);
  nor U43248(n40805,n36527,n38553);
  not U43249(n38553,G60020);
  nor U43250(n40804,n36215,n36186);
  not U43251(n36186,G60052);
  nor U43252(n40803,n38073,n35339);
  not U43253(n35339,G60179);
  not U43254(n38073,n36266);
  nor U43255(n40784,n38713,n34877);
  nor U43256(n40783,n39345,n39325);
  nor U43257(n40782,n40807,n40808);
  nor U43258(n40780,n36218,n40809);
  nor U43259(n40809,n40810,n34955);
  nand U43260(n34955,n34945,n40811);
  nand U43261(n40811,n40812,n34899);
  nand U43262(n40812,n40813,n34913,n40814);
  nand U43263(n40814,n35994,n35695);
  and U43264(n34945,n40815,n40816,n40817,n40818);
  nand U43265(n40817,n38712,n40819);
  nand U43266(n40819,n40820,n40821);
  nor U43267(n40815,n40822,n40823);
  nor U43268(n40823,n39350,n34934);
  nor U43269(n40822,n39345,n40813);
  not U43270(n39345,n34959);
  nor U43271(n40810,G60244,G60245);
  nand U43272(n40779,n40824,n39369);
  nand U43273(n40824,n40825,n40826);
  nand U43274(n40826,n40827,n40750,n40828);
  not U43275(n40828,n40808);
  nand U43276(n40825,n40829,n40751);
  nand U43277(n40829,n40808,n40830);
  nand U43278(n40830,n40831,n40827);
  nand U43279(n40827,n40832,n40833,n40834,n40835);
  nand U43280(n40835,n40836,n40837);
  nand U43281(n40837,n40838,n40839);
  nand U43282(n40839,G60009,n40840);
  nand U43283(n40834,n40841,n34867,n34877);
  nand U43284(n34867,n40842,n40843,n40844,n40845);
  nor U43285(n40845,n40846,n40847,n40848);
  nor U43286(n40848,n40849,n40054);
  nor U43287(n40847,n40850,n40851);
  nor U43288(n40850,n38200,n36989);
  not U43289(n36989,n36986);
  nor U43290(n36986,n40852,n38193);
  nor U43291(n40852,n38219,n34912);
  nor U43292(n40846,n39228,n39324);
  nor U43293(n39228,n38193,n38200);
  nand U43294(n40844,n35375,n40853);
  nand U43295(n40843,n34869,n40854);
  not U43296(n34869,n35374);
  xnor U43297(n35374,n40855,n40856);
  and U43298(n40856,n40857,n40858);
  nand U43299(n40842,n34868,n40859);
  or U43300(n40841,n34881,n40840);
  not U43301(n40840,n39748);
  nand U43302(n40833,n40860,n40861);
  nand U43303(n40860,n40862,n40863,G60015);
  nand U43304(n40863,n40836,G60010);
  nand U43305(n40862,n34881,n34877);
  nand U43306(n34881,n40864,n40865,n40866,n40867);
  nor U43307(n40867,n40868,n40869);
  nor U43308(n40869,n40870,n39314);
  not U43309(n39314,n34938);
  nor U43310(n40868,n40871,n34883);
  nand U43311(n40866,n34884,n40854);
  xor U43312(n34884,n40872,n36215);
  nand U43313(n40872,n40873,n40874);
  nand U43314(n40865,n40875,n36985);
  nand U43315(n40864,n40361,n40876);
  or U43316(n40832,n40807,G60013);
  nand U43317(n40831,G60013,n40807);
  nand U43318(n40807,n40877,n40878);
  nand U43319(n40878,n40836,n40879);
  or U43320(n40877,n34858,n40836);
  nand U43321(n34858,n40880,n40881,n40882,n40883);
  nor U43322(n40883,n40884,n40885,n40886);
  nor U43323(n40886,n39324,n39236);
  xor U43324(n39236,n40887,n40838);
  not U43325(n40838,n38192);
  nor U43326(n40885,n40849,n40283);
  nor U43327(n40884,n40871,n40888);
  nand U43328(n40882,n36958,n39187);
  xor U43329(n36958,G60008,n40889);
  nand U43330(n40881,n35364,n40853);
  nand U43331(n40880,n34860,n40854);
  not U43332(n34860,n35362);
  nand U43333(n35362,n40890,n40891);
  nand U43334(n40891,n40892,n40893);
  not U43335(n40892,n40894);
  nand U43336(n40890,n40895,n40858,n40896);
  nand U43337(n40895,n40897,n40893);
  nand U43338(n40808,n40898,n40899);
  nand U43339(n40899,n40836,n38831);
  or U43340(n40898,n34851,n40836);
  not U43341(n40836,n34877);
  nand U43342(n34877,n40900,n40901,n39341);
  and U43343(n39341,n40902,n40903,n40904,n40905);
  nor U43344(n40905,n40906,n40907);
  xnor U43345(n40907,n40821,n40908);
  not U43346(n40906,n40816);
  nor U43347(n40816,n40909,n40910,n39201,n40911);
  and U43348(n40909,n40912,n35695);
  nand U43349(n40912,n40913,n35388,n34912);
  not U43350(n40903,n40914);
  nand U43351(n40902,n35779,n40915);
  nand U43352(n40915,n35994,n39355);
  nand U43353(n40901,n40916,n34899);
  nand U43354(n40916,n40917,n40918);
  nand U43355(n40918,n40919,n34934);
  nand U43356(n40919,n39330,n40920);
  nand U43357(n40920,n34914,n40921);
  nand U43358(n40921,n35416,n39329);
  not U43359(n39329,n35894);
  not U43360(n34914,n34913);
  nand U43361(n34913,n35895,n39198);
  or U43362(n40917,n39325,n34959);
  nand U43363(n34959,n40922,n40923);
  nand U43364(n40923,n40924,n40925,n40926,n40927);
  nand U43365(n40927,n40928,n40929,n40930);
  or U43366(n40930,n40931,n34911);
  nand U43367(n40929,n40932,n40933,n40934);
  not U43368(n40934,n40935);
  not U43369(n40933,n39070);
  nand U43370(n40932,n40936,n40937);
  or U43371(n40928,n40937,n40936);
  nand U43372(n40926,n40931,n34911);
  not U43373(n40924,n40938);
  nand U43374(n40900,n40875,n34934);
  nand U43375(n34851,n40939,n40940,n40941,n40942);
  nor U43376(n40942,n40943,n40944,n40945);
  nor U43377(n40945,n39324,n39227);
  nand U43378(n39227,n40946,n40947,n40948);
  nand U43379(n40948,n40949,n35692);
  or U43380(n40947,n40950,n38831);
  nand U43381(n40946,n40951,n40950);
  nand U43382(n40950,n40887,n38192);
  xnor U43383(n40887,n34912,G60008);
  nand U43384(n40951,n40952,n40953);
  nand U43385(n40953,n34912,n38831);
  nor U43386(n40944,n40870,n36193);
  not U43387(n36193,n35352);
  not U43388(n40870,n40853);
  nand U43389(n40853,n40954,n39334,n40955,n39332);
  nand U43390(n39332,n40956,n39355);
  nor U43391(n40955,n39338,n40957);
  nor U43392(n40957,n35994,n40958);
  nor U43393(n39338,n35781,n39355);
  not U43394(n35781,n36305);
  not U43395(n40954,n39336);
  nand U43396(n39336,n35416,n40959,n40960,n40961);
  nand U43397(n40961,n39070,n34912);
  nand U43398(n40960,n40962,n35692);
  nand U43399(n40962,n40963,n40964);
  nand U43400(n40964,n35542,n40965);
  nand U43401(n40965,n40911,n40966);
  nand U43402(n40966,n40813,n34911);
  nand U43403(n40963,n39201,n40813);
  not U43404(n40813,n39350);
  nor U43405(n39350,n35695,n35994);
  nand U43406(n40959,n39201,n40967);
  nand U43407(n40967,n39320,n40908);
  nor U43408(n40943,n40871,n40968);
  not U43409(n40871,n40859);
  nand U43410(n40859,n40969,n39325);
  nand U43411(n40941,n34850,n40854);
  nand U43412(n40854,n39327,n39328,n39323,n39330);
  not U43413(n39330,n34841);
  not U43414(n39328,n40970);
  xnor U43415(n34850,n40789,n40971);
  and U43416(n40971,n40790,n40788);
  nand U43417(n40788,n40972,n40973,n40974);
  nand U43418(n40974,n35545,G60002);
  nand U43419(n40790,G60002,n40975,n35545);
  nand U43420(n40975,n40972,n40973);
  or U43421(n40973,n40976,n36215);
  nand U43422(n40972,n40976,n36215);
  nand U43423(n40976,n40977,n40978,n40979,n40980);
  nor U43424(n40980,n40981,n40982);
  nor U43425(n40982,n36214,n35348);
  nor U43426(n40981,n35998,n35351);
  not U43427(n35351,G60210);
  nand U43428(n40979,G60007,n40983);
  nand U43429(n40978,n35352,n36329);
  nor U43430(n35352,n40984,n38682);
  nor U43431(n38682,n40985,n40986);
  and U43432(n40984,n40986,n40985);
  xor U43433(n40986,n40987,n35998);
  nand U43434(n40987,n40988,n40989,n40990,n40991);
  nor U43435(n40991,n40992,n40993,n40994,n40995);
  nor U43436(n40995,n36215,n35348);
  not U43437(n35348,G60051);
  and U43438(n40994,n36266,G60178);
  nor U43439(n40993,n40996,n38831);
  nor U43440(n40992,n40516,n40745);
  not U43441(n40516,n39903);
  nor U43442(n40990,n40997,n40998);
  and U43443(n40998,n36269,G60146);
  nor U43444(n40997,n36527,n38702);
  not U43445(n38702,G60019);
  nand U43446(n40989,n34929,G60012);
  nand U43447(n40988,n39368,n34900);
  nand U43448(n40977,G60019,n36328);
  and U43449(n40789,n40893,n40894);
  nand U43450(n40894,n40897,n40999);
  nand U43451(n40999,n40896,n40858);
  nand U43452(n40858,n41000,n41001);
  nand U43453(n41001,n41002,n41003);
  nand U43454(n40896,n40855,n40857);
  nand U43455(n40857,n41002,n41003,n41004);
  not U43456(n41004,n41000);
  nand U43457(n41000,n35998,n39366,n41005,n41006);
  nor U43458(n41006,n41007,n41008,n41009);
  nor U43459(n41009,n35994,n41010);
  nor U43460(n41008,n36898,n34968);
  nand U43461(n41005,n39069,n41011,n40820,G59877);
  and U43462(n39069,n39198,n35692,n40821);
  or U43463(n41003,n41012,n36215);
  nand U43464(n41002,n36215,n41012);
  nand U43465(n41012,n41013,n41014,n41015,n41016);
  nor U43466(n41016,n41017,n41018);
  nor U43467(n41018,n36214,n35373);
  nor U43468(n41017,n35998,n34984);
  not U43469(n34984,G60208);
  nand U43470(n41015,n35375,n36329);
  not U43471(n35375,n36207);
  xor U43472(n36207,n41019,n41020);
  nand U43473(n41019,n41021,n41022);
  nand U43474(n41014,G60017,n36328);
  nand U43475(n41013,G60009,n40983);
  nand U43476(n40855,n40874,n41023);
  nand U43477(n41023,n36267,n40873);
  nand U43478(n40873,n41024,n41025,n41026);
  not U43479(n41026,n41027);
  nand U43480(n40874,n41027,n41028);
  nand U43481(n41028,n41024,n41025);
  or U43482(n41025,n41029,n36215);
  nand U43483(n41024,n41029,n36215);
  nand U43484(n41029,n41030,n41031,n41032,n41033);
  nor U43485(n41033,n41034,n41035);
  nor U43486(n41035,n36214,n35384);
  nor U43487(n41034,n35998,n34982);
  not U43488(n34982,G60207);
  nand U43489(n41032,G60010,n40983);
  nand U43490(n41031,n34938,n36329);
  nand U43491(n34938,n41036,n41037);
  nand U43492(n41037,n41038,n41039);
  nand U43493(n41038,n41040,n41041);
  nand U43494(n41041,n41042,n35998);
  or U43495(n41036,n41039,n35998);
  nand U43496(n41030,G60016,n36328);
  nand U43497(n41027,n41043,n41044,n41045,n34901);
  nand U43498(n41044,G59877,n41046);
  nand U43499(n41046,n41047,n40714,n41048,n41049);
  nor U43500(n41049,n41050,n41051,n41052,n41053);
  nor U43501(n41051,n41054,n41055);
  nor U43502(n41055,n41056,n41057);
  nor U43503(n41057,n35542,n40685);
  nor U43504(n41056,n35994,n34934);
  nor U43505(n41050,n35541,n35388);
  nand U43506(n41048,n35779,n40913);
  not U43507(n41047,n40956);
  nand U43508(n41043,n35545,G60005);
  nand U43509(n40897,n41058,n41059,n41045,n40745);
  xnor U43510(n41058,n36267,n41060);
  nand U43511(n40893,n41061,n41062);
  nand U43512(n41062,n41045,n40745,n41059);
  nand U43513(n41059,n35545,G60003);
  xnor U43514(n41061,n41060,n36215);
  nand U43515(n41060,n41063,n41064,n41065,n41066);
  nand U43516(n41066,G60008,n40983);
  nand U43517(n40983,n35789,n35785,n34901,n41067);
  nor U43518(n41067,n41068,n41069,n41070);
  nor U43519(n41070,n35994,n35385,n39322,n34934);
  not U43520(n39322,n36218);
  nor U43521(n41069,n41071,n35385);
  nor U43522(n41071,n35894,n40970);
  nor U43523(n40970,n41072,n35692);
  nor U43524(n41068,n35385,n39327);
  not U43525(n35785,n36269);
  nor U43526(n41065,n41073,n41074);
  nor U43527(n41074,n36278,n38815);
  not U43528(n36278,n36328);
  and U43529(n41076,n41077,n41078,n41045);
  nand U43530(n41045,G59877,n35388,n39349,n41079);
  and U43531(n41079,n41011,n38363);
  nor U43532(n38363,n34923,n34912);
  nand U43533(n41075,G59877,n39337);
  nand U43534(n39337,n40969,n41080);
  and U43535(n40969,n41081,n41082);
  nand U43536(n41082,n40956,n41083,n40911);
  or U43537(n41081,n41072,n34912);
  and U43538(n41073,n36329,n35364);
  not U43539(n35364,n36200);
  nand U43540(n36200,n41084,n40985);
  nand U43541(n40985,n41085,n41086);
  nand U43542(n41086,n41087,n41021);
  xnor U43543(n41085,n41088,n35998);
  nand U43544(n41084,n41087,n41021,n41089);
  xnor U43545(n41089,n34962,n41088);
  nand U43546(n41088,n41090,n41091,n41092,n41093);
  nor U43547(n41093,n41094,n41095,n41096,n41097);
  nor U43548(n41097,n40888,n39366);
  nor U43549(n41096,n40745,n40283);
  nand U43550(n40283,n41098,n41099);
  nand U43551(n41099,n41100,n41101);
  nand U43552(n41100,n41102,n41103);
  nand U43553(n41098,n41104,n34915);
  xor U43554(n41104,n41105,n41106);
  nor U43555(n41095,n40750,n34901);
  and U43556(n41094,n36269,G60145);
  nor U43557(n41092,n41107,n41108);
  nor U43558(n41108,n36527,n38815);
  not U43559(n38815,G60018);
  nor U43560(n41107,n36215,n35361);
  not U43561(n35361,G60050);
  nand U43562(n41091,G60008,n41109);
  nand U43563(n41090,G60177,n36266);
  nand U43564(n41021,n41110,n41111);
  nand U43565(n41111,n41078,n36215,n34967,n41112);
  and U43566(n41112,n41113,n41114);
  xnor U43567(n41110,n41115,n35998);
  nand U43568(n41087,n41022,n41020);
  nand U43569(n41020,n41039,n41116);
  nand U43570(n41116,n34962,n41040);
  nand U43571(n41040,n41117,n41118);
  not U43572(n41117,n41042);
  nand U43573(n41039,n41119,n41042);
  nand U43574(n41042,n36214,n41120,n34967,n34901);
  nand U43575(n41120,G59877,n41121);
  nand U43576(n41121,n41122,n41123,n41124,n41125);
  nor U43577(n41125,n41126,n41127,n41128);
  nor U43578(n41128,n35542,n41129);
  nor U43579(n41127,n39349,n41130,n41131);
  nor U43580(n41131,n35542,n40821);
  nor U43581(n41130,n41054,n40685);
  nor U43582(n41126,n35695,n39320);
  not U43583(n41124,n41052);
  nand U43584(n41052,n41132,n41133,n41134,n41135);
  nor U43585(n41135,n40914,n40910);
  nand U43586(n41134,n40821,n35695);
  nand U43587(n41133,n35542,n35692);
  nand U43588(n41132,n40820,n34912);
  nand U43589(n41123,n35779,n34911);
  nand U43590(n41122,n40911,n35994);
  not U43591(n36214,n37121);
  xnor U43592(n41119,n41118,n35998);
  nand U43593(n41118,n41136,n41137);
  nor U43594(n41137,n41138,n41139,n41140,n41141);
  nor U43595(n41141,n40745,n40284);
  not U43596(n40284,n40361);
  nor U43597(n40361,n41142,n41143);
  nor U43598(n41143,n34927,n41144);
  and U43599(n41144,G60010,n41145);
  nor U43600(n41140,n36215,n35384);
  not U43601(n35384,G60048);
  and U43602(n41139,n36266,G60175);
  nor U43603(n41138,n40996,n36985);
  nor U43604(n41136,n41146,n41147,n41148,n41149);
  nor U43605(n41149,n39366,n34883);
  nor U43606(n41148,n40439,n34901);
  and U43607(n41147,n36269,G60143);
  nor U43608(n41146,n36527,n39057);
  nand U43609(n41022,n41150,n41113,n41114,n41151);
  not U43610(n35896,n41078);
  not U43611(n41114,n41007);
  nand U43612(n41007,n35789,n41152);
  nand U43613(n41152,G59877,n35388,n41153);
  nand U43614(n41113,n40956,n41083,G59877,n39198);
  xnor U43615(n41150,n34962,n41115);
  nand U43616(n41115,n41154,n41155);
  nor U43617(n41155,n41156,n41157,n41158,n41159);
  nor U43618(n41159,n36215,n35373);
  not U43619(n35373,G60049);
  and U43620(n41158,n36266,G60176);
  nand U43621(n36266,n35998,n41160);
  nand U43622(n41160,n35546,G59877);
  nor U43623(n41157,n40996,n38219);
  not U43624(n40996,n41109);
  nand U43625(n41109,n34967,n41077,n41078,n41010);
  nand U43626(n41010,G59877,n34934,n36218);
  nand U43627(n41078,G59877,n39198,n35996);
  not U43628(n35996,n35416);
  nand U43629(n41077,G59877,n41161);
  nand U43630(n41161,n41162,n41163,n39334,n41164);
  nor U43631(n41164,n41165,n41166,n41167);
  nor U43632(n41167,n34912,n41168);
  nor U43633(n41168,n41169,n41170,n41171);
  nor U43634(n41171,n40685,n40911,n41054);
  nor U43635(n41170,n40821,n35541);
  nor U43636(n41169,n34911,n35780);
  nor U43637(n41166,n41172,n40818);
  not U43638(n40818,n35779);
  nor U43639(n35779,n35692,n35695);
  nor U43640(n41172,n41173,n40820);
  nor U43641(n41173,n41054,n34923);
  nor U43642(n41165,n41174,n41175);
  and U43643(n39334,n41176,n41177,n41178,n41179);
  nor U43644(n41179,n40910,n41180,n40914);
  nor U43645(n40914,n34911,n38981);
  not U43646(n38981,n39200);
  and U43647(n41180,n35695,n41129);
  nor U43648(n40910,n35542,n38712);
  not U43649(n41178,n41053);
  nand U43650(n41053,n41181,n41182);
  nand U43651(n41182,n41183,n40685);
  nand U43652(n41183,n40908,n40904);
  nand U43653(n40904,n39355,n35388);
  not U43654(n40908,n40820);
  nand U43655(n41181,n39355,n35541,n40821);
  nand U43656(n41177,n35780,n35388,n40821);
  nand U43657(n41176,n41184,n41185);
  nand U43658(n41185,n39349,n35542,n41186,n34923);
  nand U43659(n41184,n41187,n40714);
  nand U43660(n41187,n41153,n39349);
  not U43661(n41153,n41186);
  nand U43662(n41163,n41188,n36305);
  nand U43663(n41162,n40956,n39201);
  not U43664(n34967,n36390);
  nor U43665(n36390,n40851,n35385);
  nor U43666(n41156,n40054,n40745);
  not U43667(n40054,n39902);
  xor U43668(n39902,n41189,n41190);
  xnor U43669(n41189,n41142,n41191);
  nor U43670(n41154,n41192,n41193,n41194,n41195);
  nor U43671(n41195,n41196,n39366);
  nor U43672(n41194,n40861,n34901);
  not U43673(n34901,n34929);
  nor U43674(n34929,G59876,G59875);
  and U43675(n41193,n36269,G60144);
  nor U43676(n36269,n39323,n35385);
  nand U43677(n39323,n39199,n34912,n41197);
  nor U43678(n41192,n36527,n39059);
  not U43679(n36527,n36268);
  nand U43680(n36268,n35789,n41198);
  nand U43681(n41198,G59877,n41199);
  nand U43682(n41199,n41200,n41201,n39327,n41072);
  nand U43683(n41072,n35402,n40821,n40911,n41202);
  nor U43684(n41202,n39355,n38712,n35541);
  nand U43685(n39327,n39355,n41203);
  nand U43686(n41203,n41204,n41186);
  nand U43687(n41186,n39199,n41205);
  nor U43688(n39199,n40685,n34911);
  nand U43689(n41204,n41205,n35402);
  nor U43690(n41205,n35692,n40911,n35780);
  nand U43691(n41201,n41083,n39198,n40956);
  nand U43692(n41200,n34885,n36218);
  nor U43693(n36218,n40958,n41206);
  not U43694(n40958,n41188);
  nor U43695(n41188,n39320,n35695,n41054,n40911);
  nand U43696(n35789,n34841,G59877);
  nor U43697(n34841,n35415,n34911);
  nand U43698(n36329,n36215,n34968);
  not U43699(n34968,n35545);
  nand U43700(n41064,G60209,n34962);
  nand U43701(n39325,n41011,n39070,n40820,n35692);
  nor U43702(n40820,n35388,n39355);
  nand U43703(n41063,G60050,n37121);
  nand U43704(n37121,n39366,n40745);
  nand U43705(n40745,G60246,G59876);
  not U43706(n39366,n34900);
  nand U43707(n40940,n39903,n40876);
  not U43708(n40876,n40849);
  nor U43709(n40849,n35894,n35546);
  not U43710(n35546,n41080);
  nand U43711(n41080,n39070,n35692,n41197);
  nor U43712(n41197,n40714,n35780,n39355,n41054);
  not U43713(n35780,n39201);
  nor U43714(n39201,n35541,n35695);
  nor U43715(n35894,n35415,n35994);
  nand U43716(n39903,n41207,n41208);
  nand U43717(n41208,n41209,n41210);
  nand U43718(n41209,n41102,n41211);
  nand U43719(n41211,n41103,n41101);
  nand U43720(n41207,n41212,n41213);
  nand U43721(n41213,n41103,n41214);
  nand U43722(n41214,n34915,n41102);
  or U43723(n41102,n41106,n41105);
  nand U43724(n41103,n41105,n41106);
  nand U43725(n41106,n41215,n41216);
  nand U43726(n41216,G60008,n41145);
  nand U43727(n41215,n34859,n34898);
  nand U43728(n41105,n41217,n41218);
  nand U43729(n41218,n41219,n41220);
  or U43730(n41220,n41190,n41142);
  not U43731(n41219,n41191);
  nand U43732(n41217,n41190,n41142);
  nand U43733(n41142,n41221,n41222);
  nand U43734(n41222,n34927,n41145,G60010);
  nand U43735(n34927,n34912,G59875);
  nand U43736(n41221,n34940,n34898);
  nand U43737(n41190,n41223,n41224);
  nand U43738(n41224,G60009,n41145);
  nand U43739(n41223,n34868,n34898);
  not U43740(n41212,n41210);
  nand U43741(n41210,n41225,n41226);
  nand U43742(n41226,G60007,n41145);
  nand U43743(n41145,n41191,n41101,n41227);
  nand U43744(n41227,G59875,n35692);
  not U43745(n41101,n34915);
  nor U43746(n34915,n34911,n34898);
  nand U43747(n41191,G59875,n41228);
  nand U43748(n41228,n41206,n41229);
  nand U43749(n41229,n40956,n39198);
  nand U43750(n39198,n41230,n41231);
  nand U43751(n41231,G59839,n34951);
  nor U43752(n40956,n35692,n35994);
  not U43753(n41206,n41174);
  nor U43754(n41174,n35542,n34912);
  nand U43755(n41225,n39368,n34898);
  nand U43756(n40939,n39187,n36959);
  nand U43757(n36959,n41232,n41233);
  nand U43758(n41233,n40952,n40879,n40889);
  not U43759(n40952,n41234);
  nand U43760(n41232,n41235,n38831);
  nand U43761(n41235,n41234,n40889);
  nand U43762(n40889,n34912,n38192);
  not U43763(n39187,n40851);
  nand U43764(n40778,n34885,n41236);
  nand U43765(n41236,n35416,n35415,n41237);
  not U43766(n41237,n40875);
  nand U43767(n40875,n39324,n40851);
  nand U43768(n40851,n36305,n41129,n41238);
  nor U43769(n41238,n34923,n39349,n35695);
  not U43770(n34923,n40936);
  nor U43771(n41129,n35388,n40911);
  nand U43772(n39324,n35393,n41011,n39200,n40685);
  nand U43773(n35415,n34912,n40714,n41083);
  nor U43774(n41083,n39320,n35541,n38712,n41054);
  not U43775(n39320,n40913);
  nor U43776(n40913,n39355,n40821);
  nand U43777(n35416,n39349,n35692,n40821,n41239);
  and U43778(n41239,n41011,n35402);
  nor U43779(n35402,n35388,n34911);
  nor U43780(n41011,n35542,n40911,n35695);
  not U43781(n40911,n40714);
  nand U43782(n40714,n41240,n41241,n41242,n41243);
  nor U43783(n41243,n41244,n41245,n41246,n41247);
  nor U43784(n41247,n41248,n37004);
  nor U43785(n41246,n41249,n37002);
  nor U43786(n41245,n41250,n37020);
  nor U43787(n41244,n41251,n37016);
  nor U43788(n41242,n41252,n41253,n41254,n41255);
  nor U43789(n41255,n41256,n37014);
  nor U43790(n41254,n41257,n36388);
  nor U43791(n41253,n41258,n36384);
  nor U43792(n41252,n41259,n36382);
  nor U43793(n41241,n41260,n41261,n41262,n41263);
  nor U43794(n41263,n41264,n36376);
  nor U43795(n41262,n41265,n36372);
  nor U43796(n41261,n41266,n36370);
  nor U43797(n41260,n41267,n37008);
  nor U43798(n41240,n41268,n41269,n41270,n41271);
  nor U43799(n41271,n41272,n37006);
  nor U43800(n41270,n41273,n37018);
  nor U43801(n41269,n41274,n36386);
  nor U43802(n41268,n41275,n36374);
  not U43803(n39349,n39355);
  nand U43804(n39355,n41276,n41277,n41278,n41279);
  nor U43805(n41279,n41280,n41281,n41282,n41283);
  nor U43806(n41283,n41248,n37260);
  not U43807(n37260,G59985);
  nor U43808(n41282,n41249,n37259);
  not U43809(n37259,G59977);
  nor U43810(n41281,n41250,n37270);
  not U43811(n37270,G59969);
  nor U43812(n41280,n41251,n37268);
  not U43813(n37268,G59953);
  nor U43814(n41278,n41284,n41285,n41286,n41287);
  nor U43815(n41287,n41256,n37267);
  not U43816(n37267,G59945);
  nor U43817(n41286,n41257,n36641);
  not U43818(n36641,G59937);
  nor U43819(n41285,n41258,n36639);
  not U43820(n36639,G59921);
  nor U43821(n41284,n41259,n36638);
  not U43822(n36638,G59913);
  nor U43823(n41277,n41288,n41289,n41290,n41291);
  nor U43824(n41291,n41264,n36633);
  not U43825(n36633,G59905);
  nor U43826(n41290,n41265,n36631);
  not U43827(n36631,G59889);
  nor U43828(n41289,n41266,n36630);
  not U43829(n36630,G59881);
  nor U43830(n41288,n41267,n37262);
  not U43831(n37262,G60001);
  nor U43832(n41276,n41292,n41293,n41294,n41295);
  nor U43833(n41295,n41272,n37261);
  not U43834(n37261,G59993);
  nor U43835(n41294,n41273,n37269);
  not U43836(n37269,G59961);
  nor U43837(n41293,n41274,n36640);
  not U43838(n36640,G59929);
  nor U43839(n41292,n41275,n36632);
  not U43840(n36632,G59897);
  not U43841(n34885,n34934);
  nand U43842(n34934,n41296,n41297);
  or U43843(n41297,n41298,n41299);
  nand U43844(n41296,n41300,n41298,n41301,n41302);
  nor U43845(n41302,n41303,n41304);
  nor U43846(n41304,n41305,n40922);
  nand U43847(n40922,n41306,n41307);
  nand U43848(n41307,G60011,n41308);
  nand U43849(n41308,G60006,n41309);
  or U43850(n41306,n41309,G60006);
  nor U43851(n41303,n38713,G60244,n40749);
  not U43852(n38713,G60006);
  nand U43853(n41301,n41310,n41311,n41312,n41313);
  nor U43854(n41313,n41314,n41315);
  nor U43855(n41315,n41305,n40925);
  xnor U43856(n40925,n41309,n41316);
  xnor U43857(n41316,n39369,G60006);
  not U43858(n39369,G60011);
  nand U43859(n41309,n41317,n41318);
  nand U43860(n41318,n41319,n40751);
  nand U43861(n41319,n41320,n38831);
  nand U43862(n41317,G60007,n41321);
  nor U43863(n41314,G60007,n41322);
  nand U43864(n41312,n41323,n40938);
  nand U43865(n40938,n41324,n41325);
  nand U43866(n41325,n41326,n41321);
  xnor U43867(n41326,G60012,G60007);
  nand U43868(n41324,n41327,n41320);
  not U43869(n41320,n41321);
  nand U43870(n41321,n41328,n41329);
  nand U43871(n41329,n41330,n40750);
  nand U43872(n41330,n40879,n41331);
  or U43873(n41328,n41331,n40879);
  xnor U43874(n41327,n40751,G60007);
  nand U43875(n41311,n41332,n41333);
  nand U43876(n41333,n41334,n41335);
  nand U43877(n41335,n41336,n41337);
  nand U43878(n41337,n34897,n41338,G60008);
  nand U43879(n41332,n41322,n41339);
  nand U43880(n41310,n41340,n41341,n41342);
  nand U43881(n41342,n41343,n41344);
  nand U43882(n41344,n41322,n41345);
  not U43883(n41343,n41346);
  nand U43884(n41341,n41339,n41334,n41322);
  nand U43885(n41334,n41323,n40931);
  xor U43886(n40931,n41347,n41331);
  nand U43887(n41331,n41348,n41349);
  nand U43888(n41349,G60014,n41350);
  or U43889(n41350,n41351,n38219);
  nand U43890(n41348,n41351,n38219);
  xnor U43891(n41347,G60013,G60008);
  nand U43892(n41340,n41352,n41353,n41354);
  nand U43893(n41354,n41336,n36985);
  nand U43894(n41353,n41355,n40749);
  nand U43895(n41355,n41356,n41339);
  nand U43896(n41339,n41175,n41357);
  nand U43897(n41357,n41054,n40685);
  nand U43898(n41356,n41345,n41346);
  nand U43899(n41346,n41358,n41359,n41360);
  nand U43900(n41360,n41323,n40937);
  xnor U43901(n40937,n41351,n41361);
  xnor U43902(n41361,n40861,G60009);
  not U43903(n41359,n41362);
  nand U43904(n41358,n41363,n41336);
  nand U43905(n41363,n41364,n41365,n34897);
  not U43906(n34897,G59874);
  nand U43907(n41365,n38219,n41338);
  not U43908(n41338,G60244);
  nand U43909(n41364,G60244,n41366);
  nand U43910(n41366,G60016,n34868);
  nand U43911(n41345,n41367,n41368);
  nand U43912(n41368,n40936,n41054);
  nor U43913(n40936,n34911,n40821);
  not U43914(n41367,n41299);
  nand U43915(n41352,n41323,n40935);
  nand U43916(n40935,n41351,n41369);
  nand U43917(n41369,G60015,n36985);
  nand U43918(n41351,G60010,n40439);
  not U43919(n41323,n41305);
  nand U43920(n41305,n41322,n41370);
  nand U43921(n41370,n41299,n41175);
  not U43922(n41175,n35393);
  nor U43923(n35393,n35388,n35994);
  nor U43924(n41299,n35542,n35994,n40821);
  not U43925(n40821,n40685);
  nand U43926(n41298,n41362,n38364);
  nand U43927(n38364,n41371,n41372,n41373,n41374);
  nor U43928(n41374,n41375,n41376,n41377,n41378);
  nor U43929(n41378,n37004,n38472);
  nand U43930(n38472,n41379,n41380);
  not U43931(n37004,G59982);
  nor U43932(n41377,n37002,n38473);
  nand U43933(n38473,n41379,n41381);
  not U43934(n37002,G59974);
  nor U43935(n41376,n37020,n38474);
  nand U43936(n38474,n41382,n41383);
  not U43937(n37020,G59966);
  nor U43938(n41375,n37016,n38475);
  nand U43939(n38475,n41383,n41380);
  not U43940(n37016,G59950);
  nor U43941(n41373,n41384,n41385,n41386,n41387);
  nor U43942(n41387,n37014,n38480);
  nand U43943(n38480,n41381,n41383);
  not U43944(n37014,G59942);
  nor U43945(n41386,n36388,n38481);
  nand U43946(n38481,n41388,n41382);
  not U43947(n36388,G59934);
  nor U43948(n41385,n36384,n38482);
  nand U43949(n38482,n41388,n41380);
  not U43950(n36384,G59918);
  nor U43951(n41384,n36382,n38483);
  nand U43952(n38483,n41388,n41381);
  not U43953(n36382,G59910);
  nor U43954(n41372,n41389,n41390,n41391,n41392);
  nor U43955(n41392,n36376,n38488);
  nand U43956(n38488,n41393,n41382);
  not U43957(n36376,G59902);
  nor U43958(n41391,n36372,n38489);
  nand U43959(n38489,n41393,n41380);
  nor U43960(n41380,n41196,n34940);
  not U43961(n36372,G59886);
  nor U43962(n41390,n36370,n38490);
  nand U43963(n38490,n41393,n41381);
  nor U43964(n41381,n34883,n41196);
  not U43965(n41196,n34868);
  not U43966(n36370,G59878);
  nor U43967(n41389,n37008,n38491);
  nand U43968(n38491,n41379,n41382);
  nor U43969(n41382,n34868,n34940);
  not U43970(n34940,n34883);
  not U43971(n37008,G59998);
  nor U43972(n41371,n41394,n41395,n41396,n41397);
  nor U43973(n41397,n37006,n38496);
  nand U43974(n38496,n41398,n41379);
  nor U43975(n41379,n34859,n39368);
  not U43976(n37006,G59990);
  nor U43977(n41396,n37018,n38497);
  nand U43978(n38497,n41398,n41383);
  nor U43979(n41383,n40888,n39368);
  not U43980(n39368,n40968);
  not U43981(n37018,G59958);
  nor U43982(n41395,n36386,n38498);
  nand U43983(n38498,n41398,n41388);
  nor U43984(n41388,n40968,n34859);
  not U43985(n36386,G59926);
  nor U43986(n41394,n36374,n38499);
  nand U43987(n38499,n41398,n41393);
  nor U43988(n41393,n40968,n40888);
  not U43989(n40888,n34859);
  xor U43990(n34859,n41399,n41400);
  xnor U43991(n40968,n41401,n41402);
  nor U43992(n41402,n41399,n41400);
  and U43993(n41400,n41403,n41404);
  nand U43994(n41404,n41405,n41406);
  or U43995(n41406,n41407,n41408);
  not U43996(n41405,n41409);
  nand U43997(n41403,n41408,n41407);
  and U43998(n41399,n41410,n41411,n41412);
  nand U43999(n41412,G60013,n34900);
  nand U44000(n41411,n39746,n34898);
  xnor U44001(n39746,n39748,n40750);
  nand U44002(n41410,n36217,G60008);
  nand U44003(n41401,n41413,n41414,n41415);
  nand U44004(n41415,n34898,n39745);
  not U44005(n39745,n40359);
  nor U44006(n40359,n40046,n40129,n41416);
  nor U44007(n41416,n40751,n39748);
  nor U44008(n40129,n40751,G60013);
  not U44009(n40751,G60012);
  not U44010(n40046,n39986);
  nand U44011(n39986,n39748,n39823);
  nor U44012(n39823,n40750,G60012);
  not U44013(n40750,G60013);
  nor U44014(n39748,n40439,n40861);
  nand U44015(n41414,G60012,n34900);
  nand U44016(n41413,n36217,G60007);
  nor U44017(n41398,n34883,n34868);
  xor U44018(n34868,n41417,n41408);
  nand U44019(n41408,n41418,n41419);
  nand U44020(n41419,n40761,n41420);
  xnor U44021(n41420,n39059,n41421);
  nor U44022(n41421,n35398,n39057);
  nand U44023(n35398,n41422,n41423);
  nand U44024(n41423,G59876,n36229);
  not U44025(n36229,G60047);
  or U44026(n41422,G59876,G60206);
  not U44027(n39059,G60017);
  nand U44028(n41418,n39070,n36217);
  xnor U44029(n41417,n41409,n41407);
  nand U44030(n41407,n41424,n41425,n41426);
  nand U44031(n41426,G60014,n34900);
  nand U44032(n41425,n40438,n34898);
  not U44033(n40438,n40591);
  nor U44034(n40591,n39667,n39592);
  nor U44035(n39592,n40439,G60014);
  nor U44036(n39667,n40861,G60015);
  not U44037(n40861,G60014);
  nand U44038(n41424,n36217,G60009);
  nand U44039(n34883,n41427,n41409);
  nand U44040(n41409,n41428,n41429);
  or U44041(n41427,n41429,n41428);
  nand U44042(n41428,n41430,n41431,G59875);
  nand U44043(n41431,n40749,n34924);
  nand U44044(n34924,n38712,n35692,n39070);
  nor U44045(n39070,n40685,n35994);
  not U44046(n35994,n34911);
  nand U44047(n34911,n41432,n41433,n41434,n41435);
  nor U44048(n41435,n41436,n41437,n41438,n41439);
  nor U44049(n41439,n41248,n36896);
  not U44050(n36896,G59988);
  nor U44051(n41438,n41249,n36895);
  not U44052(n36895,G59980);
  nor U44053(n41437,n41250,n36890);
  not U44054(n36890,G59972);
  nor U44055(n41436,n41251,n36888);
  not U44056(n36888,G59956);
  nor U44057(n41434,n41440,n41441,n41442,n41443);
  nor U44058(n41443,n41256,n36887);
  not U44059(n36887,G59948);
  nor U44060(n41442,n41257,n36882);
  not U44061(n36882,G59940);
  nor U44062(n41441,n41258,n36880);
  not U44063(n36880,G59924);
  nor U44064(n41440,n41259,n36879);
  not U44065(n36879,G59916);
  nor U44066(n41433,n41444,n41445,n41446,n41447);
  nor U44067(n41447,n41264,n36874);
  not U44068(n36874,G59908);
  nor U44069(n41446,n41265,n36872);
  not U44070(n36872,G59892);
  nor U44071(n41445,n41266,n36871);
  not U44072(n36871,G59884);
  nor U44073(n41444,n41267,n36898);
  not U44074(n36898,G60004);
  nor U44075(n41432,n41448,n41449,n41450,n41451);
  nor U44076(n41451,n41272,n36897);
  not U44077(n36897,G59996);
  nor U44078(n41450,n41273,n36889);
  not U44079(n36889,G59964);
  nor U44080(n41449,n41274,n36881);
  not U44081(n36881,G59932);
  nor U44082(n41448,n41275,n36873);
  not U44083(n36873,G59900);
  nand U44084(n40685,n41452,n41453,n41454,n41455);
  nor U44085(n41455,n41456,n41457,n41458,n41459);
  nor U44086(n41459,n41248,n37178);
  not U44087(n37178,G59984);
  nor U44088(n41458,n41249,n37177);
  not U44089(n37177,G59976);
  nor U44090(n41457,n41250,n37188);
  not U44091(n37188,G59968);
  nor U44092(n41456,n41251,n37186);
  not U44093(n37186,G59952);
  nor U44094(n41454,n41460,n41461,n41462,n41463);
  nor U44095(n41463,n41256,n37185);
  not U44096(n37185,G59944);
  nor U44097(n41462,n41257,n36562);
  not U44098(n36562,G59936);
  nor U44099(n41461,n41258,n36560);
  not U44100(n36560,G59920);
  nor U44101(n41460,n41259,n36559);
  not U44102(n36559,G59912);
  nor U44103(n41453,n41464,n41465,n41466,n41467);
  nor U44104(n41467,n41264,n36554);
  not U44105(n36554,G59904);
  nor U44106(n41466,n41265,n36552);
  not U44107(n36552,G59888);
  nor U44108(n41465,n41266,n36551);
  not U44109(n36551,G59880);
  nor U44110(n41464,n41267,n37180);
  not U44111(n37180,G60000);
  nor U44112(n41452,n41468,n41469,n41470,n41471);
  nor U44113(n41471,n41272,n37179);
  not U44114(n37179,G59992);
  nor U44115(n41470,n41273,n37187);
  not U44116(n37187,G59960);
  nor U44117(n41469,n41274,n36561);
  not U44118(n36561,G59928);
  nor U44119(n41468,n41275,n36553);
  not U44120(n36553,G59896);
  nor U44121(n41475,n41476,n41477,n41478,n41479);
  nor U44122(n41479,n41248,n36987);
  not U44123(n36987,G59989);
  nor U44124(n41478,n41249,n36983);
  not U44125(n36983,G59981);
  nor U44126(n41477,n41250,n36978);
  not U44127(n36978,G59973);
  nor U44128(n41476,n41251,n36976);
  not U44129(n36976,G59957);
  nor U44130(n41474,n41480,n41481,n41482,n41483);
  nor U44131(n41483,n41256,n36974);
  not U44132(n36974,G59949);
  nor U44133(n41482,n41257,n36968);
  not U44134(n36968,G59941);
  nor U44135(n41481,n41258,n36966);
  not U44136(n36966,G59925);
  nor U44137(n41480,n41259,n36964);
  not U44138(n36964,G59917);
  nor U44139(n41473,n41484,n41485,n41486,n41487);
  nor U44140(n41487,n41264,n36956);
  not U44141(n36956,G59909);
  nor U44142(n41486,n41265,n36952);
  not U44143(n36952,G59893);
  nor U44144(n41485,n41266,n36949);
  not U44145(n36949,G59885);
  nor U44146(n41484,n41267,n36990);
  not U44147(n36990,G60005);
  nor U44148(n41472,n41488,n41489,n41490,n41491);
  nor U44149(n41491,n41272,n36988);
  not U44150(n36988,G59997);
  nor U44151(n41490,n41273,n36977);
  not U44152(n36977,G59965);
  nor U44153(n41489,n41274,n36967);
  not U44154(n36967,G59933);
  nor U44155(n41488,n41275,n36954);
  not U44156(n36954,G59901);
  not U44157(n38712,n35695);
  nand U44158(n35695,n41492,n41493,n41494,n41495);
  nor U44159(n41495,n41496,n41497,n41498,n41499);
  nor U44160(n41499,n41248,n36800);
  not U44161(n36800,G59987);
  nor U44162(n41498,n41249,n36799);
  not U44163(n36799,G59979);
  nor U44164(n41497,n41250,n36794);
  not U44165(n36794,G59971);
  nor U44166(n41496,n41251,n36792);
  not U44167(n36792,G59955);
  nor U44168(n41494,n41500,n41501,n41502,n41503);
  nor U44169(n41503,n41256,n36791);
  not U44170(n36791,G59947);
  nor U44171(n41502,n41257,n36786);
  not U44172(n36786,G59939);
  nor U44173(n41501,n41258,n36784);
  not U44174(n36784,G59923);
  nor U44175(n41500,n41259,n36783);
  not U44176(n36783,G59915);
  nor U44177(n41493,n41504,n41505,n41506,n41507);
  nor U44178(n41507,n41264,n36778);
  not U44179(n36778,G59907);
  nor U44180(n41506,n41265,n36776);
  not U44181(n36776,G59891);
  nor U44182(n41505,n41266,n36775);
  not U44183(n36775,G59883);
  nor U44184(n41504,n41267,n36802);
  not U44185(n36802,G60003);
  nor U44186(n41492,n41508,n41509,n41510,n41511);
  nor U44187(n41511,n41272,n36801);
  not U44188(n36801,G59995);
  nor U44189(n41510,n41273,n36793);
  not U44190(n36793,G59963);
  nor U44191(n41509,n41274,n36785);
  not U44192(n36785,G59931);
  nor U44193(n41508,n41275,n36777);
  not U44194(n36777,G59899);
  nand U44195(n41430,n35414,n41512);
  nand U44196(n41512,G59877,n39057);
  not U44197(n39057,G60016);
  not U44198(n35414,n36217);
  nand U44199(n41429,n36216,n41513,n41514,n41515);
  nand U44200(n41515,n34898,n40439);
  not U44201(n40439,G60015);
  nand U44202(n41514,G60015,n34900);
  nor U44203(n34900,n34898,G59877);
  nand U44204(n41513,n36217,G60010);
  nor U44205(n36217,n35385,G59876);
  not U44206(n36374,G59894);
  nor U44207(n41362,n35542,n41054,n41336);
  not U44208(n41336,n41322);
  nor U44209(n41322,G59876,G59874);
  not U44210(n41054,n35388);
  nand U44211(n35388,n41516,n41517,n41518,n41519);
  nor U44212(n41519,n41520,n41521,n41522,n41523);
  nor U44213(n41523,n41248,n36477);
  not U44214(n36477,G59983);
  nor U44215(n41522,n41249,n36475);
  not U44216(n36475,G59975);
  nor U44217(n41521,n41250,n36469);
  not U44218(n36469,G59967);
  nor U44219(n41520,n41251,n36465);
  not U44220(n36465,G59951);
  nor U44221(n41518,n41524,n41525,n41526,n41527);
  nor U44222(n41527,n41256,n36463);
  not U44223(n36463,G59943);
  nor U44224(n41526,n41257,n36458);
  not U44225(n36458,G59935);
  nor U44226(n41525,n41258,n36456);
  not U44227(n36456,G59919);
  nor U44228(n41524,n41259,n36455);
  not U44229(n36455,G59911);
  nor U44230(n41517,n41528,n41529,n41530,n41531);
  nor U44231(n41531,n41264,n36450);
  not U44232(n36450,G59903);
  nor U44233(n41530,n41265,n36448);
  not U44234(n36448,G59887);
  nor U44235(n41529,n41266,n36447);
  not U44236(n36447,G59879);
  nor U44237(n41528,n41267,n36481);
  not U44238(n36481,G59999);
  nor U44239(n41516,n41532,n41533,n41534,n41535);
  nor U44240(n41535,n41272,n36479);
  not U44241(n36479,G59991);
  nor U44242(n41534,n41273,n36467);
  not U44243(n36467,G59959);
  nor U44244(n41533,n41274,n36457);
  not U44245(n36457,G59927);
  nor U44246(n41532,n41275,n36449);
  not U44247(n36449,G59895);
  not U44248(n35542,n35541);
  nand U44249(n35541,n41536,n41537,n41538,n41539);
  nor U44250(n41539,n41540,n41541,n41542,n41543);
  nor U44251(n41543,n41248,n37343);
  not U44252(n37343,G59986);
  nand U44253(n41248,n41234,n38193);
  nor U44254(n41542,n41249,n37342);
  not U44255(n37342,G59978);
  nand U44256(n41249,n38192,n41234);
  nor U44257(n41541,n41250,n37353);
  not U44258(n37353,G59970);
  nand U44259(n41250,n38201,n38220);
  nor U44260(n41540,n41251,n37351);
  not U44261(n37351,G59954);
  nand U44262(n41251,n38220,n38193);
  nor U44263(n41538,n41544,n41545,n41546,n41547);
  nor U44264(n41547,n41256,n37350);
  not U44265(n37350,G59946);
  nand U44266(n41256,n38192,n38220);
  nor U44267(n41546,n41257,n36717);
  not U44268(n36717,G59938);
  nand U44269(n41257,n38218,n38201);
  nor U44270(n41545,n41258,n36715);
  not U44271(n36715,G59922);
  nand U44272(n41258,n38218,n38193);
  nor U44273(n41544,n41259,n36714);
  not U44274(n36714,G59914);
  nand U44275(n41259,n38218,n38192);
  nor U44276(n41537,n41548,n41549,n41550,n41551);
  nor U44277(n41551,n41264,n36709);
  not U44278(n36709,G59906);
  nand U44279(n41264,n40949,n38201);
  nor U44280(n41550,n41265,n36707);
  not U44281(n36707,G59890);
  nand U44282(n41265,n40949,n38193);
  nor U44283(n38193,n38219,G60010);
  nor U44284(n41549,n41266,n36706);
  not U44285(n36706,G59882);
  nand U44286(n41266,n40949,n38192);
  nor U44287(n38192,n36985,n38219);
  not U44288(n38219,G60009);
  nor U44289(n41548,n41267,n37345);
  not U44290(n37345,G60002);
  nand U44291(n41267,n41234,n38201);
  nor U44292(n38201,G60009,G60010);
  nor U44293(n41536,n41552,n41553,n41554,n41555);
  nor U44294(n41555,n41272,n37344);
  not U44295(n37344,G59994);
  nand U44296(n41272,n38200,n41234);
  nor U44297(n41234,G60008,G60007);
  nor U44298(n41554,n41273,n37352);
  not U44299(n37352,G59962);
  nand U44300(n41273,n38200,n38220);
  nor U44301(n38220,n40879,G60007);
  nor U44302(n41553,n41274,n36716);
  not U44303(n36716,G59930);
  nand U44304(n41274,n38200,n38218);
  nor U44305(n38218,n38831,G60008);
  nor U44306(n41552,n41275,n36708);
  not U44307(n36708,G59898);
  nand U44308(n41275,n38200,n40949);
  nor U44309(n40949,n38831,n40879);
  not U44310(n40879,G60008);
  not U44311(n38831,G60007);
  nor U44312(n38200,n36985,G60009);
  not U44313(n36985,G60010);
  nand U44314(n41300,G60006,G59874);
  nand U44315(n34873,G59874,n35385);
  not U44316(n40771,n39372);
  nor U44317(n39372,n35385,n36216);
  not U44318(n36216,n40761);
  nor U44319(n40761,n40749,n34898);
  not U44320(n34898,G59875);
  not U44321(n40749,G59876);
  not U44322(n35385,G59877);
  nor U44323(G14370,n34831,n35012);
  not U44324(n35012,G59873);
  nor U44325(G14369,n34831,n35011);
  not U44326(n35011,G59872);
  nor U44327(G14368,n34831,n35010);
  not U44328(n35010,G59871);
  nor U44329(G14367,n34831,n35009);
  not U44330(n35009,G59870);
  nor U44331(G14366,n34831,n35008);
  not U44332(n35008,G59869);
  nor U44333(G14365,n34831,n35007);
  not U44334(n35007,G59868);
  nor U44335(G14364,n34831,n35006);
  not U44336(n35006,G59867);
  nor U44337(G14363,n34831,n35005);
  not U44338(n35005,G59866);
  nor U44339(G14362,n34831,n35004);
  not U44340(n35004,G59865);
  nor U44341(G14361,n34831,n35003);
  not U44342(n35003,G59864);
  nor U44343(G14360,n34831,n35002);
  not U44344(n35002,G59863);
  nor U44345(G14359,n34831,n35001);
  not U44346(n35001,G59862);
  nor U44347(G14358,n34831,n35000);
  not U44348(n35000,G59861);
  nor U44349(G14357,n34831,n34999);
  not U44350(n34999,G59860);
  nor U44351(G14356,n34831,n34998);
  not U44352(n34998,G59859);
  nor U44353(G14355,n34831,n34997);
  not U44354(n34997,G59858);
  and U44355(G14354,n34832,G59857);
  and U44356(G14353,n34832,G59856);
  and U44357(G14352,n34832,G59855);
  and U44358(G14351,n34832,G59854);
  and U44359(G14350,n34832,G59853);
  and U44360(G14349,n34832,G59852);
  and U44361(G14348,n34832,G59851);
  and U44362(G14347,n34832,G59850);
  nor U44363(G14346,n34831,n35018);
  not U44364(n35018,G59849);
  nor U44365(G14345,n34831,n35017);
  not U44366(n35017,G59848);
  nor U44367(G14344,n34831,n35016);
  not U44368(n35016,G59847);
  nor U44369(G14343,n34831,n35015);
  not U44370(n35015,G59846);
  and U44371(G14342,n34832,G59845);
  and U44372(G14341,n34832,G59844);
  not U44373(n34832,n34831);
  nand U44374(n34831,n41556,n41557);
  nand U44375(n41557,G59841,n41558);
  nand U44376(G14340,n41559,n41560,n41561,n41562);
  nor U44377(n41562,n41563,n34836,n41564);
  nor U44378(n41564,n41230,n34899);
  not U44379(n41230,n41558);
  nor U44380(n34836,G59841,G59839);
  nor U44381(n41563,n27739,n41556);
  nand U44382(n41561,n34820,n34891);
  nand U44383(n41560,n41565,n34951);
  nand U44384(n41559,G59841,G33,G59840);
  nand U44385(G14339,n41566,n41567,n41568,n41569);
  nand U44386(n41569,n41558,G33);
  nor U44387(n41558,n34951,G59839);
  nor U44388(n41568,n41570,n41571);
  nor U44389(n41571,n34891,n41565,n35895);
  nor U44390(n41565,n41572,n27747);
  or U44391(n41567,n41556,n41572);
  nand U44392(n41556,n34951,n35895);
  nand U44393(n41566,n35790,G59840);
  nand U44394(G14338,n41573,n41574,n41575,n41576);
  nand U44395(n41576,G59839,n27739,n35895);
  not U44396(n35895,G59841);
  nand U44397(n41575,G33,n41577,G59841);
  nand U44398(n41577,n41572,n41578);
  nand U44399(n41578,n34951,n34891);
  not U44400(n41574,n41579);
  nand U44401(n41573,G59840,n41580,n35790);
  not U44402(n35790,n34899);
  nand U44403(n34899,G58906,G36);
  nand U44404(n41580,n41572,n41581);
  nand U44405(n41581,n41582,n27739,G59841);
  not U44406(n27739,G34);
  nand U44407(n41582,n34891,n27747);
  not U44408(n27747,G33);
  not U44409(n34891,G60247);
  nand U44410(G14337,n41583,n41584,n41585);
  nand U44411(n41585,G59838,n34820);
  nand U44412(n41584,n41579,G60208);
  nand U44413(n41583,n41570,G60209);
  nand U44414(G14336,n41586,n41587,n41588);
  nand U44415(n41588,G59837,n34820);
  nand U44416(n41587,n41579,G60209);
  nand U44417(n41586,n41570,G60210);
  nand U44418(G14335,n41589,n41590,n41591);
  nand U44419(n41591,G59836,n34820);
  nand U44420(n41590,n41579,G60210);
  nand U44421(n41589,n41570,G60211);
  nand U44422(G14334,n41592,n41593,n41594);
  nand U44423(n41594,G59835,n34820);
  nand U44424(n41593,n41579,G60211);
  nand U44425(n41592,n41570,G60212);
  nand U44426(G14333,n41595,n41596,n41597);
  nand U44427(n41597,G59834,n34820);
  nand U44428(n41596,n41579,G60212);
  nand U44429(n41595,n41570,G60213);
  nand U44430(G14332,n41598,n41599,n41600);
  nand U44431(n41600,G59833,n34820);
  nand U44432(n41599,n41579,G60213);
  nand U44433(n41598,n41570,G60214);
  nand U44434(G14331,n41601,n41602,n41603);
  nand U44435(n41603,G59832,n34820);
  nand U44436(n41602,n41579,G60214);
  nand U44437(n41601,n41570,G60215);
  nand U44438(G14330,n41604,n41605,n41606);
  nand U44439(n41606,G59831,n34820);
  nand U44440(n41605,n41579,G60215);
  nand U44441(n41604,n41570,G60216);
  nand U44442(G14329,n41607,n41608,n41609);
  nand U44443(n41609,G59830,n34820);
  nand U44444(n41608,n41579,G60216);
  nand U44445(n41607,n41570,G60217);
  nand U44446(G14328,n41610,n41611,n41612);
  nand U44447(n41612,G59829,n34820);
  nand U44448(n41611,n41579,G60217);
  nand U44449(n41610,n41570,G60218);
  nand U44450(G14327,n41613,n41614,n41615);
  nand U44451(n41615,G59828,n34820);
  nand U44452(n41614,n41579,G60218);
  nand U44453(n41613,n41570,G60219);
  nand U44454(G14326,n41616,n41617,n41618);
  nand U44455(n41618,G59827,n34820);
  nand U44456(n41617,n41579,G60219);
  nand U44457(n41616,n41570,G60220);
  nand U44458(G14325,n41619,n41620,n41621);
  nand U44459(n41621,G59826,n34820);
  nand U44460(n41620,n41579,G60220);
  nand U44461(n41619,n41570,G60221);
  nand U44462(G14324,n41622,n41623,n41624);
  nand U44463(n41624,G59825,n34820);
  nand U44464(n41623,n41579,G60221);
  nand U44465(n41622,n41570,G60222);
  nand U44466(G14323,n41625,n41626,n41627);
  nand U44467(n41627,G59824,n34820);
  nand U44468(n41626,n41579,G60222);
  nand U44469(n41625,n41570,G60223);
  nand U44470(G14322,n41628,n41629,n41630);
  nand U44471(n41630,G59823,n34820);
  nand U44472(n41629,n41579,G60223);
  nand U44473(n41628,n41570,G60224);
  nand U44474(G14321,n41631,n41632,n41633);
  nand U44475(n41633,G59822,n34820);
  nand U44476(n41632,n41579,G60224);
  nand U44477(n41631,n41570,G60225);
  nand U44478(G14320,n41634,n41635,n41636);
  nand U44479(n41636,G59821,n34820);
  nand U44480(n41635,n41579,G60225);
  nand U44481(n41634,n41570,G60226);
  nand U44482(G14319,n41637,n41638,n41639);
  nand U44483(n41639,G59820,n34820);
  nand U44484(n41638,n41579,G60226);
  nand U44485(n41637,n41570,G60227);
  nand U44486(G14318,n41640,n41641,n41642);
  nand U44487(n41642,G59819,n34820);
  nand U44488(n41641,n41579,G60227);
  nand U44489(n41640,n41570,G60228);
  nand U44490(G14317,n41643,n41644,n41645);
  nand U44491(n41645,G59818,n34820);
  nand U44492(n41644,n41579,G60228);
  nand U44493(n41643,n41570,G60229);
  nand U44494(G14316,n41646,n41647,n41648);
  nand U44495(n41648,G59817,n34820);
  nand U44496(n41647,n41579,G60229);
  nand U44497(n41646,n41570,G60230);
  nand U44498(G14315,n41649,n41650,n41651);
  nand U44499(n41651,G59816,n34820);
  nand U44500(n41650,n41579,G60230);
  nand U44501(n41649,n41570,G60231);
  nand U44502(G14314,n41652,n41653,n41654);
  nand U44503(n41654,G59815,n34820);
  nand U44504(n41653,n41579,G60231);
  nand U44505(n41652,n41570,G60232);
  nand U44506(G14313,n41655,n41656,n41657);
  nand U44507(n41657,G59814,n34820);
  nand U44508(n41656,n41579,G60232);
  nand U44509(n41655,n41570,G60233);
  nand U44510(G14312,n41658,n41659,n41660);
  nand U44511(n41660,G59813,n34820);
  nand U44512(n41659,n41579,G60233);
  nand U44513(n41658,n41570,G60234);
  nand U44514(G14311,n41661,n41662,n41663);
  nand U44515(n41663,G59812,n34820);
  nand U44516(n41662,n41579,G60234);
  nand U44517(n41661,n41570,G60235);
  nand U44518(G14310,n41664,n41665,n41666);
  nand U44519(n41666,G59811,n34820);
  nand U44520(n41665,n41579,G60235);
  nand U44521(n41664,n41570,G60236);
  nand U44522(G14309,n41667,n41668,n41669);
  nand U44523(n41669,G59810,n34820);
  nand U44524(n41668,n41579,G60236);
  nand U44525(n41667,n41570,G60237);
  nand U44526(G14308,n41670,n41671,n41672);
  nand U44527(n41672,G59809,n34820);
  nand U44528(n41671,n41579,G60237);
  not U44529(n41572,G59839);
  nand U44530(n41670,n41570,G60238);
  nor U44531(n34821,n34951,G59841);
  not U44532(n34951,G59840);
endmodule

