//  File   : pp2.v
//  Created: Tue Mar  1 13:59:58 2011
//  By     : lsdb version V2.9.00 (02/28/11 ) Linux_AMD64_E4
//           lsdb -verilog vip_pg_edt_controller.x
//           sdb version 330
//
//  (c) 1991-2011, SynTest Technologies, Inc.

module vip_pg_edt_controller.x ( edt_channels_out_from_controller_0 , edt_channels_out_from_controller_1 , edt_channels_out_from_controller_2 , edt_channels_out_from_controller_3 ,
        edt_channels_out_from_controller_4 , edt_channels_out_from_controller_5 , edt_channels_out_from_controller_6 , edt_channels_out_from_controller_7 ,
        edt_channels_out_from_controller_8 , edt_channels_out_from_controller_9 , edt_channels_out_from_controller_10 , edt_channels_out_from_controller_11 ,
        edt_channels_out_from_controller_12 , edt_channels_out_from_controller_13 , edt_channels_out_from_controller_14 , masks_for_compactor_0_0 ,
        masks_for_compactor_0_1 , masks_for_compactor_0_2 , masks_for_compactor_0_3 , masks_for_compactor_0_4 ,
        masks_for_compactor_0_5 , masks_for_compactor_0_6 , masks_for_compactor_0_7 , masks_for_compactor_0_8 ,
        masks_for_compactor_0_9 , masks_for_compactor_0_10 , masks_for_compactor_0_11 , masks_for_compactor_0_12 ,
        masks_for_compactor_0_13 , masks_for_compactor_0_14 , masks_for_compactor_0_15 , masks_for_compactor_0_16 ,
        masks_for_compactor_0_17 , masks_for_compactor_0_18 , masks_for_compactor_0_19 , masks_for_compactor_0_20 ,
        masks_for_compactor_0_21 , masks_for_compactor_0_22 , masks_for_compactor_0_23 , masks_for_compactor_0_24 ,
        masks_for_compactor_0_25 , masks_for_compactor_0_26 , masks_for_compactor_0_27 , masks_for_compactor_0_28 ,
        masks_for_compactor_0_29 , masks_for_compactor_0_30 , masks_for_compactor_0_31 , masks_for_compactor_0_32 ,
        masks_for_compactor_0_33 , masks_for_compactor_0_34 , masks_for_compactor_0_35 , masks_for_compactor_0_36 ,
        masks_for_compactor_0_37 , masks_for_compactor_0_38 , masks_for_compactor_0_39 , masks_for_compactor_0_40 ,
        masks_for_compactor_0_41 , masks_for_compactor_0_42 , masks_for_compactor_0_43 , masks_for_compactor_0_44 ,
        masks_for_compactor_0_45 , masks_for_compactor_0_46 , masks_for_compactor_0_47 , masks_for_compactor_0_48 ,
        masks_for_compactor_0_49 , masks_for_compactor_0_50 , masks_for_compactor_0_51 , masks_for_compactor_0_52 ,
        masks_for_compactor_0_53 , masks_for_compactor_1_0 , masks_for_compactor_1_1 , masks_for_compactor_1_2 ,
        masks_for_compactor_1_3 , masks_for_compactor_1_4 , masks_for_compactor_1_5 , masks_for_compactor_1_6 ,
        masks_for_compactor_1_7 , masks_for_compactor_1_8 , masks_for_compactor_1_9 , masks_for_compactor_1_10 ,
        masks_for_compactor_1_11 , masks_for_compactor_1_12 , masks_for_compactor_1_13 , masks_for_compactor_1_14 ,
        masks_for_compactor_1_15 , masks_for_compactor_1_16 , masks_for_compactor_1_17 , masks_for_compactor_1_18 ,
        masks_for_compactor_1_19 , masks_for_compactor_1_20 , masks_for_compactor_1_21 , masks_for_compactor_1_22 ,
        masks_for_compactor_1_23 , masks_for_compactor_1_24 , masks_for_compactor_1_25 , masks_for_compactor_1_26 ,
        masks_for_compactor_1_27 , masks_for_compactor_1_28 , masks_for_compactor_1_29 , masks_for_compactor_1_30 ,
        masks_for_compactor_1_31 , masks_for_compactor_1_32 , masks_for_compactor_1_33 , masks_for_compactor_1_34 ,
        masks_for_compactor_1_35 , masks_for_compactor_1_36 , masks_for_compactor_1_37 , masks_for_compactor_1_38 ,
        masks_for_compactor_1_39 , masks_for_compactor_1_40 , masks_for_compactor_1_41 , masks_for_compactor_1_42 ,
        masks_for_compactor_1_43 , masks_for_compactor_1_44 , masks_for_compactor_1_45 , masks_for_compactor_1_46 ,
        masks_for_compactor_1_47 , masks_for_compactor_1_48 , masks_for_compactor_1_49 , masks_for_compactor_1_50 ,
        masks_for_compactor_1_51 , masks_for_compactor_1_52 , masks_for_compactor_2_0 , masks_for_compactor_2_1 ,
        masks_for_compactor_2_2 , masks_for_compactor_2_3 , masks_for_compactor_2_4 , masks_for_compactor_2_5 ,
        masks_for_compactor_2_6 , masks_for_compactor_2_7 , masks_for_compactor_2_8 , masks_for_compactor_2_9 ,
        masks_for_compactor_2_10 , masks_for_compactor_2_11 , masks_for_compactor_2_12 , masks_for_compactor_2_13 ,
        masks_for_compactor_2_14 , masks_for_compactor_2_15 , masks_for_compactor_2_16 , masks_for_compactor_2_17 ,
        masks_for_compactor_2_18 , masks_for_compactor_2_19 , masks_for_compactor_2_20 , masks_for_compactor_2_21 ,
        masks_for_compactor_2_22 , masks_for_compactor_2_23 , masks_for_compactor_2_24 , masks_for_compactor_2_25 ,
        masks_for_compactor_2_26 , masks_for_compactor_2_27 , masks_for_compactor_2_28 , masks_for_compactor_2_29 ,
        masks_for_compactor_2_30 , masks_for_compactor_2_31 , masks_for_compactor_2_32 , masks_for_compactor_2_33 ,
        masks_for_compactor_2_34 , masks_for_compactor_2_35 , masks_for_compactor_2_36 , masks_for_compactor_2_37 ,
        masks_for_compactor_2_38 , masks_for_compactor_2_39 , masks_for_compactor_2_40 , masks_for_compactor_2_41 ,
        masks_for_compactor_2_42 , masks_for_compactor_2_43 , masks_for_compactor_2_44 , masks_for_compactor_2_45 ,
        masks_for_compactor_2_46 , masks_for_compactor_2_47 , masks_for_compactor_2_48 , masks_for_compactor_2_49 ,
        masks_for_compactor_2_50 , masks_for_compactor_2_51 , masks_for_compactor_2_52 , masks_for_compactor_3_0 ,
        masks_for_compactor_3_1 , masks_for_compactor_3_2 , masks_for_compactor_3_3 , masks_for_compactor_3_4 ,
        masks_for_compactor_3_5 , masks_for_compactor_3_6 , masks_for_compactor_3_7 , masks_for_compactor_3_8 ,
        masks_for_compactor_3_9 , masks_for_compactor_3_10 , masks_for_compactor_3_11 , masks_for_compactor_3_12 ,
        masks_for_compactor_3_13 , masks_for_compactor_3_14 , masks_for_compactor_3_15 , masks_for_compactor_3_16 ,
        masks_for_compactor_3_17 , masks_for_compactor_3_18 , masks_for_compactor_3_19 , masks_for_compactor_3_20 ,
        masks_for_compactor_3_21 , masks_for_compactor_3_22 , masks_for_compactor_3_23 , masks_for_compactor_3_24 ,
        masks_for_compactor_3_25 , masks_for_compactor_3_26 , masks_for_compactor_3_27 , masks_for_compactor_3_28 ,
        masks_for_compactor_3_29 , masks_for_compactor_3_30 , masks_for_compactor_3_31 , masks_for_compactor_3_32 ,
        masks_for_compactor_3_33 , masks_for_compactor_3_34 , masks_for_compactor_3_35 , masks_for_compactor_3_36 ,
        masks_for_compactor_3_37 , masks_for_compactor_3_38 , masks_for_compactor_3_39 , masks_for_compactor_3_40 ,
        masks_for_compactor_3_41 , masks_for_compactor_3_42 , masks_for_compactor_3_43 , masks_for_compactor_3_44 ,
        masks_for_compactor_3_45 , masks_for_compactor_3_46 , masks_for_compactor_3_47 , masks_for_compactor_3_48 ,
        masks_for_compactor_3_49 , masks_for_compactor_3_50 , masks_for_compactor_3_51 , masks_for_compactor_3_52 ,
        masks_for_compactor_4_0 , masks_for_compactor_4_1 , masks_for_compactor_4_2 , masks_for_compactor_4_3 ,
        masks_for_compactor_4_4 , masks_for_compactor_4_5 , masks_for_compactor_4_6 , masks_for_compactor_4_7 ,
        masks_for_compactor_4_8 , masks_for_compactor_4_9 , masks_for_compactor_4_10 , masks_for_compactor_4_11 ,
        masks_for_compactor_4_12 , masks_for_compactor_4_13 , masks_for_compactor_4_14 , masks_for_compactor_4_15 ,
        masks_for_compactor_4_16 , masks_for_compactor_4_17 , masks_for_compactor_4_18 , masks_for_compactor_4_19 ,
        masks_for_compactor_4_20 , masks_for_compactor_4_21 , masks_for_compactor_4_22 , masks_for_compactor_4_23 ,
        masks_for_compactor_4_24 , masks_for_compactor_4_25 , masks_for_compactor_4_26 , masks_for_compactor_4_27 ,
        masks_for_compactor_4_28 , masks_for_compactor_4_29 , masks_for_compactor_4_30 , masks_for_compactor_4_31 ,
        masks_for_compactor_4_32 , masks_for_compactor_4_33 , masks_for_compactor_4_34 , masks_for_compactor_4_35 ,
        masks_for_compactor_4_36 , masks_for_compactor_4_37 , masks_for_compactor_4_38 , masks_for_compactor_4_39 ,
        masks_for_compactor_4_40 , masks_for_compactor_4_41 , masks_for_compactor_4_42 , masks_for_compactor_4_43 ,
        masks_for_compactor_4_44 , masks_for_compactor_4_45 , masks_for_compactor_4_46 , masks_for_compactor_4_47 ,
        masks_for_compactor_4_48 , masks_for_compactor_4_49 , masks_for_compactor_4_50 , masks_for_compactor_4_51 ,
        masks_for_compactor_4_52 , masks_for_compactor_5_0 , masks_for_compactor_5_1 , masks_for_compactor_5_2 ,
        masks_for_compactor_5_3 , masks_for_compactor_5_4 , masks_for_compactor_5_5 , masks_for_compactor_5_6 ,
        masks_for_compactor_5_7 , masks_for_compactor_5_8 , masks_for_compactor_5_9 , masks_for_compactor_5_10 ,
        masks_for_compactor_5_11 , masks_for_compactor_5_12 , masks_for_compactor_5_13 , masks_for_compactor_5_14 ,
        masks_for_compactor_5_15 , masks_for_compactor_5_16 , masks_for_compactor_5_17 , masks_for_compactor_5_18 ,
        masks_for_compactor_5_19 , masks_for_compactor_5_20 , masks_for_compactor_5_21 , masks_for_compactor_5_22 ,
        masks_for_compactor_5_23 , masks_for_compactor_5_24 , masks_for_compactor_5_25 , masks_for_compactor_5_26 ,
        masks_for_compactor_5_27 , masks_for_compactor_5_28 , masks_for_compactor_5_29 , masks_for_compactor_5_30 ,
        masks_for_compactor_5_31 , masks_for_compactor_5_32 , masks_for_compactor_5_33 , masks_for_compactor_5_34 ,
        masks_for_compactor_5_35 , masks_for_compactor_5_36 , masks_for_compactor_5_37 , masks_for_compactor_5_38 ,
        masks_for_compactor_5_39 , masks_for_compactor_5_40 , masks_for_compactor_5_41 , masks_for_compactor_5_42 ,
        masks_for_compactor_5_43 , masks_for_compactor_5_44 , masks_for_compactor_5_45 , masks_for_compactor_5_46 ,
        masks_for_compactor_5_47 , masks_for_compactor_5_48 , masks_for_compactor_5_49 , masks_for_compactor_5_50 ,
        masks_for_compactor_5_51 , masks_for_compactor_5_52 , masks_for_compactor_6_0 , masks_for_compactor_6_1 ,
        masks_for_compactor_6_2 , masks_for_compactor_6_3 , masks_for_compactor_6_4 , masks_for_compactor_6_5 ,
        masks_for_compactor_6_6 , masks_for_compactor_6_7 , masks_for_compactor_6_8 , masks_for_compactor_6_9 ,
        masks_for_compactor_6_10 , masks_for_compactor_6_11 , masks_for_compactor_6_12 , masks_for_compactor_6_13 ,
        masks_for_compactor_6_14 , masks_for_compactor_6_15 , masks_for_compactor_6_16 , masks_for_compactor_6_17 ,
        masks_for_compactor_6_18 , masks_for_compactor_6_19 , masks_for_compactor_6_20 , masks_for_compactor_6_21 ,
        masks_for_compactor_6_22 , masks_for_compactor_6_23 , masks_for_compactor_6_24 , masks_for_compactor_6_25 ,
        masks_for_compactor_6_26 , masks_for_compactor_6_27 , masks_for_compactor_6_28 , masks_for_compactor_6_29 ,
        masks_for_compactor_6_30 , masks_for_compactor_6_31 , masks_for_compactor_6_32 , masks_for_compactor_6_33 ,
        masks_for_compactor_6_34 , masks_for_compactor_6_35 , masks_for_compactor_6_36 , masks_for_compactor_6_37 ,
        masks_for_compactor_6_38 , masks_for_compactor_6_39 , masks_for_compactor_6_40 , masks_for_compactor_6_41 ,
        masks_for_compactor_6_42 , masks_for_compactor_6_43 , masks_for_compactor_6_44 , masks_for_compactor_6_45 ,
        masks_for_compactor_6_46 , masks_for_compactor_6_47 , masks_for_compactor_6_48 , masks_for_compactor_6_49 ,
        masks_for_compactor_6_50 , masks_for_compactor_6_51 , masks_for_compactor_6_52 , masks_for_compactor_7_0 ,
        masks_for_compactor_7_1 , masks_for_compactor_7_2 , masks_for_compactor_7_3 , masks_for_compactor_7_4 ,
        masks_for_compactor_7_5 , masks_for_compactor_7_6 , masks_for_compactor_7_7 , masks_for_compactor_7_8 ,
        masks_for_compactor_7_9 , masks_for_compactor_7_10 , masks_for_compactor_7_11 , masks_for_compactor_7_12 ,
        masks_for_compactor_7_13 , masks_for_compactor_7_14 , masks_for_compactor_7_15 , masks_for_compactor_7_16 ,
        masks_for_compactor_7_17 , masks_for_compactor_7_18 , masks_for_compactor_7_19 , masks_for_compactor_7_20 ,
        masks_for_compactor_7_21 , masks_for_compactor_7_22 , masks_for_compactor_7_23 , masks_for_compactor_7_24 ,
        masks_for_compactor_7_25 , masks_for_compactor_7_26 , masks_for_compactor_7_27 , masks_for_compactor_7_28 ,
        masks_for_compactor_7_29 , masks_for_compactor_7_30 , masks_for_compactor_7_31 , masks_for_compactor_7_32 ,
        masks_for_compactor_7_33 , masks_for_compactor_7_34 , masks_for_compactor_7_35 , masks_for_compactor_7_36 ,
        masks_for_compactor_7_37 , masks_for_compactor_7_38 , masks_for_compactor_7_39 , masks_for_compactor_7_40 ,
        masks_for_compactor_7_41 , masks_for_compactor_7_42 , masks_for_compactor_7_43 , masks_for_compactor_7_44 ,
        masks_for_compactor_7_45 , masks_for_compactor_7_46 , masks_for_compactor_7_47 , masks_for_compactor_7_48 ,
        masks_for_compactor_7_49 , masks_for_compactor_7_50 , masks_for_compactor_7_51 , masks_for_compactor_7_52 ,
        masks_for_compactor_8_0 , masks_for_compactor_8_1 , masks_for_compactor_8_2 , masks_for_compactor_8_3 ,
        masks_for_compactor_8_4 , masks_for_compactor_8_5 , masks_for_compactor_8_6 , masks_for_compactor_8_7 ,
        masks_for_compactor_8_8 , masks_for_compactor_8_9 , masks_for_compactor_8_10 , masks_for_compactor_8_11 ,
        masks_for_compactor_8_12 , masks_for_compactor_8_13 , masks_for_compactor_8_14 , masks_for_compactor_8_15 ,
        masks_for_compactor_8_16 , masks_for_compactor_8_17 , masks_for_compactor_8_18 , masks_for_compactor_8_19 ,
        masks_for_compactor_8_20 , masks_for_compactor_8_21 , masks_for_compactor_8_22 , masks_for_compactor_8_23 ,
        masks_for_compactor_8_24 , masks_for_compactor_8_25 , masks_for_compactor_8_26 , masks_for_compactor_8_27 ,
        masks_for_compactor_8_28 , masks_for_compactor_8_29 , masks_for_compactor_8_30 , masks_for_compactor_8_31 ,
        masks_for_compactor_8_32 , masks_for_compactor_8_33 , masks_for_compactor_8_34 , masks_for_compactor_8_35 ,
        masks_for_compactor_8_36 , masks_for_compactor_8_37 , masks_for_compactor_8_38 , masks_for_compactor_8_39 ,
        masks_for_compactor_8_40 , masks_for_compactor_8_41 , masks_for_compactor_8_42 , masks_for_compactor_8_43 ,
        masks_for_compactor_8_44 , masks_for_compactor_8_45 , masks_for_compactor_8_46 , masks_for_compactor_8_47 ,
        masks_for_compactor_8_48 , masks_for_compactor_8_49 , masks_for_compactor_8_50 , masks_for_compactor_8_51 ,
        masks_for_compactor_8_52 , masks_for_compactor_9_0 , masks_for_compactor_9_1 , masks_for_compactor_9_2 ,
        masks_for_compactor_9_3 , masks_for_compactor_9_4 , masks_for_compactor_9_5 , masks_for_compactor_9_6 ,
        masks_for_compactor_9_7 , masks_for_compactor_9_8 , masks_for_compactor_9_9 , masks_for_compactor_9_10 ,
        masks_for_compactor_9_11 , masks_for_compactor_9_12 , masks_for_compactor_9_13 , masks_for_compactor_9_14 ,
        masks_for_compactor_9_15 , masks_for_compactor_9_16 , masks_for_compactor_9_17 , masks_for_compactor_9_18 ,
        masks_for_compactor_9_19 , masks_for_compactor_9_20 , masks_for_compactor_9_21 , masks_for_compactor_9_22 ,
        masks_for_compactor_9_23 , masks_for_compactor_9_24 , masks_for_compactor_9_25 , masks_for_compactor_9_26 ,
        masks_for_compactor_9_27 , masks_for_compactor_9_28 , masks_for_compactor_9_29 , masks_for_compactor_9_30 ,
        masks_for_compactor_9_31 , masks_for_compactor_9_32 , masks_for_compactor_9_33 , masks_for_compactor_9_34 ,
        masks_for_compactor_9_35 , masks_for_compactor_9_36 , masks_for_compactor_9_37 , masks_for_compactor_9_38 ,
        masks_for_compactor_9_39 , masks_for_compactor_9_40 , masks_for_compactor_9_41 , masks_for_compactor_9_42 ,
        masks_for_compactor_9_43 , masks_for_compactor_9_44 , masks_for_compactor_9_45 , masks_for_compactor_9_46 ,
        masks_for_compactor_9_47 , masks_for_compactor_9_48 , masks_for_compactor_9_49 , masks_for_compactor_9_50 ,
        masks_for_compactor_9_51 , masks_for_compactor_9_52 , masks_for_compactor_10_0 , masks_for_compactor_10_1 ,
        masks_for_compactor_10_2 , masks_for_compactor_10_3 , masks_for_compactor_10_4 , masks_for_compactor_10_5 ,
        masks_for_compactor_10_6 , masks_for_compactor_10_7 , masks_for_compactor_10_8 , masks_for_compactor_10_9 ,
        masks_for_compactor_10_10 , masks_for_compactor_10_11 , masks_for_compactor_10_12 , masks_for_compactor_10_13 ,
        masks_for_compactor_10_14 , masks_for_compactor_10_15 , masks_for_compactor_10_16 , masks_for_compactor_10_17 ,
        masks_for_compactor_10_18 , masks_for_compactor_10_19 , masks_for_compactor_10_20 , masks_for_compactor_10_21 ,
        masks_for_compactor_10_22 , masks_for_compactor_10_23 , masks_for_compactor_10_24 , masks_for_compactor_10_25 ,
        masks_for_compactor_10_26 , masks_for_compactor_10_27 , masks_for_compactor_10_28 , masks_for_compactor_10_29 ,
        masks_for_compactor_10_30 , masks_for_compactor_10_31 , masks_for_compactor_10_32 , masks_for_compactor_10_33 ,
        masks_for_compactor_10_34 , masks_for_compactor_10_35 , masks_for_compactor_10_36 , masks_for_compactor_10_37 ,
        masks_for_compactor_10_38 , masks_for_compactor_10_39 , masks_for_compactor_10_40 , masks_for_compactor_10_41 ,
        masks_for_compactor_10_42 , masks_for_compactor_10_43 , masks_for_compactor_10_44 , masks_for_compactor_10_45 ,
        masks_for_compactor_10_46 , masks_for_compactor_10_47 , masks_for_compactor_10_48 , masks_for_compactor_10_49 ,
        masks_for_compactor_10_50 , masks_for_compactor_10_51 , masks_for_compactor_10_52 , masks_for_compactor_11_0 ,
        masks_for_compactor_11_1 , masks_for_compactor_11_2 , masks_for_compactor_11_3 , masks_for_compactor_11_4 ,
        masks_for_compactor_11_5 , masks_for_compactor_11_6 , masks_for_compactor_11_7 , masks_for_compactor_11_8 ,
        masks_for_compactor_11_9 , masks_for_compactor_11_10 , masks_for_compactor_11_11 , masks_for_compactor_11_12 ,
        masks_for_compactor_11_13 , masks_for_compactor_11_14 , masks_for_compactor_11_15 , masks_for_compactor_11_16 ,
        masks_for_compactor_11_17 , masks_for_compactor_11_18 , masks_for_compactor_11_19 , masks_for_compactor_11_20 ,
        masks_for_compactor_11_21 , masks_for_compactor_11_22 , masks_for_compactor_11_23 , masks_for_compactor_11_24 ,
        masks_for_compactor_11_25 , masks_for_compactor_11_26 , masks_for_compactor_11_27 , masks_for_compactor_11_28 ,
        masks_for_compactor_11_29 , masks_for_compactor_11_30 , masks_for_compactor_11_31 , masks_for_compactor_11_32 ,
        masks_for_compactor_11_33 , masks_for_compactor_11_34 , masks_for_compactor_11_35 , masks_for_compactor_11_36 ,
        masks_for_compactor_11_37 , masks_for_compactor_11_38 , masks_for_compactor_11_39 , masks_for_compactor_11_40 ,
        masks_for_compactor_11_41 , masks_for_compactor_11_42 , masks_for_compactor_11_43 , masks_for_compactor_11_44 ,
        masks_for_compactor_11_45 , masks_for_compactor_11_46 , masks_for_compactor_11_47 , masks_for_compactor_11_48 ,
        masks_for_compactor_11_49 , masks_for_compactor_11_50 , masks_for_compactor_11_51 , masks_for_compactor_11_52 ,
        masks_for_compactor_12_0 , masks_for_compactor_12_1 , masks_for_compactor_12_2 , masks_for_compactor_12_3 ,
        masks_for_compactor_12_4 , masks_for_compactor_12_5 , masks_for_compactor_12_6 , masks_for_compactor_12_7 ,
        masks_for_compactor_12_8 , masks_for_compactor_12_9 , masks_for_compactor_12_10 , masks_for_compactor_12_11 ,
        masks_for_compactor_12_12 , masks_for_compactor_12_13 , masks_for_compactor_12_14 , masks_for_compactor_12_15 ,
        masks_for_compactor_12_16 , masks_for_compactor_12_17 , masks_for_compactor_12_18 , masks_for_compactor_12_19 ,
        masks_for_compactor_12_20 , masks_for_compactor_12_21 , masks_for_compactor_12_22 , masks_for_compactor_12_23 ,
        masks_for_compactor_12_24 , masks_for_compactor_12_25 , masks_for_compactor_12_26 , masks_for_compactor_12_27 ,
        masks_for_compactor_12_28 , masks_for_compactor_12_29 , masks_for_compactor_12_30 , masks_for_compactor_12_31 ,
        masks_for_compactor_12_32 , masks_for_compactor_12_33 , masks_for_compactor_12_34 , masks_for_compactor_12_35 ,
        masks_for_compactor_12_36 , masks_for_compactor_12_37 , masks_for_compactor_12_38 , masks_for_compactor_12_39 ,
        masks_for_compactor_12_40 , masks_for_compactor_12_41 , masks_for_compactor_12_42 , masks_for_compactor_12_43 ,
        masks_for_compactor_12_44 , masks_for_compactor_12_45 , masks_for_compactor_12_46 , masks_for_compactor_12_47 ,
        masks_for_compactor_12_48 , masks_for_compactor_12_49 , masks_for_compactor_12_50 , masks_for_compactor_12_51 ,
        masks_for_compactor_12_52 , masks_for_compactor_13_0 , masks_for_compactor_13_1 , masks_for_compactor_13_2 ,
        masks_for_compactor_13_3 , masks_for_compactor_13_4 , masks_for_compactor_13_5 , masks_for_compactor_13_6 ,
        masks_for_compactor_13_7 , masks_for_compactor_13_8 , masks_for_compactor_13_9 , masks_for_compactor_13_10 ,
        masks_for_compactor_13_11 , masks_for_compactor_13_12 , masks_for_compactor_13_13 , masks_for_compactor_13_14 ,
        masks_for_compactor_13_15 , masks_for_compactor_13_16 , masks_for_compactor_13_17 , masks_for_compactor_13_18 ,
        masks_for_compactor_13_19 , masks_for_compactor_13_20 , masks_for_compactor_13_21 , masks_for_compactor_13_22 ,
        masks_for_compactor_13_23 , masks_for_compactor_13_24 , masks_for_compactor_13_25 , masks_for_compactor_13_26 ,
        masks_for_compactor_13_27 , masks_for_compactor_13_28 , masks_for_compactor_13_29 , masks_for_compactor_13_30 ,
        masks_for_compactor_13_31 , masks_for_compactor_13_32 , masks_for_compactor_13_33 , masks_for_compactor_13_34 ,
        masks_for_compactor_13_35 , masks_for_compactor_13_36 , masks_for_compactor_13_37 , masks_for_compactor_13_38 ,
        masks_for_compactor_13_39 , masks_for_compactor_13_40 , masks_for_compactor_13_41 , masks_for_compactor_13_42 ,
        masks_for_compactor_13_43 , masks_for_compactor_13_44 , masks_for_compactor_13_45 , masks_for_compactor_13_46 ,
        masks_for_compactor_13_47 , masks_for_compactor_13_48 , masks_for_compactor_13_49 , masks_for_compactor_13_50 ,
        masks_for_compactor_13_51 , masks_for_compactor_13_52 , masks_for_compactor_14_0 , masks_for_compactor_14_1 ,
        masks_for_compactor_14_2 , masks_for_compactor_14_3 , masks_for_compactor_14_4 , masks_for_compactor_14_5 ,
        masks_for_compactor_14_6 , masks_for_compactor_14_7 , masks_for_compactor_14_8 , masks_for_compactor_14_9 ,
        masks_for_compactor_14_10 , masks_for_compactor_14_11 , masks_for_compactor_14_12 , masks_for_compactor_14_13 ,
        masks_for_compactor_14_14 , masks_for_compactor_14_15 , masks_for_compactor_14_16 , masks_for_compactor_14_17 ,
        masks_for_compactor_14_18 , masks_for_compactor_14_19 , masks_for_compactor_14_20 , masks_for_compactor_14_21 ,
        masks_for_compactor_14_22 , masks_for_compactor_14_23 , masks_for_compactor_14_24 , masks_for_compactor_14_25 ,
        masks_for_compactor_14_26 , masks_for_compactor_14_27 , masks_for_compactor_14_28 , masks_for_compactor_14_29 ,
        masks_for_compactor_14_30 , masks_for_compactor_14_31 , masks_for_compactor_14_32 , masks_for_compactor_14_33 ,
        masks_for_compactor_14_34 , masks_for_compactor_14_35 , masks_for_compactor_14_36 , masks_for_compactor_14_37 ,
        masks_for_compactor_14_38 , masks_for_compactor_14_39 , masks_for_compactor_14_40 , masks_for_compactor_14_41 ,
        masks_for_compactor_14_42 , masks_for_compactor_14_43 , masks_for_compactor_14_44 , masks_for_compactor_14_45 ,
        masks_for_compactor_14_46 , masks_for_compactor_14_47 , masks_for_compactor_14_48 , masks_for_compactor_14_49 ,
        masks_for_compactor_14_50 , masks_for_compactor_14_51 , masks_for_compactor_14_52 , edt_scan_in_0 ,
        edt_scan_in_1 , edt_scan_in_2 , edt_scan_in_3 , edt_scan_in_4 ,
        edt_scan_in_5 , edt_scan_in_6 , edt_scan_in_7 , edt_scan_in_8 ,
        edt_scan_in_9 , edt_scan_in_10 , edt_scan_in_11 , edt_scan_in_12 ,
        edt_scan_in_13 , edt_scan_in_14 , edt_scan_in_15 , edt_scan_in_16 ,
        edt_scan_in_17 , edt_scan_in_18 , edt_scan_in_19 , edt_scan_in_20 ,
        edt_scan_in_21 , edt_scan_in_22 , edt_scan_in_23 , edt_scan_in_24 ,
        edt_scan_in_25 , edt_scan_in_26 , edt_scan_in_27 , edt_scan_in_28 ,
        edt_scan_in_29 , edt_scan_in_30 , edt_scan_in_31 , edt_scan_in_32 ,
        edt_scan_in_33 , edt_scan_in_34 , edt_scan_in_35 , edt_scan_in_36 ,
        edt_scan_in_37 , edt_scan_in_38 , edt_scan_in_39 , edt_scan_in_40 ,
        edt_scan_in_41 , edt_scan_in_42 , edt_scan_in_43 , edt_scan_in_44 ,
        edt_scan_in_45 , edt_scan_in_46 , edt_scan_in_47 , edt_scan_in_48 ,
        edt_scan_in_49 , edt_scan_in_50 , edt_scan_in_51 , edt_scan_in_52 ,
        edt_scan_in_53 , edt_scan_in_54 , edt_scan_in_55 , edt_scan_in_56 ,
        edt_scan_in_57 , edt_scan_in_58 , edt_scan_in_59 , edt_scan_in_60 ,
        edt_scan_in_61 , edt_scan_in_62 , edt_scan_in_63 , edt_scan_in_64 ,
        edt_scan_in_65 , edt_scan_in_66 , edt_scan_in_67 , edt_scan_in_68 ,
        edt_scan_in_69 , edt_scan_in_70 , edt_scan_in_71 , edt_scan_in_72 ,
        edt_scan_in_73 , edt_scan_in_74 , edt_scan_in_75 , edt_scan_in_76 ,
        edt_scan_in_77 , edt_scan_in_78 , edt_scan_in_79 , edt_scan_in_80 ,
        edt_scan_in_81 , edt_scan_in_82 , edt_scan_in_83 , edt_scan_in_84 ,
        edt_scan_in_85 , edt_scan_in_86 , edt_scan_in_87 , edt_scan_in_88 ,
        edt_scan_in_89 , edt_scan_in_90 , edt_scan_in_91 , edt_scan_in_92 ,
        edt_scan_in_93 , edt_scan_in_94 , edt_scan_in_95 , edt_scan_in_96 ,
        edt_scan_in_97 , edt_scan_in_98 , edt_scan_in_99 , edt_scan_in_100 ,
        edt_scan_in_101 , edt_scan_in_102 , edt_scan_in_103 , edt_scan_in_104 ,
        edt_scan_in_105 , edt_scan_in_106 , edt_scan_in_107 , edt_scan_in_108 ,
        edt_scan_in_109 , edt_scan_in_110 , edt_scan_in_111 , edt_scan_in_112 ,
        edt_scan_in_113 , edt_scan_in_114 , edt_scan_in_115 , edt_scan_in_116 ,
        edt_scan_in_117 , edt_scan_in_118 , edt_scan_in_119 , edt_scan_in_120 ,
        edt_scan_in_121 , edt_scan_in_122 , edt_scan_in_123 , edt_scan_in_124 ,
        edt_scan_in_125 , edt_scan_in_126 , edt_scan_in_127 , edt_scan_in_128 ,
        edt_scan_in_129 , edt_scan_in_130 , edt_scan_in_131 , edt_scan_in_132 ,
        edt_scan_in_133 , edt_scan_in_134 , edt_scan_in_135 , edt_scan_in_136 ,
        edt_scan_in_137 , edt_scan_in_138 , edt_scan_in_139 , edt_scan_in_140 ,
        edt_scan_in_141 , edt_scan_in_142 , edt_scan_in_143 , edt_scan_in_144 ,
        edt_scan_in_145 , edt_scan_in_146 , edt_scan_in_147 , edt_scan_in_148 ,
        edt_scan_in_149 , edt_scan_in_150 , edt_scan_in_151 , edt_scan_in_152 ,
        edt_scan_in_153 , edt_scan_in_154 , edt_scan_in_155 , edt_scan_in_156 ,
        edt_scan_in_157 , edt_scan_in_158 , edt_scan_in_159 , edt_scan_in_160 ,
        edt_scan_in_161 , edt_scan_in_162 , edt_scan_in_163 , edt_scan_in_164 ,
        edt_scan_in_165 , edt_scan_in_166 , edt_scan_in_167 , edt_scan_in_168 ,
        edt_scan_in_169 , edt_scan_in_170 , edt_scan_in_171 , edt_scan_in_172 ,
        edt_scan_in_173 , edt_scan_in_174 , edt_scan_in_175 , edt_scan_in_176 ,
        edt_scan_in_177 , edt_scan_in_178 , edt_scan_in_179 , edt_scan_in_180 ,
        edt_scan_in_181 , edt_scan_in_182 , edt_scan_in_183 , edt_scan_in_184 ,
        edt_scan_in_185 , edt_scan_in_186 , edt_scan_in_187 , edt_scan_in_188 ,
        edt_scan_in_189 , edt_scan_in_190 , edt_scan_in_191 , edt_scan_in_192 ,
        edt_scan_in_193 , edt_scan_in_194 , edt_scan_in_195 , edt_scan_in_196 ,
        edt_scan_in_197 , edt_scan_in_198 , edt_scan_in_199 , edt_scan_in_200 ,
        edt_scan_in_201 , edt_scan_in_202 , edt_scan_in_203 , edt_scan_in_204 ,
        edt_scan_in_205 , edt_scan_in_206 , edt_scan_in_207 , edt_scan_in_208 ,
        edt_scan_in_209 , edt_scan_in_210 , edt_scan_in_211 , edt_scan_in_212 ,
        edt_scan_in_213 , edt_scan_in_214 , edt_scan_in_215 , edt_scan_in_216 ,
        edt_scan_in_217 , edt_scan_in_218 , edt_scan_in_219 , edt_scan_in_220 ,
        edt_scan_in_221 , edt_scan_in_222 , edt_scan_in_223 , edt_scan_in_224 ,
        edt_scan_in_225 , edt_scan_in_226 , edt_scan_in_227 , edt_scan_in_228 ,
        edt_scan_in_229 , edt_scan_in_230 , edt_scan_in_231 , edt_scan_in_232 ,
        edt_scan_in_233 , edt_scan_in_234 , edt_scan_in_235 , edt_scan_in_236 ,
        edt_scan_in_237 , edt_scan_in_238 , edt_scan_in_239 , edt_scan_in_240 ,
        edt_scan_in_241 , edt_scan_in_242 , edt_scan_in_243 , edt_scan_in_244 ,
        edt_scan_in_245 , edt_scan_in_246 , edt_scan_in_247 , edt_scan_in_248 ,
        edt_scan_in_249 , edt_scan_in_250 , edt_scan_in_251 , edt_scan_in_252 ,
        edt_scan_in_253 , edt_scan_in_254 , edt_scan_in_255 , edt_scan_in_256 ,
        edt_scan_in_257 , edt_scan_in_258 , edt_scan_in_259 , edt_scan_in_260 ,
        edt_scan_in_261 , edt_scan_in_262 , edt_scan_in_263 , edt_scan_in_264 ,
        edt_scan_in_265 , edt_scan_in_266 , edt_scan_in_267 , edt_scan_in_268 ,
        edt_scan_in_269 , edt_scan_in_270 , edt_scan_in_271 , edt_scan_in_272 ,
        edt_scan_in_273 , edt_scan_in_274 , edt_scan_in_275 , edt_scan_in_276 ,
        edt_scan_in_277 , edt_scan_in_278 , edt_scan_in_279 , edt_scan_in_280 ,
        edt_scan_in_281 , edt_scan_in_282 , edt_scan_in_283 , edt_scan_in_284 ,
        edt_scan_in_285 , edt_scan_in_286 , edt_scan_in_287 , edt_scan_in_288 ,
        edt_scan_in_289 , edt_scan_in_290 , edt_scan_in_291 , edt_scan_in_292 ,
        edt_scan_in_293 , edt_scan_in_294 , edt_scan_in_295 , edt_scan_in_296 ,
        edt_scan_in_297 , edt_scan_in_298 , edt_scan_in_299 , edt_scan_in_300 ,
        edt_scan_in_301 , edt_scan_in_302 , edt_scan_in_303 , edt_scan_in_304 ,
        edt_scan_in_305 , edt_scan_in_306 , edt_scan_in_307 , edt_scan_in_308 ,
        edt_scan_in_309 , edt_scan_in_310 , edt_scan_in_311 , edt_scan_in_312 ,
        edt_scan_in_313 , edt_scan_in_314 , edt_scan_in_315 , edt_scan_in_316 ,
        edt_scan_in_317 , edt_scan_in_318 , edt_scan_in_319 , edt_scan_in_320 ,
        edt_scan_in_321 , edt_scan_in_322 , edt_scan_in_323 , edt_scan_in_324 ,
        edt_scan_in_325 , edt_scan_in_326 , edt_scan_in_327 , edt_scan_in_328 ,
        edt_scan_in_329 , edt_scan_in_330 , edt_scan_in_331 , edt_scan_in_332 ,
        edt_scan_in_333 , edt_scan_in_334 , edt_scan_in_335 , edt_scan_in_336 ,
        edt_scan_in_337 , edt_scan_in_338 , edt_scan_in_339 , edt_scan_in_340 ,
        edt_scan_in_341 , edt_scan_in_342 , edt_scan_in_343 , edt_scan_in_344 ,
        edt_scan_in_345 , edt_scan_in_346 , edt_scan_in_347 , edt_scan_in_348 ,
        edt_scan_in_349 , edt_scan_in_350 , edt_scan_in_351 , edt_scan_in_352 ,
        edt_scan_in_353 , edt_scan_in_354 , edt_scan_in_355 , edt_scan_in_356 ,
        edt_scan_in_357 , edt_scan_in_358 , edt_scan_in_359 , edt_scan_in_360 ,
        edt_scan_in_361 , edt_scan_in_362 , edt_scan_in_363 , edt_scan_in_364 ,
        edt_scan_in_365 , edt_scan_in_366 , edt_scan_in_367 , edt_scan_in_368 ,
        edt_scan_in_369 , edt_scan_in_370 , edt_scan_in_371 , edt_scan_in_372 ,
        edt_scan_in_373 , edt_scan_in_374 , edt_scan_in_375 , edt_scan_in_376 ,
        edt_scan_in_377 , edt_scan_in_378 , edt_scan_in_379 , edt_scan_in_380 ,
        edt_scan_in_381 , edt_scan_in_382 , edt_scan_in_383 , edt_scan_in_384 ,
        edt_scan_in_385 , edt_scan_in_386 , edt_scan_in_387 , edt_scan_in_388 ,
        edt_scan_in_389 , edt_scan_in_390 , edt_scan_in_391 , edt_scan_in_392 ,
        edt_scan_in_393 , edt_scan_in_394 , edt_scan_in_395 , edt_scan_in_396 ,
        edt_scan_in_397 , edt_scan_in_398 , edt_scan_in_399 , edt_scan_in_400 ,
        edt_scan_in_401 , edt_scan_in_402 , edt_scan_in_403 , edt_scan_in_404 ,
        edt_scan_in_405 , edt_scan_in_406 , edt_scan_in_407 , edt_scan_in_408 ,
        edt_scan_in_409 , edt_scan_in_410 , edt_scan_in_411 , edt_scan_in_412 ,
        edt_scan_in_413 , edt_scan_in_414 , edt_scan_in_415 , edt_scan_in_416 ,
        edt_scan_in_417 , edt_scan_in_418 , edt_scan_in_419 , edt_scan_in_420 ,
        edt_scan_in_421 , edt_scan_in_422 , edt_scan_in_423 , edt_scan_in_424 ,
        edt_scan_in_425 , edt_scan_in_426 , edt_scan_in_427 , edt_scan_in_428 ,
        edt_scan_in_429 , edt_scan_in_430 , edt_scan_in_431 , edt_scan_in_432 ,
        edt_scan_in_433 , edt_scan_in_434 , edt_scan_in_435 , edt_scan_in_436 ,
        edt_scan_in_437 , edt_scan_in_438 , edt_scan_in_439 , edt_scan_in_440 ,
        edt_scan_in_441 , edt_scan_in_442 , edt_scan_in_443 , edt_scan_in_444 ,
        edt_scan_in_445 , edt_scan_in_446 , edt_scan_in_447 , edt_scan_in_448 ,
        edt_scan_in_449 , edt_scan_in_450 , edt_scan_in_451 , edt_scan_in_452 ,
        edt_scan_in_453 , edt_scan_in_454 , edt_scan_in_455 , edt_scan_in_456 ,
        edt_scan_in_457 , edt_scan_in_458 , edt_scan_in_459 , edt_scan_in_460 ,
        edt_scan_in_461 , edt_scan_in_462 , edt_scan_in_463 , edt_scan_in_464 ,
        edt_scan_in_465 , edt_scan_in_466 , edt_scan_in_467 , edt_scan_in_468 ,
        edt_scan_in_469 , edt_scan_in_470 , edt_scan_in_471 , edt_scan_in_472 ,
        edt_scan_in_473 , edt_scan_in_474 , edt_scan_in_475 , edt_scan_in_476 ,
        edt_scan_in_477 , edt_scan_in_478 , edt_scan_in_479 , edt_scan_in_480 ,
        edt_scan_in_481 , edt_scan_in_482 , edt_scan_in_483 , edt_scan_in_484 ,
        edt_scan_in_485 , edt_scan_in_486 , edt_scan_in_487 , edt_scan_in_488 ,
        edt_scan_in_489 , edt_scan_in_490 , edt_scan_in_491 , edt_scan_in_492 ,
        edt_scan_in_493 , edt_scan_in_494 , edt_scan_in_495 , edt_scan_in_496 ,
        edt_scan_in_497 , edt_scan_in_498 , edt_scan_in_499 , edt_scan_in_500 ,
        edt_scan_in_501 , edt_scan_in_502 , edt_scan_in_503 , edt_scan_in_504 ,
        edt_scan_in_505 , edt_scan_in_506 , edt_scan_in_507 , edt_scan_in_508 ,
        edt_scan_in_509 , edt_scan_in_510 , edt_scan_in_511 , edt_scan_in_512 ,
        edt_scan_in_513 , edt_scan_in_514 , edt_scan_in_515 , edt_scan_in_516 ,
        edt_scan_in_517 , edt_scan_in_518 , edt_scan_in_519 , edt_scan_in_520 ,
        edt_scan_in_521 , edt_scan_in_522 , edt_scan_in_523 , edt_scan_in_524 ,
        edt_scan_in_525 , edt_scan_in_526 , edt_scan_in_527 , edt_scan_in_528 ,
        edt_scan_in_529 , edt_scan_in_530 , edt_scan_in_531 , edt_scan_in_532 ,
        edt_scan_in_533 , edt_scan_in_534 , edt_scan_in_535 , edt_scan_in_536 ,
        edt_scan_in_537 , edt_scan_in_538 , edt_scan_in_539 , edt_scan_in_540 ,
        edt_scan_in_541 , edt_scan_in_542 , edt_scan_in_543 , edt_scan_in_544 ,
        edt_scan_in_545 , edt_scan_in_546 , edt_scan_in_547 , edt_scan_in_548 ,
        edt_scan_in_549 , edt_scan_in_550 , edt_scan_in_551 , edt_scan_in_552 ,
        edt_scan_in_553 , edt_scan_in_554 , edt_scan_in_555 , edt_scan_in_556 ,
        edt_scan_in_557 , edt_scan_in_558 , edt_scan_in_559 , edt_scan_in_560 ,
        edt_scan_in_561 , edt_scan_in_562 , edt_scan_in_563 , edt_scan_in_564 ,
        edt_scan_in_565 , edt_scan_in_566 , edt_scan_in_567 , edt_scan_in_568 ,
        edt_scan_in_569 , edt_scan_in_570 , edt_scan_in_571 , edt_scan_in_572 ,
        edt_scan_in_573 , edt_scan_in_574 , edt_scan_in_575 , edt_scan_in_576 ,
        edt_scan_in_577 , edt_scan_in_578 , edt_scan_in_579 , edt_scan_in_580 ,
        edt_scan_in_581 , edt_scan_in_582 , edt_scan_in_583 , edt_scan_in_584 ,
        edt_scan_in_585 , edt_scan_in_586 , edt_scan_in_587 , edt_scan_in_588 ,
        edt_scan_in_589 , edt_scan_in_590 , edt_scan_in_591 , edt_scan_in_592 ,
        edt_scan_in_593 , edt_scan_in_594 , edt_scan_in_595 , edt_scan_in_596 ,
        edt_scan_in_597 , edt_scan_in_598 , edt_scan_in_599 , edt_scan_in_600 ,
        edt_scan_in_601 , edt_scan_in_602 , edt_scan_in_603 , edt_scan_in_604 ,
        edt_scan_in_605 , edt_scan_in_606 , edt_scan_in_607 , edt_scan_in_608 ,
        edt_scan_in_609 , edt_scan_in_610 , edt_scan_in_611 , edt_scan_in_612 ,
        edt_scan_in_613 , edt_scan_in_614 , edt_scan_in_615 , edt_scan_in_616 ,
        edt_scan_in_617 , edt_scan_in_618 , edt_scan_in_619 , edt_scan_in_620 ,
        edt_scan_in_621 , edt_scan_in_622 , edt_scan_in_623 , edt_scan_in_624 ,
        edt_scan_in_625 , edt_scan_in_626 , edt_scan_in_627 , edt_scan_in_628 ,
        edt_scan_in_629 , edt_scan_in_630 , edt_scan_in_631 , edt_scan_in_632 ,
        edt_scan_in_633 , edt_scan_in_634 , edt_scan_in_635 , edt_scan_in_636 ,
        edt_scan_in_637 , edt_scan_in_638 , edt_scan_in_639 , edt_scan_in_640 ,
        edt_scan_in_641 , edt_scan_in_642 , edt_scan_in_643 , edt_scan_in_644 ,
        edt_scan_in_645 , edt_scan_in_646 , edt_scan_in_647 , edt_scan_in_648 ,
        edt_scan_in_649 , edt_scan_in_650 , edt_scan_in_651 , edt_scan_in_652 ,
        edt_scan_in_653 , edt_scan_in_654 , edt_scan_in_655 , edt_scan_in_656 ,
        edt_scan_in_657 , edt_scan_in_658 , edt_scan_in_659 , edt_scan_in_660 ,
        edt_scan_in_661 , edt_scan_in_662 , edt_scan_in_663 , edt_scan_in_664 ,
        edt_scan_in_665 , edt_scan_in_666 , edt_scan_in_667 , edt_scan_in_668 ,
        edt_scan_in_669 , edt_scan_in_670 , edt_scan_in_671 , edt_scan_in_672 ,
        edt_scan_in_673 , edt_scan_in_674 , edt_scan_in_675 , edt_scan_in_676 ,
        edt_scan_in_677 , edt_scan_in_678 , edt_scan_in_679 , edt_scan_in_680 ,
        edt_scan_in_681 , edt_scan_in_682 , edt_scan_in_683 , edt_scan_in_684 ,
        edt_scan_in_685 , edt_scan_in_686 , edt_scan_in_687 , edt_scan_in_688 ,
        edt_scan_in_689 , edt_scan_in_690 , edt_scan_in_691 , edt_scan_in_692 ,
        edt_scan_in_693 , edt_scan_in_694 , edt_scan_in_695 , edt_scan_in_696 ,
        edt_scan_in_697 , edt_scan_in_698 , edt_scan_in_699 , edt_scan_in_700 ,
        edt_scan_in_701 , edt_scan_in_702 , edt_scan_in_703 , edt_scan_in_704 ,
        edt_scan_in_705 , edt_scan_in_706 , edt_scan_in_707 , edt_scan_in_708 ,
        edt_scan_in_709 , edt_scan_in_710 , edt_scan_in_711 , edt_scan_in_712 ,
        edt_scan_in_713 , edt_scan_in_714 , edt_scan_in_715 , edt_scan_in_716 ,
        edt_scan_in_717 , edt_scan_in_718 , edt_scan_in_719 , edt_scan_in_720 ,
        edt_scan_in_721 , edt_scan_in_722 , edt_scan_in_723 , edt_scan_in_724 ,
        edt_scan_in_725 , edt_scan_in_726 , edt_scan_in_727 , edt_scan_in_728 ,
        edt_scan_in_729 , edt_scan_in_730 , edt_scan_in_731 , edt_scan_in_732 ,
        edt_scan_in_733 , edt_scan_in_734 , edt_scan_in_735 , edt_scan_in_736 ,
        edt_scan_in_737 , edt_scan_in_738 , edt_scan_in_739 , edt_scan_in_740 ,
        edt_scan_in_741 , edt_scan_in_742 , edt_scan_in_743 , edt_scan_in_744 ,
        edt_scan_in_745 , edt_scan_in_746 , edt_scan_in_747 , edt_scan_in_748 ,
        edt_scan_in_749 , edt_scan_in_750 , edt_scan_in_751 , edt_scan_in_752 ,
        edt_scan_in_753 , edt_scan_in_754 , edt_scan_in_755 , edt_scan_in_756 ,
        edt_scan_in_757 , edt_scan_in_758 , edt_scan_in_759 , edt_scan_in_760 ,
        edt_scan_in_761 , edt_scan_in_762 , edt_scan_in_763 , edt_scan_in_764 ,
        edt_scan_in_765 , edt_scan_in_766 , edt_scan_in_767 , edt_scan_in_768 ,
        edt_scan_in_769 , edt_scan_in_770 , edt_scan_in_771 , edt_scan_in_772 ,
        edt_scan_in_773 , edt_scan_in_774 , edt_scan_in_775 , edt_scan_in_776 ,
        edt_scan_in_777 , edt_scan_in_778 , edt_scan_in_779 , edt_scan_in_780 ,
        edt_scan_in_781 , edt_scan_in_782 , edt_scan_in_783 , edt_scan_in_784 ,
        edt_scan_in_785 , edt_scan_in_786 , edt_scan_in_787 , edt_scan_in_788 ,
        edt_scan_in_789 , edt_scan_in_790 , edt_scan_in_791 , edt_scan_in_792 ,
        edt_scan_in_793 , edt_scan_in_794 , edt_scan_in_795 , edt_channels_in_0 ,
        edt_channels_in_1 , edt_channels_in_2 , edt_channels_in_3 , edt_channels_in_4 ,
        edt_channels_in_5 , edt_channels_in_6 , edt_channels_in_7 , edt_channels_in_8 ,
        edt_channels_in_9 , edt_channels_in_10 , edt_channels_in_11 , edt_channels_in_12 ,
        edt_channels_in_13 , edt_channels_in_14 , edt_clock , edt_update ,
        edt_configuration , edt_shift_const_en , edt_decompressor_out_0 , edt_decompressor_out_1 ,
        edt_decompressor_out_2 , edt_decompressor_out_3 , edt_decompressor_out_4 , edt_decompressor_out_5 ,
        edt_decompressor_out_6 , edt_decompressor_out_7 , edt_decompressor_out_8 , edt_decompressor_out_9 ,
        edt_decompressor_out_10 , edt_decompressor_out_11 , edt_decompressor_out_12 , edt_decompressor_out_13 ,
        edt_decompressor_out_14 , edt_decompressor_out_15 , edt_decompressor_out_16 , edt_decompressor_out_17 ,
        edt_decompressor_out_18 , edt_decompressor_out_19 , edt_decompressor_out_20 , edt_decompressor_out_21 ,
        edt_decompressor_out_22 , edt_decompressor_out_23 , edt_decompressor_out_24 , edt_decompressor_out_25 ,
        edt_decompressor_out_26 , edt_decompressor_out_27 , edt_decompressor_out_28 , edt_decompressor_out_29 ,
        edt_decompressor_out_30 , edt_decompressor_out_31 , edt_decompressor_out_32 , edt_decompressor_out_33 ,
        edt_decompressor_out_34 , edt_decompressor_out_35 , edt_decompressor_out_36 , edt_decompressor_out_37 ,
        edt_decompressor_out_38 , edt_decompressor_out_39 , edt_decompressor_out_40 , edt_decompressor_out_41 ,
        edt_decompressor_out_42 , edt_decompressor_out_43 , edt_decompressor_out_44 , edt_decompressor_out_45 ,
        edt_decompressor_out_46 , edt_decompressor_out_47 , edt_decompressor_out_48 , edt_decompressor_out_49 ,
        edt_decompressor_out_50 , edt_decompressor_out_51 , edt_decompressor_out_52 , edt_decompressor_out_53 ,
        edt_decompressor_out_54 , edt_decompressor_out_55 , edt_decompressor_out_56 , edt_decompressor_out_57 ,
        edt_decompressor_out_58 , edt_decompressor_out_59 , edt_decompressor_out_60 , edt_decompressor_out_61 ,
        edt_decompressor_out_62 , edt_decompressor_out_63 , edt_decompressor_out_64 , edt_decompressor_out_65 ,
        edt_decompressor_out_66 , edt_decompressor_out_67 , edt_decompressor_out_68 , edt_decompressor_out_69 ,
        edt_decompressor_out_70 , edt_decompressor_out_71 , edt_decompressor_out_72 , edt_decompressor_out_73 ,
        edt_decompressor_out_74 , edt_decompressor_out_75 , edt_decompressor_out_76 , edt_decompressor_out_77 ,
        edt_decompressor_out_78 , edt_decompressor_out_79 , edt_decompressor_out_80 , edt_decompressor_out_81 ,
        edt_decompressor_out_82 , edt_decompressor_out_83 , edt_decompressor_out_84 , edt_decompressor_out_85 ,
        edt_decompressor_out_86 , edt_decompressor_out_87 , edt_decompressor_out_88 , edt_decompressor_out_89 ,
        edt_decompressor_out_90 , edt_decompressor_out_91 , edt_decompressor_out_92 , edt_decompressor_out_93 ,
        edt_decompressor_out_94 , edt_decompressor_out_95 , edt_decompressor_out_96 , edt_decompressor_out_97 ,
        edt_decompressor_out_98 , edt_decompressor_out_99 , edt_decompressor_out_100 , edt_decompressor_out_101 ,
        edt_decompressor_out_102 , edt_decompressor_out_103 , edt_decompressor_out_104 , edt_decompressor_out_105 ,
        edt_decompressor_out_106 , edt_decompressor_out_107 , edt_decompressor_out_108 , edt_decompressor_out_109 ,
        edt_decompressor_out_110 , edt_decompressor_out_111 , edt_decompressor_out_112 , edt_decompressor_out_113 ,
        edt_decompressor_out_114 , edt_decompressor_out_115 , edt_decompressor_out_116 , edt_decompressor_out_117 ,
        edt_decompressor_out_118 , edt_decompressor_out_119 , edt_decompressor_out_120 , edt_decompressor_out_121 ,
        edt_decompressor_out_122 , edt_decompressor_out_123 , edt_decompressor_out_124 , edt_decompressor_out_125 ,
        edt_decompressor_out_126 , edt_decompressor_out_127 , edt_decompressor_out_128 , edt_decompressor_out_129 ,
        edt_decompressor_out_130 , edt_decompressor_out_131 , edt_decompressor_out_132 , edt_decompressor_out_133 ,
        edt_decompressor_out_134 , edt_decompressor_out_135 , edt_decompressor_out_136 , edt_decompressor_out_137 ,
        edt_decompressor_out_138 , edt_decompressor_out_139 , edt_decompressor_out_140 , edt_decompressor_out_141 ,
        edt_decompressor_out_142 , edt_decompressor_out_143 , edt_decompressor_out_144 , edt_decompressor_out_145 ,
        edt_decompressor_out_146 , edt_decompressor_out_147 , edt_decompressor_out_148 , edt_decompressor_out_149 ,
        edt_decompressor_out_150 , edt_decompressor_out_151 , edt_decompressor_out_152 , edt_decompressor_out_153 ,
        edt_decompressor_out_154 , edt_decompressor_out_155 , edt_decompressor_out_156 , edt_decompressor_out_157 ,
        edt_decompressor_out_158 , edt_decompressor_out_159 , edt_decompressor_out_160 , edt_decompressor_out_161 ,
        edt_decompressor_out_162 , edt_decompressor_out_163 , edt_decompressor_out_164 , edt_decompressor_out_165 ,
        edt_decompressor_out_166 , edt_decompressor_out_167 , edt_decompressor_out_168 , edt_decompressor_out_169 ,
        edt_decompressor_out_170 , edt_decompressor_out_171 , edt_decompressor_out_172 , edt_decompressor_out_173 ,
        edt_decompressor_out_174 , edt_decompressor_out_175 , edt_decompressor_out_176 , edt_decompressor_out_177 ,
        edt_decompressor_out_178 , edt_decompressor_out_179 , edt_decompressor_out_180 , edt_decompressor_out_181 ,
        edt_decompressor_out_182 , edt_decompressor_out_183 , edt_decompressor_out_184 , edt_decompressor_out_185 ,
        edt_decompressor_out_186 , edt_decompressor_out_187 , edt_decompressor_out_188 , edt_decompressor_out_189 ,
        edt_decompressor_out_190 , edt_decompressor_out_191 , edt_decompressor_out_192 , edt_decompressor_out_193 ,
        edt_decompressor_out_194 , edt_decompressor_out_195 , edt_decompressor_out_196 , edt_decompressor_out_197 ,
        edt_decompressor_out_198 , edt_decompressor_out_199 , edt_decompressor_out_200 , edt_decompressor_out_201 ,
        edt_decompressor_out_202 , edt_decompressor_out_203 , edt_decompressor_out_204 , edt_decompressor_out_205 ,
        edt_decompressor_out_206 , edt_decompressor_out_207 , edt_decompressor_out_208 , edt_decompressor_out_209 ,
        edt_decompressor_out_210 , edt_decompressor_out_211 , edt_decompressor_out_212 , edt_decompressor_out_213 ,
        edt_decompressor_out_214 , edt_decompressor_out_215 , edt_decompressor_out_216 , edt_decompressor_out_217 ,
        edt_decompressor_out_218 , edt_decompressor_out_219 , edt_decompressor_out_220 , edt_decompressor_out_221 ,
        edt_decompressor_out_222 , edt_decompressor_out_223 , edt_decompressor_out_224 , edt_decompressor_out_225 ,
        edt_decompressor_out_226 , edt_decompressor_out_227 , edt_decompressor_out_228 , edt_decompressor_out_229 ,
        edt_decompressor_out_230 , edt_decompressor_out_231 , edt_decompressor_out_232 , edt_decompressor_out_233 ,
        edt_decompressor_out_234 , edt_decompressor_out_235 , edt_decompressor_out_236 , edt_decompressor_out_237 ,
        edt_decompressor_out_238 , edt_decompressor_out_239 , edt_decompressor_out_240 , edt_decompressor_out_241 ,
        edt_decompressor_out_242 , edt_decompressor_out_243 , edt_decompressor_out_244 , edt_decompressor_out_245 ,
        edt_decompressor_out_246 , edt_decompressor_out_247 , edt_decompressor_out_248 , edt_decompressor_out_249 ,
        edt_decompressor_out_250 , edt_decompressor_out_251 , edt_decompressor_out_252 , edt_decompressor_out_253 ,
        edt_decompressor_out_254 , edt_decompressor_out_255 , edt_decompressor_out_256 , edt_decompressor_out_257 ,
        edt_decompressor_out_258 , edt_decompressor_out_259 , edt_decompressor_out_260 , edt_decompressor_out_261 ,
        edt_decompressor_out_262 , edt_decompressor_out_263 , edt_decompressor_out_264 , edt_decompressor_out_265 ,
        edt_decompressor_out_266 , edt_decompressor_out_267 , edt_decompressor_out_268 , edt_decompressor_out_269 ,
        edt_decompressor_out_270 , edt_decompressor_out_271 , edt_decompressor_out_272 , edt_decompressor_out_273 ,
        edt_decompressor_out_274 , edt_decompressor_out_275 , edt_decompressor_out_276 , edt_decompressor_out_277 ,
        edt_decompressor_out_278 , edt_decompressor_out_279 , edt_decompressor_out_280 , edt_decompressor_out_281 ,
        edt_decompressor_out_282 , edt_decompressor_out_283 , edt_decompressor_out_284 , edt_decompressor_out_285 ,
        edt_decompressor_out_286 , edt_decompressor_out_287 , edt_decompressor_out_288 , edt_decompressor_out_289 ,
        edt_decompressor_out_290 , edt_decompressor_out_291 , edt_decompressor_out_292 , edt_decompressor_out_293 ,
        edt_decompressor_out_294 , edt_decompressor_out_295 , edt_decompressor_out_296 , edt_decompressor_out_297 ,
        edt_decompressor_out_298 , edt_decompressor_out_299 , edt_decompressor_out_300 , edt_decompressor_out_301 ,
        edt_decompressor_out_302 , edt_decompressor_out_303 , edt_decompressor_out_304 , edt_decompressor_out_305 ,
        edt_decompressor_out_306 , edt_decompressor_out_307 , edt_decompressor_out_308 , edt_decompressor_out_309 ,
        edt_decompressor_out_310 , edt_decompressor_out_311 , edt_decompressor_out_312 , edt_decompressor_out_313 ,
        edt_decompressor_out_314 , edt_decompressor_out_315 , edt_decompressor_out_316 , edt_decompressor_out_317 ,
        edt_decompressor_out_318 , edt_decompressor_out_319 , edt_decompressor_out_320 , edt_decompressor_out_321 ,
        edt_decompressor_out_322 , edt_decompressor_out_323 , edt_decompressor_out_324 , edt_decompressor_out_325 ,
        edt_decompressor_out_326 , edt_decompressor_out_327 , edt_decompressor_out_328 , edt_decompressor_out_329 ,
        edt_decompressor_out_330 , edt_decompressor_out_331 , edt_decompressor_out_332 , edt_decompressor_out_333 ,
        edt_decompressor_out_334 , edt_decompressor_out_335 , edt_decompressor_out_336 , edt_decompressor_out_337 ,
        edt_decompressor_out_338 , edt_decompressor_out_339 , edt_decompressor_out_340 , edt_decompressor_out_341 ,
        edt_decompressor_out_342 , edt_decompressor_out_343 , edt_decompressor_out_344 , edt_decompressor_out_345 ,
        edt_decompressor_out_346 , edt_decompressor_out_347 , edt_decompressor_out_348 , edt_decompressor_out_349 ,
        edt_decompressor_out_350 , edt_decompressor_out_351 , edt_decompressor_out_352 , edt_decompressor_out_353 ,
        edt_decompressor_out_354 , edt_decompressor_out_355 , edt_decompressor_out_356 , edt_decompressor_out_357 ,
        edt_decompressor_out_358 , edt_decompressor_out_359 , edt_decompressor_out_360 , edt_decompressor_out_361 ,
        edt_decompressor_out_362 , edt_decompressor_out_363 , edt_decompressor_out_364 , edt_decompressor_out_365 ,
        edt_decompressor_out_366 , edt_decompressor_out_367 , edt_decompressor_out_368 , edt_decompressor_out_369 ,
        edt_decompressor_out_370 , edt_decompressor_out_371 , edt_decompressor_out_372 , edt_decompressor_out_373 ,
        edt_decompressor_out_374 , edt_decompressor_out_375 , edt_decompressor_out_376 , edt_decompressor_out_377 ,
        edt_decompressor_out_378 , edt_decompressor_out_379 , edt_decompressor_out_380 , edt_decompressor_out_381 ,
        edt_decompressor_out_382 , edt_decompressor_out_383 , edt_decompressor_out_384 , edt_decompressor_out_385 ,
        edt_decompressor_out_386 , edt_decompressor_out_387 , edt_decompressor_out_388 , edt_decompressor_out_389 ,
        edt_decompressor_out_390 , edt_decompressor_out_391 , edt_decompressor_out_392 , edt_decompressor_out_393 ,
        edt_decompressor_out_394 , edt_decompressor_out_395 , edt_decompressor_out_396 , edt_decompressor_out_397 ,
        edt_decompressor_out_398 , edt_decompressor_out_399 , edt_decompressor_out_400 , edt_decompressor_out_401 ,
        edt_decompressor_out_402 , edt_decompressor_out_403 , edt_decompressor_out_404 , edt_decompressor_out_405 ,
        edt_decompressor_out_406 , edt_decompressor_out_407 , edt_decompressor_out_408 , edt_decompressor_out_409 ,
        edt_decompressor_out_410 , edt_decompressor_out_411 , edt_decompressor_out_412 , edt_decompressor_out_413 ,
        edt_decompressor_out_414 , edt_decompressor_out_415 , edt_decompressor_out_416 , edt_decompressor_out_417 ,
        edt_decompressor_out_418 , edt_decompressor_out_419 , edt_decompressor_out_420 , edt_decompressor_out_421 ,
        edt_decompressor_out_422 , edt_decompressor_out_423 , edt_decompressor_out_424 , edt_decompressor_out_425 ,
        edt_decompressor_out_426 , edt_decompressor_out_427 , edt_decompressor_out_428 , edt_decompressor_out_429 ,
        edt_decompressor_out_430 , edt_decompressor_out_431 , edt_decompressor_out_432 , edt_decompressor_out_433 ,
        edt_decompressor_out_434 , edt_decompressor_out_435 , edt_decompressor_out_436 , edt_decompressor_out_437 ,
        edt_decompressor_out_438 , edt_decompressor_out_439 , edt_decompressor_out_440 , edt_decompressor_out_441 ,
        edt_decompressor_out_442 , edt_decompressor_out_443 , edt_decompressor_out_444 , edt_decompressor_out_445 ,
        edt_decompressor_out_446 , edt_decompressor_out_447 , edt_decompressor_out_448 , edt_decompressor_out_449 ,
        edt_decompressor_out_450 , edt_decompressor_out_451 , edt_decompressor_out_452 , edt_decompressor_out_453 ,
        edt_decompressor_out_454 , edt_decompressor_out_455 , edt_decompressor_out_456 , edt_decompressor_out_457 ,
        edt_decompressor_out_458 , edt_decompressor_out_459 , edt_decompressor_out_460 , edt_decompressor_out_461 ,
        edt_decompressor_out_462 , edt_decompressor_out_463 , edt_decompressor_out_464 , edt_decompressor_out_465 ,
        edt_decompressor_out_466 , edt_decompressor_out_467 , edt_decompressor_out_468 , edt_decompressor_out_469 ,
        edt_decompressor_out_470 , edt_decompressor_out_471 , edt_decompressor_out_472 , edt_decompressor_out_473 ,
        edt_decompressor_out_474 , edt_decompressor_out_475 , edt_decompressor_out_476 , edt_decompressor_out_477 ,
        edt_decompressor_out_478 , edt_decompressor_out_479 , edt_decompressor_out_480 , edt_decompressor_out_481 ,
        edt_decompressor_out_482 , edt_decompressor_out_483 , edt_decompressor_out_484 , edt_decompressor_out_485 ,
        edt_decompressor_out_486 , edt_decompressor_out_487 , edt_decompressor_out_488 , edt_decompressor_out_489 ,
        edt_decompressor_out_490 , edt_decompressor_out_491 , edt_decompressor_out_492 , edt_decompressor_out_493 ,
        edt_decompressor_out_494 , edt_decompressor_out_495 , edt_decompressor_out_496 , edt_decompressor_out_497 ,
        edt_decompressor_out_498 , edt_decompressor_out_499 , edt_decompressor_out_500 , edt_decompressor_out_501 ,
        edt_decompressor_out_502 , edt_decompressor_out_503 , edt_decompressor_out_504 , edt_decompressor_out_505 ,
        edt_decompressor_out_506 , edt_decompressor_out_507 , edt_decompressor_out_508 , edt_decompressor_out_509 ,
        edt_decompressor_out_510 , edt_decompressor_out_511 , edt_decompressor_out_512 , edt_decompressor_out_513 ,
        edt_decompressor_out_514 , edt_decompressor_out_515 , edt_decompressor_out_516 , edt_decompressor_out_517 ,
        edt_decompressor_out_518 , edt_decompressor_out_519 , edt_decompressor_out_520 , edt_decompressor_out_521 ,
        edt_decompressor_out_522 , edt_decompressor_out_523 , edt_decompressor_out_524 , edt_decompressor_out_525 ,
        edt_decompressor_out_526 , edt_decompressor_out_527 , edt_decompressor_out_528 , edt_decompressor_out_529 ,
        edt_decompressor_out_530 , edt_decompressor_out_531 , edt_decompressor_out_532 , edt_decompressor_out_533 ,
        edt_decompressor_out_534 , edt_decompressor_out_535 , edt_decompressor_out_536 , edt_decompressor_out_537 ,
        edt_decompressor_out_538 , edt_decompressor_out_539 , edt_decompressor_out_540 , edt_decompressor_out_541 ,
        edt_decompressor_out_542 , edt_decompressor_out_543 , edt_decompressor_out_544 , edt_decompressor_out_545 ,
        edt_decompressor_out_546 , edt_decompressor_out_547 , edt_decompressor_out_548 , edt_decompressor_out_549 ,
        edt_decompressor_out_550 , edt_decompressor_out_551 , edt_decompressor_out_552 , edt_decompressor_out_553 ,
        edt_decompressor_out_554 , edt_decompressor_out_555 , edt_decompressor_out_556 , edt_decompressor_out_557 ,
        edt_decompressor_out_558 , edt_decompressor_out_559 , edt_decompressor_out_560 , edt_decompressor_out_561 ,
        edt_decompressor_out_562 , edt_decompressor_out_563 , edt_decompressor_out_564 , edt_decompressor_out_565 ,
        edt_decompressor_out_566 , edt_decompressor_out_567 , edt_decompressor_out_568 , edt_decompressor_out_569 ,
        edt_decompressor_out_570 , edt_decompressor_out_571 , edt_decompressor_out_572 , edt_decompressor_out_573 ,
        edt_decompressor_out_574 , edt_decompressor_out_575 , edt_decompressor_out_576 , edt_decompressor_out_577 ,
        edt_decompressor_out_578 , edt_decompressor_out_579 , edt_decompressor_out_580 , edt_decompressor_out_581 ,
        edt_decompressor_out_582 , edt_decompressor_out_583 , edt_decompressor_out_584 , edt_decompressor_out_585 ,
        edt_decompressor_out_586 , edt_decompressor_out_587 , edt_decompressor_out_588 , edt_decompressor_out_589 ,
        edt_decompressor_out_590 , edt_decompressor_out_591 , edt_decompressor_out_592 , edt_decompressor_out_593 ,
        edt_decompressor_out_594 , edt_decompressor_out_595 , edt_decompressor_out_596 , edt_decompressor_out_597 ,
        edt_decompressor_out_598 , edt_decompressor_out_599 , edt_decompressor_out_600 , edt_decompressor_out_601 ,
        edt_decompressor_out_602 , edt_decompressor_out_603 , edt_decompressor_out_604 , edt_decompressor_out_605 ,
        edt_decompressor_out_606 , edt_decompressor_out_607 , edt_decompressor_out_608 , edt_decompressor_out_609 ,
        edt_decompressor_out_610 , edt_decompressor_out_611 , edt_decompressor_out_612 , edt_decompressor_out_613 ,
        edt_decompressor_out_614 , edt_decompressor_out_615 , edt_decompressor_out_616 , edt_decompressor_out_617 ,
        edt_decompressor_out_618 , edt_decompressor_out_619 , edt_decompressor_out_620 , edt_decompressor_out_621 ,
        edt_decompressor_out_622 , edt_decompressor_out_623 , edt_decompressor_out_624 , edt_decompressor_out_625 ,
        edt_decompressor_out_626 , edt_decompressor_out_627 , edt_decompressor_out_628 , edt_decompressor_out_629 ,
        edt_decompressor_out_630 , edt_decompressor_out_631 , edt_decompressor_out_632 , edt_decompressor_out_633 ,
        edt_decompressor_out_634 , edt_decompressor_out_635 , edt_decompressor_out_636 , edt_decompressor_out_637 ,
        edt_decompressor_out_638 , edt_decompressor_out_639 , edt_decompressor_out_640 , edt_decompressor_out_641 ,
        edt_decompressor_out_642 , edt_decompressor_out_643 , edt_decompressor_out_644 , edt_decompressor_out_645 ,
        edt_decompressor_out_646 , edt_decompressor_out_647 , edt_decompressor_out_648 , edt_decompressor_out_649 ,
        edt_decompressor_out_650 , edt_decompressor_out_651 , edt_decompressor_out_652 , edt_decompressor_out_653 ,
        edt_decompressor_out_654 , edt_decompressor_out_655 , edt_decompressor_out_656 , edt_decompressor_out_657 ,
        edt_decompressor_out_658 , edt_decompressor_out_659 , edt_decompressor_out_660 , edt_decompressor_out_661 ,
        edt_decompressor_out_662 , edt_decompressor_out_663 , edt_decompressor_out_664 , edt_decompressor_out_665 ,
        edt_decompressor_out_666 , edt_decompressor_out_667 , edt_decompressor_out_668 , edt_decompressor_out_669 ,
        edt_decompressor_out_670 , edt_decompressor_out_671 , edt_decompressor_out_672 , edt_decompressor_out_673 ,
        edt_decompressor_out_674 , edt_decompressor_out_675 , edt_decompressor_out_676 , edt_decompressor_out_677 ,
        edt_decompressor_out_678 , edt_decompressor_out_679 , edt_decompressor_out_680 , edt_decompressor_out_681 ,
        edt_decompressor_out_682 , edt_decompressor_out_683 , edt_decompressor_out_684 , edt_decompressor_out_685 ,
        edt_decompressor_out_686 , edt_decompressor_out_687 , edt_decompressor_out_688 , edt_decompressor_out_689 ,
        edt_decompressor_out_690 , edt_decompressor_out_691 , edt_decompressor_out_692 , edt_decompressor_out_693 ,
        edt_decompressor_out_694 , edt_decompressor_out_695 , edt_decompressor_out_696 , edt_decompressor_out_697 ,
        edt_decompressor_out_698 , edt_decompressor_out_699 , edt_decompressor_out_700 , edt_decompressor_out_701 ,
        edt_decompressor_out_702 , edt_decompressor_out_703 , edt_decompressor_out_704 , edt_decompressor_out_705 ,
        edt_decompressor_out_706 , edt_decompressor_out_707 , edt_decompressor_out_708 , edt_decompressor_out_709 ,
        edt_decompressor_out_710 , edt_decompressor_out_711 , edt_decompressor_out_712 , edt_decompressor_out_713 ,
        edt_decompressor_out_714 , edt_decompressor_out_715 , edt_decompressor_out_716 , edt_decompressor_out_717 ,
        edt_decompressor_out_718 , edt_decompressor_out_719 , edt_decompressor_out_720 , edt_decompressor_out_721 ,
        edt_decompressor_out_722 , edt_decompressor_out_723 , edt_decompressor_out_724 , edt_decompressor_out_725 ,
        edt_decompressor_out_726 , edt_decompressor_out_727 , edt_decompressor_out_728 , edt_decompressor_out_729 ,
        edt_decompressor_out_730 , edt_decompressor_out_731 , edt_decompressor_out_732 , edt_decompressor_out_733 ,
        edt_decompressor_out_734 , edt_decompressor_out_735 , edt_decompressor_out_736 , edt_decompressor_out_737 ,
        edt_decompressor_out_738 , edt_decompressor_out_739 , edt_decompressor_out_740 , edt_decompressor_out_741 ,
        edt_decompressor_out_742 , edt_decompressor_out_743 , edt_decompressor_out_744 , edt_decompressor_out_745 ,
        edt_decompressor_out_746 , edt_decompressor_out_747 , edt_decompressor_out_748 , edt_decompressor_out_749 ,
        edt_decompressor_out_750 , edt_decompressor_out_751 , edt_decompressor_out_752 , edt_decompressor_out_753 ,
        edt_decompressor_out_754 , edt_decompressor_out_755 , edt_decompressor_out_756 , edt_decompressor_out_757 ,
        edt_decompressor_out_758 , edt_decompressor_out_759 , edt_decompressor_out_760 , edt_decompressor_out_761 ,
        edt_decompressor_out_762 , edt_decompressor_out_763 , edt_decompressor_out_764 , edt_decompressor_out_765 ,
        edt_decompressor_out_766 , edt_decompressor_out_767 , edt_decompressor_out_768 , edt_decompressor_out_769 ,
        edt_decompressor_out_770 , edt_decompressor_out_771 , edt_decompressor_out_772 , edt_decompressor_out_773 ,
        edt_decompressor_out_774 , edt_decompressor_out_775 , edt_decompressor_out_776 , edt_decompressor_out_777 ,
        edt_decompressor_out_778 , edt_decompressor_out_779 , edt_decompressor_out_780 , edt_decompressor_out_781 ,
        edt_decompressor_out_782 , edt_decompressor_out_783 , edt_decompressor_out_784 , edt_decompressor_out_785 ,
        edt_decompressor_out_786 , edt_decompressor_out_787 , edt_decompressor_out_788 , edt_decompressor_out_789 ,
        edt_decompressor_out_790 , edt_decompressor_out_791 , edt_decompressor_out_792 , edt_decompressor_out_793 ,
        edt_decompressor_out_794 , edt_decompressor_out_795 , edt_update_hfs_netlink_29280 , edt_update_hfs_netlink_29281 ,
        edt_update_hfs_netlink_29282 , edt_update_hfs_netlink_29283 , edt_update_hfs_netlink_29284 , edt_update_hfs_netlink_29285 ,
        edt_update_hfs_netlink_29286 , edt_update_hfs_netlink_29287 , edt_update_hfs_netlink_29288 , edt_update_hfs_netlink_29289 ,
        edt_configuration_hfs_netlink_29290 , edt_configuration_hfs_netlink_29291 , edt_configuration_hfs_netlink_29292 , edt_clock_cts_1 ,
        edt_clock_cts_2 , edt_clock_cts_3 , edt_clock_cts_4 , edt_clock_cts_5 ,
        edt_clock_cts_6 , edt_clock_cts_7 , edt_clock_cts_8 , edt_clock_cts_9 ,
        edt_clock_cts_0_1 , edt_clock_cts_1_1 , edt_clock_cts_2_1 , edt_clock_cts_3_1 ,
        edt_clock_cts_4_1 , edt_clock_cts_5_1 , edt_clock_cts_6_1 , edt_clock_cts_7_1 ) ;
output  edt_channels_out_from_controller_0 , edt_channels_out_from_controller_1 , edt_channels_out_from_controller_2 , edt_channels_out_from_controller_3 ,
        edt_channels_out_from_controller_4 , edt_channels_out_from_controller_5 , edt_channels_out_from_controller_6 , edt_channels_out_from_controller_7 ,
        edt_channels_out_from_controller_8 , edt_channels_out_from_controller_9 , edt_channels_out_from_controller_10 , edt_channels_out_from_controller_11 ,
        edt_channels_out_from_controller_12 , edt_channels_out_from_controller_13 , edt_channels_out_from_controller_14 , masks_for_compactor_0_0 ,
        masks_for_compactor_0_1 , masks_for_compactor_0_2 , masks_for_compactor_0_3 , masks_for_compactor_0_4 ,
        masks_for_compactor_0_5 , masks_for_compactor_0_6 , masks_for_compactor_0_7 , masks_for_compactor_0_8 ,
        masks_for_compactor_0_9 , masks_for_compactor_0_10 , masks_for_compactor_0_11 , masks_for_compactor_0_12 ,
        masks_for_compactor_0_13 , masks_for_compactor_0_14 , masks_for_compactor_0_15 , masks_for_compactor_0_16 ,
        masks_for_compactor_0_17 , masks_for_compactor_0_18 , masks_for_compactor_0_19 , masks_for_compactor_0_20 ,
        masks_for_compactor_0_21 , masks_for_compactor_0_22 , masks_for_compactor_0_23 , masks_for_compactor_0_24 ,
        masks_for_compactor_0_25 , masks_for_compactor_0_26 , masks_for_compactor_0_27 , masks_for_compactor_0_28 ,
        masks_for_compactor_0_29 , masks_for_compactor_0_30 , masks_for_compactor_0_31 , masks_for_compactor_0_32 ,
        masks_for_compactor_0_33 , masks_for_compactor_0_34 , masks_for_compactor_0_35 , masks_for_compactor_0_36 ,
        masks_for_compactor_0_37 , masks_for_compactor_0_38 , masks_for_compactor_0_39 , masks_for_compactor_0_40 ,
        masks_for_compactor_0_41 , masks_for_compactor_0_42 , masks_for_compactor_0_43 , masks_for_compactor_0_44 ,
        masks_for_compactor_0_45 , masks_for_compactor_0_46 , masks_for_compactor_0_47 , masks_for_compactor_0_48 ,
        masks_for_compactor_0_49 , masks_for_compactor_0_50 , masks_for_compactor_0_51 , masks_for_compactor_0_52 ,
        masks_for_compactor_0_53 , masks_for_compactor_1_0 , masks_for_compactor_1_1 , masks_for_compactor_1_2 ,
        masks_for_compactor_1_3 , masks_for_compactor_1_4 , masks_for_compactor_1_5 , masks_for_compactor_1_6 ,
        masks_for_compactor_1_7 , masks_for_compactor_1_8 , masks_for_compactor_1_9 , masks_for_compactor_1_10 ,
        masks_for_compactor_1_11 , masks_for_compactor_1_12 , masks_for_compactor_1_13 , masks_for_compactor_1_14 ,
        masks_for_compactor_1_15 , masks_for_compactor_1_16 , masks_for_compactor_1_17 , masks_for_compactor_1_18 ,
        masks_for_compactor_1_19 , masks_for_compactor_1_20 , masks_for_compactor_1_21 , masks_for_compactor_1_22 ,
        masks_for_compactor_1_23 , masks_for_compactor_1_24 , masks_for_compactor_1_25 , masks_for_compactor_1_26 ,
        masks_for_compactor_1_27 , masks_for_compactor_1_28 , masks_for_compactor_1_29 , masks_for_compactor_1_30 ,
        masks_for_compactor_1_31 , masks_for_compactor_1_32 , masks_for_compactor_1_33 , masks_for_compactor_1_34 ,
        masks_for_compactor_1_35 , masks_for_compactor_1_36 , masks_for_compactor_1_37 , masks_for_compactor_1_38 ,
        masks_for_compactor_1_39 , masks_for_compactor_1_40 , masks_for_compactor_1_41 , masks_for_compactor_1_42 ,
        masks_for_compactor_1_43 , masks_for_compactor_1_44 , masks_for_compactor_1_45 , masks_for_compactor_1_46 ,
        masks_for_compactor_1_47 , masks_for_compactor_1_48 , masks_for_compactor_1_49 , masks_for_compactor_1_50 ,
        masks_for_compactor_1_51 , masks_for_compactor_1_52 , masks_for_compactor_2_0 , masks_for_compactor_2_1 ,
        masks_for_compactor_2_2 , masks_for_compactor_2_3 , masks_for_compactor_2_4 , masks_for_compactor_2_5 ,
        masks_for_compactor_2_6 , masks_for_compactor_2_7 , masks_for_compactor_2_8 , masks_for_compactor_2_9 ,
        masks_for_compactor_2_10 , masks_for_compactor_2_11 , masks_for_compactor_2_12 , masks_for_compactor_2_13 ,
        masks_for_compactor_2_14 , masks_for_compactor_2_15 , masks_for_compactor_2_16 , masks_for_compactor_2_17 ,
        masks_for_compactor_2_18 , masks_for_compactor_2_19 , masks_for_compactor_2_20 , masks_for_compactor_2_21 ,
        masks_for_compactor_2_22 , masks_for_compactor_2_23 , masks_for_compactor_2_24 , masks_for_compactor_2_25 ,
        masks_for_compactor_2_26 , masks_for_compactor_2_27 , masks_for_compactor_2_28 , masks_for_compactor_2_29 ,
        masks_for_compactor_2_30 , masks_for_compactor_2_31 , masks_for_compactor_2_32 , masks_for_compactor_2_33 ,
        masks_for_compactor_2_34 , masks_for_compactor_2_35 , masks_for_compactor_2_36 , masks_for_compactor_2_37 ,
        masks_for_compactor_2_38 , masks_for_compactor_2_39 , masks_for_compactor_2_40 , masks_for_compactor_2_41 ,
        masks_for_compactor_2_42 , masks_for_compactor_2_43 , masks_for_compactor_2_44 , masks_for_compactor_2_45 ,
        masks_for_compactor_2_46 , masks_for_compactor_2_47 , masks_for_compactor_2_48 , masks_for_compactor_2_49 ,
        masks_for_compactor_2_50 , masks_for_compactor_2_51 , masks_for_compactor_2_52 , masks_for_compactor_3_0 ,
        masks_for_compactor_3_1 , masks_for_compactor_3_2 , masks_for_compactor_3_3 , masks_for_compactor_3_4 ,
        masks_for_compactor_3_5 , masks_for_compactor_3_6 , masks_for_compactor_3_7 , masks_for_compactor_3_8 ,
        masks_for_compactor_3_9 , masks_for_compactor_3_10 , masks_for_compactor_3_11 , masks_for_compactor_3_12 ,
        masks_for_compactor_3_13 , masks_for_compactor_3_14 , masks_for_compactor_3_15 , masks_for_compactor_3_16 ,
        masks_for_compactor_3_17 , masks_for_compactor_3_18 , masks_for_compactor_3_19 , masks_for_compactor_3_20 ,
        masks_for_compactor_3_21 , masks_for_compactor_3_22 , masks_for_compactor_3_23 , masks_for_compactor_3_24 ,
        masks_for_compactor_3_25 , masks_for_compactor_3_26 , masks_for_compactor_3_27 , masks_for_compactor_3_28 ,
        masks_for_compactor_3_29 , masks_for_compactor_3_30 , masks_for_compactor_3_31 , masks_for_compactor_3_32 ,
        masks_for_compactor_3_33 , masks_for_compactor_3_34 , masks_for_compactor_3_35 , masks_for_compactor_3_36 ,
        masks_for_compactor_3_37 , masks_for_compactor_3_38 , masks_for_compactor_3_39 , masks_for_compactor_3_40 ,
        masks_for_compactor_3_41 , masks_for_compactor_3_42 , masks_for_compactor_3_43 , masks_for_compactor_3_44 ,
        masks_for_compactor_3_45 , masks_for_compactor_3_46 , masks_for_compactor_3_47 , masks_for_compactor_3_48 ,
        masks_for_compactor_3_49 , masks_for_compactor_3_50 , masks_for_compactor_3_51 , masks_for_compactor_3_52 ,
        masks_for_compactor_4_0 , masks_for_compactor_4_1 , masks_for_compactor_4_2 , masks_for_compactor_4_3 ,
        masks_for_compactor_4_4 , masks_for_compactor_4_5 , masks_for_compactor_4_6 , masks_for_compactor_4_7 ,
        masks_for_compactor_4_8 , masks_for_compactor_4_9 , masks_for_compactor_4_10 , masks_for_compactor_4_11 ,
        masks_for_compactor_4_12 , masks_for_compactor_4_13 , masks_for_compactor_4_14 , masks_for_compactor_4_15 ,
        masks_for_compactor_4_16 , masks_for_compactor_4_17 , masks_for_compactor_4_18 , masks_for_compactor_4_19 ,
        masks_for_compactor_4_20 , masks_for_compactor_4_21 , masks_for_compactor_4_22 , masks_for_compactor_4_23 ,
        masks_for_compactor_4_24 , masks_for_compactor_4_25 , masks_for_compactor_4_26 , masks_for_compactor_4_27 ,
        masks_for_compactor_4_28 , masks_for_compactor_4_29 , masks_for_compactor_4_30 , masks_for_compactor_4_31 ,
        masks_for_compactor_4_32 , masks_for_compactor_4_33 , masks_for_compactor_4_34 , masks_for_compactor_4_35 ,
        masks_for_compactor_4_36 , masks_for_compactor_4_37 , masks_for_compactor_4_38 , masks_for_compactor_4_39 ,
        masks_for_compactor_4_40 , masks_for_compactor_4_41 , masks_for_compactor_4_42 , masks_for_compactor_4_43 ,
        masks_for_compactor_4_44 , masks_for_compactor_4_45 , masks_for_compactor_4_46 , masks_for_compactor_4_47 ,
        masks_for_compactor_4_48 , masks_for_compactor_4_49 , masks_for_compactor_4_50 , masks_for_compactor_4_51 ,
        masks_for_compactor_4_52 , masks_for_compactor_5_0 , masks_for_compactor_5_1 , masks_for_compactor_5_2 ,
        masks_for_compactor_5_3 , masks_for_compactor_5_4 , masks_for_compactor_5_5 , masks_for_compactor_5_6 ,
        masks_for_compactor_5_7 , masks_for_compactor_5_8 , masks_for_compactor_5_9 , masks_for_compactor_5_10 ,
        masks_for_compactor_5_11 , masks_for_compactor_5_12 , masks_for_compactor_5_13 , masks_for_compactor_5_14 ,
        masks_for_compactor_5_15 , masks_for_compactor_5_16 , masks_for_compactor_5_17 , masks_for_compactor_5_18 ,
        masks_for_compactor_5_19 , masks_for_compactor_5_20 , masks_for_compactor_5_21 , masks_for_compactor_5_22 ,
        masks_for_compactor_5_23 , masks_for_compactor_5_24 , masks_for_compactor_5_25 , masks_for_compactor_5_26 ,
        masks_for_compactor_5_27 , masks_for_compactor_5_28 , masks_for_compactor_5_29 , masks_for_compactor_5_30 ,
        masks_for_compactor_5_31 , masks_for_compactor_5_32 , masks_for_compactor_5_33 , masks_for_compactor_5_34 ,
        masks_for_compactor_5_35 , masks_for_compactor_5_36 , masks_for_compactor_5_37 , masks_for_compactor_5_38 ,
        masks_for_compactor_5_39 , masks_for_compactor_5_40 , masks_for_compactor_5_41 , masks_for_compactor_5_42 ,
        masks_for_compactor_5_43 , masks_for_compactor_5_44 , masks_for_compactor_5_45 , masks_for_compactor_5_46 ,
        masks_for_compactor_5_47 , masks_for_compactor_5_48 , masks_for_compactor_5_49 , masks_for_compactor_5_50 ,
        masks_for_compactor_5_51 , masks_for_compactor_5_52 , masks_for_compactor_6_0 , masks_for_compactor_6_1 ,
        masks_for_compactor_6_2 , masks_for_compactor_6_3 , masks_for_compactor_6_4 , masks_for_compactor_6_5 ,
        masks_for_compactor_6_6 , masks_for_compactor_6_7 , masks_for_compactor_6_8 , masks_for_compactor_6_9 ,
        masks_for_compactor_6_10 , masks_for_compactor_6_11 , masks_for_compactor_6_12 , masks_for_compactor_6_13 ,
        masks_for_compactor_6_14 , masks_for_compactor_6_15 , masks_for_compactor_6_16 , masks_for_compactor_6_17 ,
        masks_for_compactor_6_18 , masks_for_compactor_6_19 , masks_for_compactor_6_20 , masks_for_compactor_6_21 ,
        masks_for_compactor_6_22 , masks_for_compactor_6_23 , masks_for_compactor_6_24 , masks_for_compactor_6_25 ,
        masks_for_compactor_6_26 , masks_for_compactor_6_27 , masks_for_compactor_6_28 , masks_for_compactor_6_29 ,
        masks_for_compactor_6_30 , masks_for_compactor_6_31 , masks_for_compactor_6_32 , masks_for_compactor_6_33 ,
        masks_for_compactor_6_34 , masks_for_compactor_6_35 , masks_for_compactor_6_36 , masks_for_compactor_6_37 ,
        masks_for_compactor_6_38 , masks_for_compactor_6_39 , masks_for_compactor_6_40 , masks_for_compactor_6_41 ,
        masks_for_compactor_6_42 , masks_for_compactor_6_43 , masks_for_compactor_6_44 , masks_for_compactor_6_45 ,
        masks_for_compactor_6_46 , masks_for_compactor_6_47 , masks_for_compactor_6_48 , masks_for_compactor_6_49 ,
        masks_for_compactor_6_50 , masks_for_compactor_6_51 , masks_for_compactor_6_52 , masks_for_compactor_7_0 ,
        masks_for_compactor_7_1 , masks_for_compactor_7_2 , masks_for_compactor_7_3 , masks_for_compactor_7_4 ,
        masks_for_compactor_7_5 , masks_for_compactor_7_6 , masks_for_compactor_7_7 , masks_for_compactor_7_8 ,
        masks_for_compactor_7_9 , masks_for_compactor_7_10 , masks_for_compactor_7_11 , masks_for_compactor_7_12 ,
        masks_for_compactor_7_13 , masks_for_compactor_7_14 , masks_for_compactor_7_15 , masks_for_compactor_7_16 ,
        masks_for_compactor_7_17 , masks_for_compactor_7_18 , masks_for_compactor_7_19 , masks_for_compactor_7_20 ,
        masks_for_compactor_7_21 , masks_for_compactor_7_22 , masks_for_compactor_7_23 , masks_for_compactor_7_24 ,
        masks_for_compactor_7_25 , masks_for_compactor_7_26 , masks_for_compactor_7_27 , masks_for_compactor_7_28 ,
        masks_for_compactor_7_29 , masks_for_compactor_7_30 , masks_for_compactor_7_31 , masks_for_compactor_7_32 ,
        masks_for_compactor_7_33 , masks_for_compactor_7_34 , masks_for_compactor_7_35 , masks_for_compactor_7_36 ,
        masks_for_compactor_7_37 , masks_for_compactor_7_38 , masks_for_compactor_7_39 , masks_for_compactor_7_40 ,
        masks_for_compactor_7_41 , masks_for_compactor_7_42 , masks_for_compactor_7_43 , masks_for_compactor_7_44 ,
        masks_for_compactor_7_45 , masks_for_compactor_7_46 , masks_for_compactor_7_47 , masks_for_compactor_7_48 ,
        masks_for_compactor_7_49 , masks_for_compactor_7_50 , masks_for_compactor_7_51 , masks_for_compactor_7_52 ,
        masks_for_compactor_8_0 , masks_for_compactor_8_1 , masks_for_compactor_8_2 , masks_for_compactor_8_3 ,
        masks_for_compactor_8_4 , masks_for_compactor_8_5 , masks_for_compactor_8_6 , masks_for_compactor_8_7 ,
        masks_for_compactor_8_8 , masks_for_compactor_8_9 , masks_for_compactor_8_10 , masks_for_compactor_8_11 ,
        masks_for_compactor_8_12 , masks_for_compactor_8_13 , masks_for_compactor_8_14 , masks_for_compactor_8_15 ,
        masks_for_compactor_8_16 , masks_for_compactor_8_17 , masks_for_compactor_8_18 , masks_for_compactor_8_19 ,
        masks_for_compactor_8_20 , masks_for_compactor_8_21 , masks_for_compactor_8_22 , masks_for_compactor_8_23 ,
        masks_for_compactor_8_24 , masks_for_compactor_8_25 , masks_for_compactor_8_26 , masks_for_compactor_8_27 ,
        masks_for_compactor_8_28 , masks_for_compactor_8_29 , masks_for_compactor_8_30 , masks_for_compactor_8_31 ,
        masks_for_compactor_8_32 , masks_for_compactor_8_33 , masks_for_compactor_8_34 , masks_for_compactor_8_35 ,
        masks_for_compactor_8_36 , masks_for_compactor_8_37 , masks_for_compactor_8_38 , masks_for_compactor_8_39 ,
        masks_for_compactor_8_40 , masks_for_compactor_8_41 , masks_for_compactor_8_42 , masks_for_compactor_8_43 ,
        masks_for_compactor_8_44 , masks_for_compactor_8_45 , masks_for_compactor_8_46 , masks_for_compactor_8_47 ,
        masks_for_compactor_8_48 , masks_for_compactor_8_49 , masks_for_compactor_8_50 , masks_for_compactor_8_51 ,
        masks_for_compactor_8_52 , masks_for_compactor_9_0 , masks_for_compactor_9_1 , masks_for_compactor_9_2 ,
        masks_for_compactor_9_3 , masks_for_compactor_9_4 , masks_for_compactor_9_5 , masks_for_compactor_9_6 ,
        masks_for_compactor_9_7 , masks_for_compactor_9_8 , masks_for_compactor_9_9 , masks_for_compactor_9_10 ,
        masks_for_compactor_9_11 , masks_for_compactor_9_12 , masks_for_compactor_9_13 , masks_for_compactor_9_14 ,
        masks_for_compactor_9_15 , masks_for_compactor_9_16 , masks_for_compactor_9_17 , masks_for_compactor_9_18 ,
        masks_for_compactor_9_19 , masks_for_compactor_9_20 , masks_for_compactor_9_21 , masks_for_compactor_9_22 ,
        masks_for_compactor_9_23 , masks_for_compactor_9_24 , masks_for_compactor_9_25 , masks_for_compactor_9_26 ,
        masks_for_compactor_9_27 , masks_for_compactor_9_28 , masks_for_compactor_9_29 , masks_for_compactor_9_30 ,
        masks_for_compactor_9_31 , masks_for_compactor_9_32 , masks_for_compactor_9_33 , masks_for_compactor_9_34 ,
        masks_for_compactor_9_35 , masks_for_compactor_9_36 , masks_for_compactor_9_37 , masks_for_compactor_9_38 ,
        masks_for_compactor_9_39 , masks_for_compactor_9_40 , masks_for_compactor_9_41 , masks_for_compactor_9_42 ,
        masks_for_compactor_9_43 , masks_for_compactor_9_44 , masks_for_compactor_9_45 , masks_for_compactor_9_46 ,
        masks_for_compactor_9_47 , masks_for_compactor_9_48 , masks_for_compactor_9_49 , masks_for_compactor_9_50 ,
        masks_for_compactor_9_51 , masks_for_compactor_9_52 , masks_for_compactor_10_0 , masks_for_compactor_10_1 ,
        masks_for_compactor_10_2 , masks_for_compactor_10_3 , masks_for_compactor_10_4 , masks_for_compactor_10_5 ,
        masks_for_compactor_10_6 , masks_for_compactor_10_7 , masks_for_compactor_10_8 , masks_for_compactor_10_9 ,
        masks_for_compactor_10_10 , masks_for_compactor_10_11 , masks_for_compactor_10_12 , masks_for_compactor_10_13 ,
        masks_for_compactor_10_14 , masks_for_compactor_10_15 , masks_for_compactor_10_16 , masks_for_compactor_10_17 ,
        masks_for_compactor_10_18 , masks_for_compactor_10_19 , masks_for_compactor_10_20 , masks_for_compactor_10_21 ,
        masks_for_compactor_10_22 , masks_for_compactor_10_23 , masks_for_compactor_10_24 , masks_for_compactor_10_25 ,
        masks_for_compactor_10_26 , masks_for_compactor_10_27 , masks_for_compactor_10_28 , masks_for_compactor_10_29 ,
        masks_for_compactor_10_30 , masks_for_compactor_10_31 , masks_for_compactor_10_32 , masks_for_compactor_10_33 ,
        masks_for_compactor_10_34 , masks_for_compactor_10_35 , masks_for_compactor_10_36 , masks_for_compactor_10_37 ,
        masks_for_compactor_10_38 , masks_for_compactor_10_39 , masks_for_compactor_10_40 , masks_for_compactor_10_41 ,
        masks_for_compactor_10_42 , masks_for_compactor_10_43 , masks_for_compactor_10_44 , masks_for_compactor_10_45 ,
        masks_for_compactor_10_46 , masks_for_compactor_10_47 , masks_for_compactor_10_48 , masks_for_compactor_10_49 ,
        masks_for_compactor_10_50 , masks_for_compactor_10_51 , masks_for_compactor_10_52 , masks_for_compactor_11_0 ,
        masks_for_compactor_11_1 , masks_for_compactor_11_2 , masks_for_compactor_11_3 , masks_for_compactor_11_4 ,
        masks_for_compactor_11_5 , masks_for_compactor_11_6 , masks_for_compactor_11_7 , masks_for_compactor_11_8 ,
        masks_for_compactor_11_9 , masks_for_compactor_11_10 , masks_for_compactor_11_11 , masks_for_compactor_11_12 ,
        masks_for_compactor_11_13 , masks_for_compactor_11_14 , masks_for_compactor_11_15 , masks_for_compactor_11_16 ,
        masks_for_compactor_11_17 , masks_for_compactor_11_18 , masks_for_compactor_11_19 , masks_for_compactor_11_20 ,
        masks_for_compactor_11_21 , masks_for_compactor_11_22 , masks_for_compactor_11_23 , masks_for_compactor_11_24 ,
        masks_for_compactor_11_25 , masks_for_compactor_11_26 , masks_for_compactor_11_27 , masks_for_compactor_11_28 ,
        masks_for_compactor_11_29 , masks_for_compactor_11_30 , masks_for_compactor_11_31 , masks_for_compactor_11_32 ,
        masks_for_compactor_11_33 , masks_for_compactor_11_34 , masks_for_compactor_11_35 , masks_for_compactor_11_36 ,
        masks_for_compactor_11_37 , masks_for_compactor_11_38 , masks_for_compactor_11_39 , masks_for_compactor_11_40 ,
        masks_for_compactor_11_41 , masks_for_compactor_11_42 , masks_for_compactor_11_43 , masks_for_compactor_11_44 ,
        masks_for_compactor_11_45 , masks_for_compactor_11_46 , masks_for_compactor_11_47 , masks_for_compactor_11_48 ,
        masks_for_compactor_11_49 , masks_for_compactor_11_50 , masks_for_compactor_11_51 , masks_for_compactor_11_52 ,
        masks_for_compactor_12_0 , masks_for_compactor_12_1 , masks_for_compactor_12_2 , masks_for_compactor_12_3 ,
        masks_for_compactor_12_4 , masks_for_compactor_12_5 , masks_for_compactor_12_6 , masks_for_compactor_12_7 ,
        masks_for_compactor_12_8 , masks_for_compactor_12_9 , masks_for_compactor_12_10 , masks_for_compactor_12_11 ,
        masks_for_compactor_12_12 , masks_for_compactor_12_13 , masks_for_compactor_12_14 , masks_for_compactor_12_15 ,
        masks_for_compactor_12_16 , masks_for_compactor_12_17 , masks_for_compactor_12_18 , masks_for_compactor_12_19 ,
        masks_for_compactor_12_20 , masks_for_compactor_12_21 , masks_for_compactor_12_22 , masks_for_compactor_12_23 ,
        masks_for_compactor_12_24 , masks_for_compactor_12_25 , masks_for_compactor_12_26 , masks_for_compactor_12_27 ,
        masks_for_compactor_12_28 , masks_for_compactor_12_29 , masks_for_compactor_12_30 , masks_for_compactor_12_31 ,
        masks_for_compactor_12_32 , masks_for_compactor_12_33 , masks_for_compactor_12_34 , masks_for_compactor_12_35 ,
        masks_for_compactor_12_36 , masks_for_compactor_12_37 , masks_for_compactor_12_38 , masks_for_compactor_12_39 ,
        masks_for_compactor_12_40 , masks_for_compactor_12_41 , masks_for_compactor_12_42 , masks_for_compactor_12_43 ,
        masks_for_compactor_12_44 , masks_for_compactor_12_45 , masks_for_compactor_12_46 , masks_for_compactor_12_47 ,
        masks_for_compactor_12_48 , masks_for_compactor_12_49 , masks_for_compactor_12_50 , masks_for_compactor_12_51 ,
        masks_for_compactor_12_52 , masks_for_compactor_13_0 , masks_for_compactor_13_1 , masks_for_compactor_13_2 ,
        masks_for_compactor_13_3 , masks_for_compactor_13_4 , masks_for_compactor_13_5 , masks_for_compactor_13_6 ,
        masks_for_compactor_13_7 , masks_for_compactor_13_8 , masks_for_compactor_13_9 , masks_for_compactor_13_10 ,
        masks_for_compactor_13_11 , masks_for_compactor_13_12 , masks_for_compactor_13_13 , masks_for_compactor_13_14 ,
        masks_for_compactor_13_15 , masks_for_compactor_13_16 , masks_for_compactor_13_17 , masks_for_compactor_13_18 ,
        masks_for_compactor_13_19 , masks_for_compactor_13_20 , masks_for_compactor_13_21 , masks_for_compactor_13_22 ,
        masks_for_compactor_13_23 , masks_for_compactor_13_24 , masks_for_compactor_13_25 , masks_for_compactor_13_26 ,
        masks_for_compactor_13_27 , masks_for_compactor_13_28 , masks_for_compactor_13_29 , masks_for_compactor_13_30 ,
        masks_for_compactor_13_31 , masks_for_compactor_13_32 , masks_for_compactor_13_33 , masks_for_compactor_13_34 ,
        masks_for_compactor_13_35 , masks_for_compactor_13_36 , masks_for_compactor_13_37 , masks_for_compactor_13_38 ,
        masks_for_compactor_13_39 , masks_for_compactor_13_40 , masks_for_compactor_13_41 , masks_for_compactor_13_42 ,
        masks_for_compactor_13_43 , masks_for_compactor_13_44 , masks_for_compactor_13_45 , masks_for_compactor_13_46 ,
        masks_for_compactor_13_47 , masks_for_compactor_13_48 , masks_for_compactor_13_49 , masks_for_compactor_13_50 ,
        masks_for_compactor_13_51 , masks_for_compactor_13_52 , masks_for_compactor_14_0 , masks_for_compactor_14_1 ,
        masks_for_compactor_14_2 , masks_for_compactor_14_3 , masks_for_compactor_14_4 , masks_for_compactor_14_5 ,
        masks_for_compactor_14_6 , masks_for_compactor_14_7 , masks_for_compactor_14_8 , masks_for_compactor_14_9 ,
        masks_for_compactor_14_10 , masks_for_compactor_14_11 , masks_for_compactor_14_12 , masks_for_compactor_14_13 ,
        masks_for_compactor_14_14 , masks_for_compactor_14_15 , masks_for_compactor_14_16 , masks_for_compactor_14_17 ,
        masks_for_compactor_14_18 , masks_for_compactor_14_19 , masks_for_compactor_14_20 , masks_for_compactor_14_21 ,
        masks_for_compactor_14_22 , masks_for_compactor_14_23 , masks_for_compactor_14_24 , masks_for_compactor_14_25 ,
        masks_for_compactor_14_26 , masks_for_compactor_14_27 , masks_for_compactor_14_28 , masks_for_compactor_14_29 ,
        masks_for_compactor_14_30 , masks_for_compactor_14_31 , masks_for_compactor_14_32 , masks_for_compactor_14_33 ,
        masks_for_compactor_14_34 , masks_for_compactor_14_35 , masks_for_compactor_14_36 , masks_for_compactor_14_37 ,
        masks_for_compactor_14_38 , masks_for_compactor_14_39 , masks_for_compactor_14_40 , masks_for_compactor_14_41 ,
        masks_for_compactor_14_42 , masks_for_compactor_14_43 , masks_for_compactor_14_44 , masks_for_compactor_14_45 ,
        masks_for_compactor_14_46 , masks_for_compactor_14_47 , masks_for_compactor_14_48 , masks_for_compactor_14_49 ,
        masks_for_compactor_14_50 , masks_for_compactor_14_51 , masks_for_compactor_14_52 , edt_scan_in_0 ,
        edt_scan_in_1 , edt_scan_in_2 , edt_scan_in_3 , edt_scan_in_4 ,
        edt_scan_in_5 , edt_scan_in_6 , edt_scan_in_7 , edt_scan_in_8 ,
        edt_scan_in_9 , edt_scan_in_10 , edt_scan_in_11 , edt_scan_in_12 ,
        edt_scan_in_13 , edt_scan_in_14 , edt_scan_in_15 , edt_scan_in_16 ,
        edt_scan_in_17 , edt_scan_in_18 , edt_scan_in_19 , edt_scan_in_20 ,
        edt_scan_in_21 , edt_scan_in_22 , edt_scan_in_23 , edt_scan_in_24 ,
        edt_scan_in_25 , edt_scan_in_26 , edt_scan_in_27 , edt_scan_in_28 ,
        edt_scan_in_29 , edt_scan_in_30 , edt_scan_in_31 , edt_scan_in_32 ,
        edt_scan_in_33 , edt_scan_in_34 , edt_scan_in_35 , edt_scan_in_36 ,
        edt_scan_in_37 , edt_scan_in_38 , edt_scan_in_39 , edt_scan_in_40 ,
        edt_scan_in_41 , edt_scan_in_42 , edt_scan_in_43 , edt_scan_in_44 ,
        edt_scan_in_45 , edt_scan_in_46 , edt_scan_in_47 , edt_scan_in_48 ,
        edt_scan_in_49 , edt_scan_in_50 , edt_scan_in_51 , edt_scan_in_52 ,
        edt_scan_in_53 , edt_scan_in_54 , edt_scan_in_55 , edt_scan_in_56 ,
        edt_scan_in_57 , edt_scan_in_58 , edt_scan_in_59 , edt_scan_in_60 ,
        edt_scan_in_61 , edt_scan_in_62 , edt_scan_in_63 , edt_scan_in_64 ,
        edt_scan_in_65 , edt_scan_in_66 , edt_scan_in_67 , edt_scan_in_68 ,
        edt_scan_in_69 , edt_scan_in_70 , edt_scan_in_71 , edt_scan_in_72 ,
        edt_scan_in_73 , edt_scan_in_74 , edt_scan_in_75 , edt_scan_in_76 ,
        edt_scan_in_77 , edt_scan_in_78 , edt_scan_in_79 , edt_scan_in_80 ,
        edt_scan_in_81 , edt_scan_in_82 , edt_scan_in_83 , edt_scan_in_84 ,
        edt_scan_in_85 , edt_scan_in_86 , edt_scan_in_87 , edt_scan_in_88 ,
        edt_scan_in_89 , edt_scan_in_90 , edt_scan_in_91 , edt_scan_in_92 ,
        edt_scan_in_93 , edt_scan_in_94 , edt_scan_in_95 , edt_scan_in_96 ,
        edt_scan_in_97 , edt_scan_in_98 , edt_scan_in_99 , edt_scan_in_100 ,
        edt_scan_in_101 , edt_scan_in_102 , edt_scan_in_103 , edt_scan_in_104 ,
        edt_scan_in_105 , edt_scan_in_106 , edt_scan_in_107 , edt_scan_in_108 ,
        edt_scan_in_109 , edt_scan_in_110 , edt_scan_in_111 , edt_scan_in_112 ,
        edt_scan_in_113 , edt_scan_in_114 , edt_scan_in_115 , edt_scan_in_116 ,
        edt_scan_in_117 , edt_scan_in_118 , edt_scan_in_119 , edt_scan_in_120 ,
        edt_scan_in_121 , edt_scan_in_122 , edt_scan_in_123 , edt_scan_in_124 ,
        edt_scan_in_125 , edt_scan_in_126 , edt_scan_in_127 , edt_scan_in_128 ,
        edt_scan_in_129 , edt_scan_in_130 , edt_scan_in_131 , edt_scan_in_132 ,
        edt_scan_in_133 , edt_scan_in_134 , edt_scan_in_135 , edt_scan_in_136 ,
        edt_scan_in_137 , edt_scan_in_138 , edt_scan_in_139 , edt_scan_in_140 ,
        edt_scan_in_141 , edt_scan_in_142 , edt_scan_in_143 , edt_scan_in_144 ,
        edt_scan_in_145 , edt_scan_in_146 , edt_scan_in_147 , edt_scan_in_148 ,
        edt_scan_in_149 , edt_scan_in_150 , edt_scan_in_151 , edt_scan_in_152 ,
        edt_scan_in_153 , edt_scan_in_154 , edt_scan_in_155 , edt_scan_in_156 ,
        edt_scan_in_157 , edt_scan_in_158 , edt_scan_in_159 , edt_scan_in_160 ,
        edt_scan_in_161 , edt_scan_in_162 , edt_scan_in_163 , edt_scan_in_164 ,
        edt_scan_in_165 , edt_scan_in_166 , edt_scan_in_167 , edt_scan_in_168 ,
        edt_scan_in_169 , edt_scan_in_170 , edt_scan_in_171 , edt_scan_in_172 ,
        edt_scan_in_173 , edt_scan_in_174 , edt_scan_in_175 , edt_scan_in_176 ,
        edt_scan_in_177 , edt_scan_in_178 , edt_scan_in_179 , edt_scan_in_180 ,
        edt_scan_in_181 , edt_scan_in_182 , edt_scan_in_183 , edt_scan_in_184 ,
        edt_scan_in_185 , edt_scan_in_186 , edt_scan_in_187 , edt_scan_in_188 ,
        edt_scan_in_189 , edt_scan_in_190 , edt_scan_in_191 , edt_scan_in_192 ,
        edt_scan_in_193 , edt_scan_in_194 , edt_scan_in_195 , edt_scan_in_196 ,
        edt_scan_in_197 , edt_scan_in_198 , edt_scan_in_199 , edt_scan_in_200 ,
        edt_scan_in_201 , edt_scan_in_202 , edt_scan_in_203 , edt_scan_in_204 ,
        edt_scan_in_205 , edt_scan_in_206 , edt_scan_in_207 , edt_scan_in_208 ,
        edt_scan_in_209 , edt_scan_in_210 , edt_scan_in_211 , edt_scan_in_212 ,
        edt_scan_in_213 , edt_scan_in_214 , edt_scan_in_215 , edt_scan_in_216 ,
        edt_scan_in_217 , edt_scan_in_218 , edt_scan_in_219 , edt_scan_in_220 ,
        edt_scan_in_221 , edt_scan_in_222 , edt_scan_in_223 , edt_scan_in_224 ,
        edt_scan_in_225 , edt_scan_in_226 , edt_scan_in_227 , edt_scan_in_228 ,
        edt_scan_in_229 , edt_scan_in_230 , edt_scan_in_231 , edt_scan_in_232 ,
        edt_scan_in_233 , edt_scan_in_234 , edt_scan_in_235 , edt_scan_in_236 ,
        edt_scan_in_237 , edt_scan_in_238 , edt_scan_in_239 , edt_scan_in_240 ,
        edt_scan_in_241 , edt_scan_in_242 , edt_scan_in_243 , edt_scan_in_244 ,
        edt_scan_in_245 , edt_scan_in_246 , edt_scan_in_247 , edt_scan_in_248 ,
        edt_scan_in_249 , edt_scan_in_250 , edt_scan_in_251 , edt_scan_in_252 ,
        edt_scan_in_253 , edt_scan_in_254 , edt_scan_in_255 , edt_scan_in_256 ,
        edt_scan_in_257 , edt_scan_in_258 , edt_scan_in_259 , edt_scan_in_260 ,
        edt_scan_in_261 , edt_scan_in_262 , edt_scan_in_263 , edt_scan_in_264 ,
        edt_scan_in_265 , edt_scan_in_266 , edt_scan_in_267 , edt_scan_in_268 ,
        edt_scan_in_269 , edt_scan_in_270 , edt_scan_in_271 , edt_scan_in_272 ,
        edt_scan_in_273 , edt_scan_in_274 , edt_scan_in_275 , edt_scan_in_276 ,
        edt_scan_in_277 , edt_scan_in_278 , edt_scan_in_279 , edt_scan_in_280 ,
        edt_scan_in_281 , edt_scan_in_282 , edt_scan_in_283 , edt_scan_in_284 ,
        edt_scan_in_285 , edt_scan_in_286 , edt_scan_in_287 , edt_scan_in_288 ,
        edt_scan_in_289 , edt_scan_in_290 , edt_scan_in_291 , edt_scan_in_292 ,
        edt_scan_in_293 , edt_scan_in_294 , edt_scan_in_295 , edt_scan_in_296 ,
        edt_scan_in_297 , edt_scan_in_298 , edt_scan_in_299 , edt_scan_in_300 ,
        edt_scan_in_301 , edt_scan_in_302 , edt_scan_in_303 , edt_scan_in_304 ,
        edt_scan_in_305 , edt_scan_in_306 , edt_scan_in_307 , edt_scan_in_308 ,
        edt_scan_in_309 , edt_scan_in_310 , edt_scan_in_311 , edt_scan_in_312 ,
        edt_scan_in_313 , edt_scan_in_314 , edt_scan_in_315 , edt_scan_in_316 ,
        edt_scan_in_317 , edt_scan_in_318 , edt_scan_in_319 , edt_scan_in_320 ,
        edt_scan_in_321 , edt_scan_in_322 , edt_scan_in_323 , edt_scan_in_324 ,
        edt_scan_in_325 , edt_scan_in_326 , edt_scan_in_327 , edt_scan_in_328 ,
        edt_scan_in_329 , edt_scan_in_330 , edt_scan_in_331 , edt_scan_in_332 ,
        edt_scan_in_333 , edt_scan_in_334 , edt_scan_in_335 , edt_scan_in_336 ,
        edt_scan_in_337 , edt_scan_in_338 , edt_scan_in_339 , edt_scan_in_340 ,
        edt_scan_in_341 , edt_scan_in_342 , edt_scan_in_343 , edt_scan_in_344 ,
        edt_scan_in_345 , edt_scan_in_346 , edt_scan_in_347 , edt_scan_in_348 ,
        edt_scan_in_349 , edt_scan_in_350 , edt_scan_in_351 , edt_scan_in_352 ,
        edt_scan_in_353 , edt_scan_in_354 , edt_scan_in_355 , edt_scan_in_356 ,
        edt_scan_in_357 , edt_scan_in_358 , edt_scan_in_359 , edt_scan_in_360 ,
        edt_scan_in_361 , edt_scan_in_362 , edt_scan_in_363 , edt_scan_in_364 ,
        edt_scan_in_365 , edt_scan_in_366 , edt_scan_in_367 , edt_scan_in_368 ,
        edt_scan_in_369 , edt_scan_in_370 , edt_scan_in_371 , edt_scan_in_372 ,
        edt_scan_in_373 , edt_scan_in_374 , edt_scan_in_375 , edt_scan_in_376 ,
        edt_scan_in_377 , edt_scan_in_378 , edt_scan_in_379 , edt_scan_in_380 ,
        edt_scan_in_381 , edt_scan_in_382 , edt_scan_in_383 , edt_scan_in_384 ,
        edt_scan_in_385 , edt_scan_in_386 , edt_scan_in_387 , edt_scan_in_388 ,
        edt_scan_in_389 , edt_scan_in_390 , edt_scan_in_391 , edt_scan_in_392 ,
        edt_scan_in_393 , edt_scan_in_394 , edt_scan_in_395 , edt_scan_in_396 ,
        edt_scan_in_397 , edt_scan_in_398 , edt_scan_in_399 , edt_scan_in_400 ,
        edt_scan_in_401 , edt_scan_in_402 , edt_scan_in_403 , edt_scan_in_404 ,
        edt_scan_in_405 , edt_scan_in_406 , edt_scan_in_407 , edt_scan_in_408 ,
        edt_scan_in_409 , edt_scan_in_410 , edt_scan_in_411 , edt_scan_in_412 ,
        edt_scan_in_413 , edt_scan_in_414 , edt_scan_in_415 , edt_scan_in_416 ,
        edt_scan_in_417 , edt_scan_in_418 , edt_scan_in_419 , edt_scan_in_420 ,
        edt_scan_in_421 , edt_scan_in_422 , edt_scan_in_423 , edt_scan_in_424 ,
        edt_scan_in_425 , edt_scan_in_426 , edt_scan_in_427 , edt_scan_in_428 ,
        edt_scan_in_429 , edt_scan_in_430 , edt_scan_in_431 , edt_scan_in_432 ,
        edt_scan_in_433 , edt_scan_in_434 , edt_scan_in_435 , edt_scan_in_436 ,
        edt_scan_in_437 , edt_scan_in_438 , edt_scan_in_439 , edt_scan_in_440 ,
        edt_scan_in_441 , edt_scan_in_442 , edt_scan_in_443 , edt_scan_in_444 ,
        edt_scan_in_445 , edt_scan_in_446 , edt_scan_in_447 , edt_scan_in_448 ,
        edt_scan_in_449 , edt_scan_in_450 , edt_scan_in_451 , edt_scan_in_452 ,
        edt_scan_in_453 , edt_scan_in_454 , edt_scan_in_455 , edt_scan_in_456 ,
        edt_scan_in_457 , edt_scan_in_458 , edt_scan_in_459 , edt_scan_in_460 ,
        edt_scan_in_461 , edt_scan_in_462 , edt_scan_in_463 , edt_scan_in_464 ,
        edt_scan_in_465 , edt_scan_in_466 , edt_scan_in_467 , edt_scan_in_468 ,
        edt_scan_in_469 , edt_scan_in_470 , edt_scan_in_471 , edt_scan_in_472 ,
        edt_scan_in_473 , edt_scan_in_474 , edt_scan_in_475 , edt_scan_in_476 ,
        edt_scan_in_477 , edt_scan_in_478 , edt_scan_in_479 , edt_scan_in_480 ,
        edt_scan_in_481 , edt_scan_in_482 , edt_scan_in_483 , edt_scan_in_484 ,
        edt_scan_in_485 , edt_scan_in_486 , edt_scan_in_487 , edt_scan_in_488 ,
        edt_scan_in_489 , edt_scan_in_490 , edt_scan_in_491 , edt_scan_in_492 ,
        edt_scan_in_493 , edt_scan_in_494 , edt_scan_in_495 , edt_scan_in_496 ,
        edt_scan_in_497 , edt_scan_in_498 , edt_scan_in_499 , edt_scan_in_500 ,
        edt_scan_in_501 , edt_scan_in_502 , edt_scan_in_503 , edt_scan_in_504 ,
        edt_scan_in_505 , edt_scan_in_506 , edt_scan_in_507 , edt_scan_in_508 ,
        edt_scan_in_509 , edt_scan_in_510 , edt_scan_in_511 , edt_scan_in_512 ,
        edt_scan_in_513 , edt_scan_in_514 , edt_scan_in_515 , edt_scan_in_516 ,
        edt_scan_in_517 , edt_scan_in_518 , edt_scan_in_519 , edt_scan_in_520 ,
        edt_scan_in_521 , edt_scan_in_522 , edt_scan_in_523 , edt_scan_in_524 ,
        edt_scan_in_525 , edt_scan_in_526 , edt_scan_in_527 , edt_scan_in_528 ,
        edt_scan_in_529 , edt_scan_in_530 , edt_scan_in_531 , edt_scan_in_532 ,
        edt_scan_in_533 , edt_scan_in_534 , edt_scan_in_535 , edt_scan_in_536 ,
        edt_scan_in_537 , edt_scan_in_538 , edt_scan_in_539 , edt_scan_in_540 ,
        edt_scan_in_541 , edt_scan_in_542 , edt_scan_in_543 , edt_scan_in_544 ,
        edt_scan_in_545 , edt_scan_in_546 , edt_scan_in_547 , edt_scan_in_548 ,
        edt_scan_in_549 , edt_scan_in_550 , edt_scan_in_551 , edt_scan_in_552 ,
        edt_scan_in_553 , edt_scan_in_554 , edt_scan_in_555 , edt_scan_in_556 ,
        edt_scan_in_557 , edt_scan_in_558 , edt_scan_in_559 , edt_scan_in_560 ,
        edt_scan_in_561 , edt_scan_in_562 , edt_scan_in_563 , edt_scan_in_564 ,
        edt_scan_in_565 , edt_scan_in_566 , edt_scan_in_567 , edt_scan_in_568 ,
        edt_scan_in_569 , edt_scan_in_570 , edt_scan_in_571 , edt_scan_in_572 ,
        edt_scan_in_573 , edt_scan_in_574 , edt_scan_in_575 , edt_scan_in_576 ,
        edt_scan_in_577 , edt_scan_in_578 , edt_scan_in_579 , edt_scan_in_580 ,
        edt_scan_in_581 , edt_scan_in_582 , edt_scan_in_583 , edt_scan_in_584 ,
        edt_scan_in_585 , edt_scan_in_586 , edt_scan_in_587 , edt_scan_in_588 ,
        edt_scan_in_589 , edt_scan_in_590 , edt_scan_in_591 , edt_scan_in_592 ,
        edt_scan_in_593 , edt_scan_in_594 , edt_scan_in_595 , edt_scan_in_596 ,
        edt_scan_in_597 , edt_scan_in_598 , edt_scan_in_599 , edt_scan_in_600 ,
        edt_scan_in_601 , edt_scan_in_602 , edt_scan_in_603 , edt_scan_in_604 ,
        edt_scan_in_605 , edt_scan_in_606 , edt_scan_in_607 , edt_scan_in_608 ,
        edt_scan_in_609 , edt_scan_in_610 , edt_scan_in_611 , edt_scan_in_612 ,
        edt_scan_in_613 , edt_scan_in_614 , edt_scan_in_615 , edt_scan_in_616 ,
        edt_scan_in_617 , edt_scan_in_618 , edt_scan_in_619 , edt_scan_in_620 ,
        edt_scan_in_621 , edt_scan_in_622 , edt_scan_in_623 , edt_scan_in_624 ,
        edt_scan_in_625 , edt_scan_in_626 , edt_scan_in_627 , edt_scan_in_628 ,
        edt_scan_in_629 , edt_scan_in_630 , edt_scan_in_631 , edt_scan_in_632 ,
        edt_scan_in_633 , edt_scan_in_634 , edt_scan_in_635 , edt_scan_in_636 ,
        edt_scan_in_637 , edt_scan_in_638 , edt_scan_in_639 , edt_scan_in_640 ,
        edt_scan_in_641 , edt_scan_in_642 , edt_scan_in_643 , edt_scan_in_644 ,
        edt_scan_in_645 , edt_scan_in_646 , edt_scan_in_647 , edt_scan_in_648 ,
        edt_scan_in_649 , edt_scan_in_650 , edt_scan_in_651 , edt_scan_in_652 ,
        edt_scan_in_653 , edt_scan_in_654 , edt_scan_in_655 , edt_scan_in_656 ,
        edt_scan_in_657 , edt_scan_in_658 , edt_scan_in_659 , edt_scan_in_660 ,
        edt_scan_in_661 , edt_scan_in_662 , edt_scan_in_663 , edt_scan_in_664 ,
        edt_scan_in_665 , edt_scan_in_666 , edt_scan_in_667 , edt_scan_in_668 ,
        edt_scan_in_669 , edt_scan_in_670 , edt_scan_in_671 , edt_scan_in_672 ,
        edt_scan_in_673 , edt_scan_in_674 , edt_scan_in_675 , edt_scan_in_676 ,
        edt_scan_in_677 , edt_scan_in_678 , edt_scan_in_679 , edt_scan_in_680 ,
        edt_scan_in_681 , edt_scan_in_682 , edt_scan_in_683 , edt_scan_in_684 ,
        edt_scan_in_685 , edt_scan_in_686 , edt_scan_in_687 , edt_scan_in_688 ,
        edt_scan_in_689 , edt_scan_in_690 , edt_scan_in_691 , edt_scan_in_692 ,
        edt_scan_in_693 , edt_scan_in_694 , edt_scan_in_695 , edt_scan_in_696 ,
        edt_scan_in_697 , edt_scan_in_698 , edt_scan_in_699 , edt_scan_in_700 ,
        edt_scan_in_701 , edt_scan_in_702 , edt_scan_in_703 , edt_scan_in_704 ,
        edt_scan_in_705 , edt_scan_in_706 , edt_scan_in_707 , edt_scan_in_708 ,
        edt_scan_in_709 , edt_scan_in_710 , edt_scan_in_711 , edt_scan_in_712 ,
        edt_scan_in_713 , edt_scan_in_714 , edt_scan_in_715 , edt_scan_in_716 ,
        edt_scan_in_717 , edt_scan_in_718 , edt_scan_in_719 , edt_scan_in_720 ,
        edt_scan_in_721 , edt_scan_in_722 , edt_scan_in_723 , edt_scan_in_724 ,
        edt_scan_in_725 , edt_scan_in_726 , edt_scan_in_727 , edt_scan_in_728 ,
        edt_scan_in_729 , edt_scan_in_730 , edt_scan_in_731 , edt_scan_in_732 ,
        edt_scan_in_733 , edt_scan_in_734 , edt_scan_in_735 , edt_scan_in_736 ,
        edt_scan_in_737 , edt_scan_in_738 , edt_scan_in_739 , edt_scan_in_740 ,
        edt_scan_in_741 , edt_scan_in_742 , edt_scan_in_743 , edt_scan_in_744 ,
        edt_scan_in_745 , edt_scan_in_746 , edt_scan_in_747 , edt_scan_in_748 ,
        edt_scan_in_749 , edt_scan_in_750 , edt_scan_in_751 , edt_scan_in_752 ,
        edt_scan_in_753 , edt_scan_in_754 , edt_scan_in_755 , edt_scan_in_756 ,
        edt_scan_in_757 , edt_scan_in_758 , edt_scan_in_759 , edt_scan_in_760 ,
        edt_scan_in_761 , edt_scan_in_762 , edt_scan_in_763 , edt_scan_in_764 ,
        edt_scan_in_765 , edt_scan_in_766 , edt_scan_in_767 , edt_scan_in_768 ,
        edt_scan_in_769 , edt_scan_in_770 , edt_scan_in_771 , edt_scan_in_772 ,
        edt_scan_in_773 , edt_scan_in_774 , edt_scan_in_775 , edt_scan_in_776 ,
        edt_scan_in_777 , edt_scan_in_778 , edt_scan_in_779 , edt_scan_in_780 ,
        edt_scan_in_781 , edt_scan_in_782 , edt_scan_in_783 , edt_scan_in_784 ,
        edt_scan_in_785 , edt_scan_in_786 , edt_scan_in_787 , edt_scan_in_788 ,
        edt_scan_in_789 , edt_scan_in_790 , edt_scan_in_791 , edt_scan_in_792 ,
        edt_scan_in_793 , edt_scan_in_794 , edt_scan_in_795 ;
input   edt_channels_in_0 , edt_channels_in_1 , edt_channels_in_2 , edt_channels_in_3 ,
        edt_channels_in_4 , edt_channels_in_5 , edt_channels_in_6 , edt_channels_in_7 ,
        edt_channels_in_8 , edt_channels_in_9 , edt_channels_in_10 , edt_channels_in_11 ,
        edt_channels_in_12 , edt_channels_in_13 , edt_channels_in_14 , edt_clock ,
        edt_update , edt_configuration , edt_shift_const_en , edt_decompressor_out_0 ,
        edt_decompressor_out_1 , edt_decompressor_out_2 , edt_decompressor_out_3 , edt_decompressor_out_4 ,
        edt_decompressor_out_5 , edt_decompressor_out_6 , edt_decompressor_out_7 , edt_decompressor_out_8 ,
        edt_decompressor_out_9 , edt_decompressor_out_10 , edt_decompressor_out_11 , edt_decompressor_out_12 ,
        edt_decompressor_out_13 , edt_decompressor_out_14 , edt_decompressor_out_15 , edt_decompressor_out_16 ,
        edt_decompressor_out_17 , edt_decompressor_out_18 , edt_decompressor_out_19 , edt_decompressor_out_20 ,
        edt_decompressor_out_21 , edt_decompressor_out_22 , edt_decompressor_out_23 , edt_decompressor_out_24 ,
        edt_decompressor_out_25 , edt_decompressor_out_26 , edt_decompressor_out_27 , edt_decompressor_out_28 ,
        edt_decompressor_out_29 , edt_decompressor_out_30 , edt_decompressor_out_31 , edt_decompressor_out_32 ,
        edt_decompressor_out_33 , edt_decompressor_out_34 , edt_decompressor_out_35 , edt_decompressor_out_36 ,
        edt_decompressor_out_37 , edt_decompressor_out_38 , edt_decompressor_out_39 , edt_decompressor_out_40 ,
        edt_decompressor_out_41 , edt_decompressor_out_42 , edt_decompressor_out_43 , edt_decompressor_out_44 ,
        edt_decompressor_out_45 , edt_decompressor_out_46 , edt_decompressor_out_47 , edt_decompressor_out_48 ,
        edt_decompressor_out_49 , edt_decompressor_out_50 , edt_decompressor_out_51 , edt_decompressor_out_52 ,
        edt_decompressor_out_53 , edt_decompressor_out_54 , edt_decompressor_out_55 , edt_decompressor_out_56 ,
        edt_decompressor_out_57 , edt_decompressor_out_58 , edt_decompressor_out_59 , edt_decompressor_out_60 ,
        edt_decompressor_out_61 , edt_decompressor_out_62 , edt_decompressor_out_63 , edt_decompressor_out_64 ,
        edt_decompressor_out_65 , edt_decompressor_out_66 , edt_decompressor_out_67 , edt_decompressor_out_68 ,
        edt_decompressor_out_69 , edt_decompressor_out_70 , edt_decompressor_out_71 , edt_decompressor_out_72 ,
        edt_decompressor_out_73 , edt_decompressor_out_74 , edt_decompressor_out_75 , edt_decompressor_out_76 ,
        edt_decompressor_out_77 , edt_decompressor_out_78 , edt_decompressor_out_79 , edt_decompressor_out_80 ,
        edt_decompressor_out_81 , edt_decompressor_out_82 , edt_decompressor_out_83 , edt_decompressor_out_84 ,
        edt_decompressor_out_85 , edt_decompressor_out_86 , edt_decompressor_out_87 , edt_decompressor_out_88 ,
        edt_decompressor_out_89 , edt_decompressor_out_90 , edt_decompressor_out_91 , edt_decompressor_out_92 ,
        edt_decompressor_out_93 , edt_decompressor_out_94 , edt_decompressor_out_95 , edt_decompressor_out_96 ,
        edt_decompressor_out_97 , edt_decompressor_out_98 , edt_decompressor_out_99 , edt_decompressor_out_100 ,
        edt_decompressor_out_101 , edt_decompressor_out_102 , edt_decompressor_out_103 , edt_decompressor_out_104 ,
        edt_decompressor_out_105 , edt_decompressor_out_106 , edt_decompressor_out_107 , edt_decompressor_out_108 ,
        edt_decompressor_out_109 , edt_decompressor_out_110 , edt_decompressor_out_111 , edt_decompressor_out_112 ,
        edt_decompressor_out_113 , edt_decompressor_out_114 , edt_decompressor_out_115 , edt_decompressor_out_116 ,
        edt_decompressor_out_117 , edt_decompressor_out_118 , edt_decompressor_out_119 , edt_decompressor_out_120 ,
        edt_decompressor_out_121 , edt_decompressor_out_122 , edt_decompressor_out_123 , edt_decompressor_out_124 ,
        edt_decompressor_out_125 , edt_decompressor_out_126 , edt_decompressor_out_127 , edt_decompressor_out_128 ,
        edt_decompressor_out_129 , edt_decompressor_out_130 , edt_decompressor_out_131 , edt_decompressor_out_132 ,
        edt_decompressor_out_133 , edt_decompressor_out_134 , edt_decompressor_out_135 , edt_decompressor_out_136 ,
        edt_decompressor_out_137 , edt_decompressor_out_138 , edt_decompressor_out_139 , edt_decompressor_out_140 ,
        edt_decompressor_out_141 , edt_decompressor_out_142 , edt_decompressor_out_143 , edt_decompressor_out_144 ,
        edt_decompressor_out_145 , edt_decompressor_out_146 , edt_decompressor_out_147 , edt_decompressor_out_148 ,
        edt_decompressor_out_149 , edt_decompressor_out_150 , edt_decompressor_out_151 , edt_decompressor_out_152 ,
        edt_decompressor_out_153 , edt_decompressor_out_154 , edt_decompressor_out_155 , edt_decompressor_out_156 ,
        edt_decompressor_out_157 , edt_decompressor_out_158 , edt_decompressor_out_159 , edt_decompressor_out_160 ,
        edt_decompressor_out_161 , edt_decompressor_out_162 , edt_decompressor_out_163 , edt_decompressor_out_164 ,
        edt_decompressor_out_165 , edt_decompressor_out_166 , edt_decompressor_out_167 , edt_decompressor_out_168 ,
        edt_decompressor_out_169 , edt_decompressor_out_170 , edt_decompressor_out_171 , edt_decompressor_out_172 ,
        edt_decompressor_out_173 , edt_decompressor_out_174 , edt_decompressor_out_175 , edt_decompressor_out_176 ,
        edt_decompressor_out_177 , edt_decompressor_out_178 , edt_decompressor_out_179 , edt_decompressor_out_180 ,
        edt_decompressor_out_181 , edt_decompressor_out_182 , edt_decompressor_out_183 , edt_decompressor_out_184 ,
        edt_decompressor_out_185 , edt_decompressor_out_186 , edt_decompressor_out_187 , edt_decompressor_out_188 ,
        edt_decompressor_out_189 , edt_decompressor_out_190 , edt_decompressor_out_191 , edt_decompressor_out_192 ,
        edt_decompressor_out_193 , edt_decompressor_out_194 , edt_decompressor_out_195 , edt_decompressor_out_196 ,
        edt_decompressor_out_197 , edt_decompressor_out_198 , edt_decompressor_out_199 , edt_decompressor_out_200 ,
        edt_decompressor_out_201 , edt_decompressor_out_202 , edt_decompressor_out_203 , edt_decompressor_out_204 ,
        edt_decompressor_out_205 , edt_decompressor_out_206 , edt_decompressor_out_207 , edt_decompressor_out_208 ,
        edt_decompressor_out_209 , edt_decompressor_out_210 , edt_decompressor_out_211 , edt_decompressor_out_212 ,
        edt_decompressor_out_213 , edt_decompressor_out_214 , edt_decompressor_out_215 , edt_decompressor_out_216 ,
        edt_decompressor_out_217 , edt_decompressor_out_218 , edt_decompressor_out_219 , edt_decompressor_out_220 ,
        edt_decompressor_out_221 , edt_decompressor_out_222 , edt_decompressor_out_223 , edt_decompressor_out_224 ,
        edt_decompressor_out_225 , edt_decompressor_out_226 , edt_decompressor_out_227 , edt_decompressor_out_228 ,
        edt_decompressor_out_229 , edt_decompressor_out_230 , edt_decompressor_out_231 , edt_decompressor_out_232 ,
        edt_decompressor_out_233 , edt_decompressor_out_234 , edt_decompressor_out_235 , edt_decompressor_out_236 ,
        edt_decompressor_out_237 , edt_decompressor_out_238 , edt_decompressor_out_239 , edt_decompressor_out_240 ,
        edt_decompressor_out_241 , edt_decompressor_out_242 , edt_decompressor_out_243 , edt_decompressor_out_244 ,
        edt_decompressor_out_245 , edt_decompressor_out_246 , edt_decompressor_out_247 , edt_decompressor_out_248 ,
        edt_decompressor_out_249 , edt_decompressor_out_250 , edt_decompressor_out_251 , edt_decompressor_out_252 ,
        edt_decompressor_out_253 , edt_decompressor_out_254 , edt_decompressor_out_255 , edt_decompressor_out_256 ,
        edt_decompressor_out_257 , edt_decompressor_out_258 , edt_decompressor_out_259 , edt_decompressor_out_260 ,
        edt_decompressor_out_261 , edt_decompressor_out_262 , edt_decompressor_out_263 , edt_decompressor_out_264 ,
        edt_decompressor_out_265 , edt_decompressor_out_266 , edt_decompressor_out_267 , edt_decompressor_out_268 ,
        edt_decompressor_out_269 , edt_decompressor_out_270 , edt_decompressor_out_271 , edt_decompressor_out_272 ,
        edt_decompressor_out_273 , edt_decompressor_out_274 , edt_decompressor_out_275 , edt_decompressor_out_276 ,
        edt_decompressor_out_277 , edt_decompressor_out_278 , edt_decompressor_out_279 , edt_decompressor_out_280 ,
        edt_decompressor_out_281 , edt_decompressor_out_282 , edt_decompressor_out_283 , edt_decompressor_out_284 ,
        edt_decompressor_out_285 , edt_decompressor_out_286 , edt_decompressor_out_287 , edt_decompressor_out_288 ,
        edt_decompressor_out_289 , edt_decompressor_out_290 , edt_decompressor_out_291 , edt_decompressor_out_292 ,
        edt_decompressor_out_293 , edt_decompressor_out_294 , edt_decompressor_out_295 , edt_decompressor_out_296 ,
        edt_decompressor_out_297 , edt_decompressor_out_298 , edt_decompressor_out_299 , edt_decompressor_out_300 ,
        edt_decompressor_out_301 , edt_decompressor_out_302 , edt_decompressor_out_303 , edt_decompressor_out_304 ,
        edt_decompressor_out_305 , edt_decompressor_out_306 , edt_decompressor_out_307 , edt_decompressor_out_308 ,
        edt_decompressor_out_309 , edt_decompressor_out_310 , edt_decompressor_out_311 , edt_decompressor_out_312 ,
        edt_decompressor_out_313 , edt_decompressor_out_314 , edt_decompressor_out_315 , edt_decompressor_out_316 ,
        edt_decompressor_out_317 , edt_decompressor_out_318 , edt_decompressor_out_319 , edt_decompressor_out_320 ,
        edt_decompressor_out_321 , edt_decompressor_out_322 , edt_decompressor_out_323 , edt_decompressor_out_324 ,
        edt_decompressor_out_325 , edt_decompressor_out_326 , edt_decompressor_out_327 , edt_decompressor_out_328 ,
        edt_decompressor_out_329 , edt_decompressor_out_330 , edt_decompressor_out_331 , edt_decompressor_out_332 ,
        edt_decompressor_out_333 , edt_decompressor_out_334 , edt_decompressor_out_335 , edt_decompressor_out_336 ,
        edt_decompressor_out_337 , edt_decompressor_out_338 , edt_decompressor_out_339 , edt_decompressor_out_340 ,
        edt_decompressor_out_341 , edt_decompressor_out_342 , edt_decompressor_out_343 , edt_decompressor_out_344 ,
        edt_decompressor_out_345 , edt_decompressor_out_346 , edt_decompressor_out_347 , edt_decompressor_out_348 ,
        edt_decompressor_out_349 , edt_decompressor_out_350 , edt_decompressor_out_351 , edt_decompressor_out_352 ,
        edt_decompressor_out_353 , edt_decompressor_out_354 , edt_decompressor_out_355 , edt_decompressor_out_356 ,
        edt_decompressor_out_357 , edt_decompressor_out_358 , edt_decompressor_out_359 , edt_decompressor_out_360 ,
        edt_decompressor_out_361 , edt_decompressor_out_362 , edt_decompressor_out_363 , edt_decompressor_out_364 ,
        edt_decompressor_out_365 , edt_decompressor_out_366 , edt_decompressor_out_367 , edt_decompressor_out_368 ,
        edt_decompressor_out_369 , edt_decompressor_out_370 , edt_decompressor_out_371 , edt_decompressor_out_372 ,
        edt_decompressor_out_373 , edt_decompressor_out_374 , edt_decompressor_out_375 , edt_decompressor_out_376 ,
        edt_decompressor_out_377 , edt_decompressor_out_378 , edt_decompressor_out_379 , edt_decompressor_out_380 ,
        edt_decompressor_out_381 , edt_decompressor_out_382 , edt_decompressor_out_383 , edt_decompressor_out_384 ,
        edt_decompressor_out_385 , edt_decompressor_out_386 , edt_decompressor_out_387 , edt_decompressor_out_388 ,
        edt_decompressor_out_389 , edt_decompressor_out_390 , edt_decompressor_out_391 , edt_decompressor_out_392 ,
        edt_decompressor_out_393 , edt_decompressor_out_394 , edt_decompressor_out_395 , edt_decompressor_out_396 ,
        edt_decompressor_out_397 , edt_decompressor_out_398 , edt_decompressor_out_399 , edt_decompressor_out_400 ,
        edt_decompressor_out_401 , edt_decompressor_out_402 , edt_decompressor_out_403 , edt_decompressor_out_404 ,
        edt_decompressor_out_405 , edt_decompressor_out_406 , edt_decompressor_out_407 , edt_decompressor_out_408 ,
        edt_decompressor_out_409 , edt_decompressor_out_410 , edt_decompressor_out_411 , edt_decompressor_out_412 ,
        edt_decompressor_out_413 , edt_decompressor_out_414 , edt_decompressor_out_415 , edt_decompressor_out_416 ,
        edt_decompressor_out_417 , edt_decompressor_out_418 , edt_decompressor_out_419 , edt_decompressor_out_420 ,
        edt_decompressor_out_421 , edt_decompressor_out_422 , edt_decompressor_out_423 , edt_decompressor_out_424 ,
        edt_decompressor_out_425 , edt_decompressor_out_426 , edt_decompressor_out_427 , edt_decompressor_out_428 ,
        edt_decompressor_out_429 , edt_decompressor_out_430 , edt_decompressor_out_431 , edt_decompressor_out_432 ,
        edt_decompressor_out_433 , edt_decompressor_out_434 , edt_decompressor_out_435 , edt_decompressor_out_436 ,
        edt_decompressor_out_437 , edt_decompressor_out_438 , edt_decompressor_out_439 , edt_decompressor_out_440 ,
        edt_decompressor_out_441 , edt_decompressor_out_442 , edt_decompressor_out_443 , edt_decompressor_out_444 ,
        edt_decompressor_out_445 , edt_decompressor_out_446 , edt_decompressor_out_447 , edt_decompressor_out_448 ,
        edt_decompressor_out_449 , edt_decompressor_out_450 , edt_decompressor_out_451 , edt_decompressor_out_452 ,
        edt_decompressor_out_453 , edt_decompressor_out_454 , edt_decompressor_out_455 , edt_decompressor_out_456 ,
        edt_decompressor_out_457 , edt_decompressor_out_458 , edt_decompressor_out_459 , edt_decompressor_out_460 ,
        edt_decompressor_out_461 , edt_decompressor_out_462 , edt_decompressor_out_463 , edt_decompressor_out_464 ,
        edt_decompressor_out_465 , edt_decompressor_out_466 , edt_decompressor_out_467 , edt_decompressor_out_468 ,
        edt_decompressor_out_469 , edt_decompressor_out_470 , edt_decompressor_out_471 , edt_decompressor_out_472 ,
        edt_decompressor_out_473 , edt_decompressor_out_474 , edt_decompressor_out_475 , edt_decompressor_out_476 ,
        edt_decompressor_out_477 , edt_decompressor_out_478 , edt_decompressor_out_479 , edt_decompressor_out_480 ,
        edt_decompressor_out_481 , edt_decompressor_out_482 , edt_decompressor_out_483 , edt_decompressor_out_484 ,
        edt_decompressor_out_485 , edt_decompressor_out_486 , edt_decompressor_out_487 , edt_decompressor_out_488 ,
        edt_decompressor_out_489 , edt_decompressor_out_490 , edt_decompressor_out_491 , edt_decompressor_out_492 ,
        edt_decompressor_out_493 , edt_decompressor_out_494 , edt_decompressor_out_495 , edt_decompressor_out_496 ,
        edt_decompressor_out_497 , edt_decompressor_out_498 , edt_decompressor_out_499 , edt_decompressor_out_500 ,
        edt_decompressor_out_501 , edt_decompressor_out_502 , edt_decompressor_out_503 , edt_decompressor_out_504 ,
        edt_decompressor_out_505 , edt_decompressor_out_506 , edt_decompressor_out_507 , edt_decompressor_out_508 ,
        edt_decompressor_out_509 , edt_decompressor_out_510 , edt_decompressor_out_511 , edt_decompressor_out_512 ,
        edt_decompressor_out_513 , edt_decompressor_out_514 , edt_decompressor_out_515 , edt_decompressor_out_516 ,
        edt_decompressor_out_517 , edt_decompressor_out_518 , edt_decompressor_out_519 , edt_decompressor_out_520 ,
        edt_decompressor_out_521 , edt_decompressor_out_522 , edt_decompressor_out_523 , edt_decompressor_out_524 ,
        edt_decompressor_out_525 , edt_decompressor_out_526 , edt_decompressor_out_527 , edt_decompressor_out_528 ,
        edt_decompressor_out_529 , edt_decompressor_out_530 , edt_decompressor_out_531 , edt_decompressor_out_532 ,
        edt_decompressor_out_533 , edt_decompressor_out_534 , edt_decompressor_out_535 , edt_decompressor_out_536 ,
        edt_decompressor_out_537 , edt_decompressor_out_538 , edt_decompressor_out_539 , edt_decompressor_out_540 ,
        edt_decompressor_out_541 , edt_decompressor_out_542 , edt_decompressor_out_543 , edt_decompressor_out_544 ,
        edt_decompressor_out_545 , edt_decompressor_out_546 , edt_decompressor_out_547 , edt_decompressor_out_548 ,
        edt_decompressor_out_549 , edt_decompressor_out_550 , edt_decompressor_out_551 , edt_decompressor_out_552 ,
        edt_decompressor_out_553 , edt_decompressor_out_554 , edt_decompressor_out_555 , edt_decompressor_out_556 ,
        edt_decompressor_out_557 , edt_decompressor_out_558 , edt_decompressor_out_559 , edt_decompressor_out_560 ,
        edt_decompressor_out_561 , edt_decompressor_out_562 , edt_decompressor_out_563 , edt_decompressor_out_564 ,
        edt_decompressor_out_565 , edt_decompressor_out_566 , edt_decompressor_out_567 , edt_decompressor_out_568 ,
        edt_decompressor_out_569 , edt_decompressor_out_570 , edt_decompressor_out_571 , edt_decompressor_out_572 ,
        edt_decompressor_out_573 , edt_decompressor_out_574 , edt_decompressor_out_575 , edt_decompressor_out_576 ,
        edt_decompressor_out_577 , edt_decompressor_out_578 , edt_decompressor_out_579 , edt_decompressor_out_580 ,
        edt_decompressor_out_581 , edt_decompressor_out_582 , edt_decompressor_out_583 , edt_decompressor_out_584 ,
        edt_decompressor_out_585 , edt_decompressor_out_586 , edt_decompressor_out_587 , edt_decompressor_out_588 ,
        edt_decompressor_out_589 , edt_decompressor_out_590 , edt_decompressor_out_591 , edt_decompressor_out_592 ,
        edt_decompressor_out_593 , edt_decompressor_out_594 , edt_decompressor_out_595 , edt_decompressor_out_596 ,
        edt_decompressor_out_597 , edt_decompressor_out_598 , edt_decompressor_out_599 , edt_decompressor_out_600 ,
        edt_decompressor_out_601 , edt_decompressor_out_602 , edt_decompressor_out_603 , edt_decompressor_out_604 ,
        edt_decompressor_out_605 , edt_decompressor_out_606 , edt_decompressor_out_607 , edt_decompressor_out_608 ,
        edt_decompressor_out_609 , edt_decompressor_out_610 , edt_decompressor_out_611 , edt_decompressor_out_612 ,
        edt_decompressor_out_613 , edt_decompressor_out_614 , edt_decompressor_out_615 , edt_decompressor_out_616 ,
        edt_decompressor_out_617 , edt_decompressor_out_618 , edt_decompressor_out_619 , edt_decompressor_out_620 ,
        edt_decompressor_out_621 , edt_decompressor_out_622 , edt_decompressor_out_623 , edt_decompressor_out_624 ,
        edt_decompressor_out_625 , edt_decompressor_out_626 , edt_decompressor_out_627 , edt_decompressor_out_628 ,
        edt_decompressor_out_629 , edt_decompressor_out_630 , edt_decompressor_out_631 , edt_decompressor_out_632 ,
        edt_decompressor_out_633 , edt_decompressor_out_634 , edt_decompressor_out_635 , edt_decompressor_out_636 ,
        edt_decompressor_out_637 , edt_decompressor_out_638 , edt_decompressor_out_639 , edt_decompressor_out_640 ,
        edt_decompressor_out_641 , edt_decompressor_out_642 , edt_decompressor_out_643 , edt_decompressor_out_644 ,
        edt_decompressor_out_645 , edt_decompressor_out_646 , edt_decompressor_out_647 , edt_decompressor_out_648 ,
        edt_decompressor_out_649 , edt_decompressor_out_650 , edt_decompressor_out_651 , edt_decompressor_out_652 ,
        edt_decompressor_out_653 , edt_decompressor_out_654 , edt_decompressor_out_655 , edt_decompressor_out_656 ,
        edt_decompressor_out_657 , edt_decompressor_out_658 , edt_decompressor_out_659 , edt_decompressor_out_660 ,
        edt_decompressor_out_661 , edt_decompressor_out_662 , edt_decompressor_out_663 , edt_decompressor_out_664 ,
        edt_decompressor_out_665 , edt_decompressor_out_666 , edt_decompressor_out_667 , edt_decompressor_out_668 ,
        edt_decompressor_out_669 , edt_decompressor_out_670 , edt_decompressor_out_671 , edt_decompressor_out_672 ,
        edt_decompressor_out_673 , edt_decompressor_out_674 , edt_decompressor_out_675 , edt_decompressor_out_676 ,
        edt_decompressor_out_677 , edt_decompressor_out_678 , edt_decompressor_out_679 , edt_decompressor_out_680 ,
        edt_decompressor_out_681 , edt_decompressor_out_682 , edt_decompressor_out_683 , edt_decompressor_out_684 ,
        edt_decompressor_out_685 , edt_decompressor_out_686 , edt_decompressor_out_687 , edt_decompressor_out_688 ,
        edt_decompressor_out_689 , edt_decompressor_out_690 , edt_decompressor_out_691 , edt_decompressor_out_692 ,
        edt_decompressor_out_693 , edt_decompressor_out_694 , edt_decompressor_out_695 , edt_decompressor_out_696 ,
        edt_decompressor_out_697 , edt_decompressor_out_698 , edt_decompressor_out_699 , edt_decompressor_out_700 ,
        edt_decompressor_out_701 , edt_decompressor_out_702 , edt_decompressor_out_703 , edt_decompressor_out_704 ,
        edt_decompressor_out_705 , edt_decompressor_out_706 , edt_decompressor_out_707 , edt_decompressor_out_708 ,
        edt_decompressor_out_709 , edt_decompressor_out_710 , edt_decompressor_out_711 , edt_decompressor_out_712 ,
        edt_decompressor_out_713 , edt_decompressor_out_714 , edt_decompressor_out_715 , edt_decompressor_out_716 ,
        edt_decompressor_out_717 , edt_decompressor_out_718 , edt_decompressor_out_719 , edt_decompressor_out_720 ,
        edt_decompressor_out_721 , edt_decompressor_out_722 , edt_decompressor_out_723 , edt_decompressor_out_724 ,
        edt_decompressor_out_725 , edt_decompressor_out_726 , edt_decompressor_out_727 , edt_decompressor_out_728 ,
        edt_decompressor_out_729 , edt_decompressor_out_730 , edt_decompressor_out_731 , edt_decompressor_out_732 ,
        edt_decompressor_out_733 , edt_decompressor_out_734 , edt_decompressor_out_735 , edt_decompressor_out_736 ,
        edt_decompressor_out_737 , edt_decompressor_out_738 , edt_decompressor_out_739 , edt_decompressor_out_740 ,
        edt_decompressor_out_741 , edt_decompressor_out_742 , edt_decompressor_out_743 , edt_decompressor_out_744 ,
        edt_decompressor_out_745 , edt_decompressor_out_746 , edt_decompressor_out_747 , edt_decompressor_out_748 ,
        edt_decompressor_out_749 , edt_decompressor_out_750 , edt_decompressor_out_751 , edt_decompressor_out_752 ,
        edt_decompressor_out_753 , edt_decompressor_out_754 , edt_decompressor_out_755 , edt_decompressor_out_756 ,
        edt_decompressor_out_757 , edt_decompressor_out_758 , edt_decompressor_out_759 , edt_decompressor_out_760 ,
        edt_decompressor_out_761 , edt_decompressor_out_762 , edt_decompressor_out_763 , edt_decompressor_out_764 ,
        edt_decompressor_out_765 , edt_decompressor_out_766 , edt_decompressor_out_767 , edt_decompressor_out_768 ,
        edt_decompressor_out_769 , edt_decompressor_out_770 , edt_decompressor_out_771 , edt_decompressor_out_772 ,
        edt_decompressor_out_773 , edt_decompressor_out_774 , edt_decompressor_out_775 , edt_decompressor_out_776 ,
        edt_decompressor_out_777 , edt_decompressor_out_778 , edt_decompressor_out_779 , edt_decompressor_out_780 ,
        edt_decompressor_out_781 , edt_decompressor_out_782 , edt_decompressor_out_783 , edt_decompressor_out_784 ,
        edt_decompressor_out_785 , edt_decompressor_out_786 , edt_decompressor_out_787 , edt_decompressor_out_788 ,
        edt_decompressor_out_789 , edt_decompressor_out_790 , edt_decompressor_out_791 , edt_decompressor_out_792 ,
        edt_decompressor_out_793 , edt_decompressor_out_794 , edt_decompressor_out_795 , edt_update_hfs_netlink_29280 ,
        edt_update_hfs_netlink_29281 , edt_update_hfs_netlink_29282 , edt_update_hfs_netlink_29283 , edt_update_hfs_netlink_29284 ,
        edt_update_hfs_netlink_29285 , edt_update_hfs_netlink_29286 , edt_update_hfs_netlink_29287 , edt_update_hfs_netlink_29288 ,
        edt_update_hfs_netlink_29289 , edt_configuration_hfs_netlink_29290 , edt_configuration_hfs_netlink_29291 , edt_configuration_hfs_netlink_29292 ,
        edt_clock_cts_1 , edt_clock_cts_2 , edt_clock_cts_3 , edt_clock_cts_4 ,
        edt_clock_cts_5 , edt_clock_cts_6 , edt_clock_cts_7 , edt_clock_cts_8 ,
        edt_clock_cts_9 , edt_clock_cts_0_1 , edt_clock_cts_1_1 , edt_clock_cts_2_1 ,
        edt_clock_cts_3_1 , edt_clock_cts_4_1 , edt_clock_cts_5_1 , edt_clock_cts_6_1 , GND,
        edt_clock_cts_7_1 ;
wire    masks_hold_reg_10_0 , masks_hold_reg_10_1 , masks_hold_reg_10_2 , masks_hold_reg_10_3 ,
        masks_hold_reg_10_4 , masks_hold_reg_10_5 , masks_hold_reg_10_6 , masks_hold_reg_10_7 ,
        masks_hold_reg_10_8 , masks_hold_reg_10_9 , masks_hold_reg_10_10 , config0_onehot_decoded_masks_11_0 ,
        config0_onehot_decoded_masks_11_1 , config0_onehot_decoded_masks_11_2 , config0_onehot_decoded_masks_11_3 , config0_onehot_decoded_masks_11_4 ,
        config0_onehot_decoded_masks_11_5 , config0_onehot_decoded_masks_11_6 , config0_onehot_decoded_masks_11_7 , config0_onehot_decoded_masks_11_8 ,
        config0_onehot_decoded_masks_11_9 , config0_onehot_decoded_masks_11_10 , config0_onehot_decoded_masks_11_11 , config0_onehot_decoded_masks_11_12 ,
        config0_onehot_decoded_masks_11_13 , config0_onehot_decoded_masks_11_14 , config0_onehot_decoded_masks_11_15 , config0_onehot_decoded_masks_11_16 ,
        config0_onehot_decoded_masks_11_17 , config0_onehot_decoded_masks_11_18 , config0_onehot_decoded_masks_11_19 , config0_onehot_decoded_masks_11_20 ,
        config0_onehot_decoded_masks_11_21 , config0_onehot_decoded_masks_11_22 , config0_onehot_decoded_masks_11_23 , config0_onehot_decoded_masks_11_24 ,
        config0_onehot_decoded_masks_11_25 , config0_onehot_decoded_masks_11_26 , config0_onehot_decoded_masks_11_27 , config0_onehot_decoded_masks_11_28 ,
        config0_onehot_decoded_masks_11_29 , config0_onehot_decoded_masks_11_30 , config0_onehot_decoded_masks_11_31 , config0_onehot_decoded_masks_11_32 ,
        config0_onehot_decoded_masks_11_33 , config0_onehot_decoded_masks_11_34 , config0_onehot_decoded_masks_11_35 , config0_onehot_decoded_masks_11_36 ,
        config0_onehot_decoded_masks_11_37 , config0_onehot_decoded_masks_11_38 , config0_onehot_decoded_masks_11_39 , config0_onehot_decoded_masks_11_40 ,
        config0_onehot_decoded_masks_11_41 , config0_onehot_decoded_masks_11_42 , config0_onehot_decoded_masks_11_43 , config0_onehot_decoded_masks_11_44 ,
        config0_onehot_decoded_masks_11_45 , config0_onehot_decoded_masks_11_46 , config0_onehot_decoded_masks_11_47 , config0_onehot_decoded_masks_11_48 ,
        config0_onehot_decoded_masks_11_49 , config0_onehot_decoded_masks_11_50 , config0_onehot_decoded_masks_11_51 , config0_onehot_decoded_masks_11_52 ,
        masks_hold_reg_11_0 , masks_hold_reg_11_1 , masks_hold_reg_11_2 , masks_hold_reg_11_3 ,
        masks_hold_reg_11_4 , masks_hold_reg_11_5 , masks_hold_reg_11_6 , masks_hold_reg_11_7 ,
        masks_hold_reg_11_8 , masks_hold_reg_11_9 , masks_hold_reg_11_10 , config0_onehot_decoded_masks_12_0 ,
        config0_onehot_decoded_masks_12_1 , config0_onehot_decoded_masks_12_2 , config0_onehot_decoded_masks_12_3 , config0_onehot_decoded_masks_12_4 ,
        config0_onehot_decoded_masks_12_5 , config0_onehot_decoded_masks_12_6 , config0_onehot_decoded_masks_12_7 , config0_onehot_decoded_masks_12_8 ,
        config0_onehot_decoded_masks_12_9 , config0_onehot_decoded_masks_12_10 , config0_onehot_decoded_masks_12_11 , config0_onehot_decoded_masks_12_12 ,
        config0_onehot_decoded_masks_12_13 , config0_onehot_decoded_masks_12_14 , config0_onehot_decoded_masks_12_15 , config0_onehot_decoded_masks_12_16 ,
        config0_onehot_decoded_masks_12_17 , config0_onehot_decoded_masks_12_18 , config0_onehot_decoded_masks_12_19 , config0_onehot_decoded_masks_12_20 ,
        config0_onehot_decoded_masks_12_21 , config0_onehot_decoded_masks_12_22 , config0_onehot_decoded_masks_12_23 , config0_onehot_decoded_masks_12_24 ,
        config0_onehot_decoded_masks_12_25 , config0_onehot_decoded_masks_12_26 , config0_onehot_decoded_masks_12_27 , config0_onehot_decoded_masks_12_28 ,
        config0_onehot_decoded_masks_12_29 , config0_onehot_decoded_masks_12_30 , config0_onehot_decoded_masks_12_31 , config0_onehot_decoded_masks_12_32 ,
        config0_onehot_decoded_masks_12_33 , config0_onehot_decoded_masks_12_34 , config0_onehot_decoded_masks_12_35 , config0_onehot_decoded_masks_12_36 ,
        config0_onehot_decoded_masks_12_37 , config0_onehot_decoded_masks_12_38 , config0_onehot_decoded_masks_12_39 , config0_onehot_decoded_masks_12_40 ,
        config0_onehot_decoded_masks_12_41 , config0_onehot_decoded_masks_12_42 , config0_onehot_decoded_masks_12_43 , config0_onehot_decoded_masks_12_44 ,
        config0_onehot_decoded_masks_12_45 , config0_onehot_decoded_masks_12_46 , config0_onehot_decoded_masks_12_47 , config0_onehot_decoded_masks_12_48 ,
        config0_onehot_decoded_masks_12_49 , config0_onehot_decoded_masks_12_50 , config0_onehot_decoded_masks_12_51 , config0_onehot_decoded_masks_12_52 ,
        masks_hold_reg_8_0 , masks_hold_reg_8_1 , masks_hold_reg_8_2 , masks_hold_reg_8_3 ,
        masks_hold_reg_8_4 , masks_hold_reg_8_5 , masks_hold_reg_8_6 , masks_hold_reg_8_7 ,
        masks_hold_reg_8_8 , masks_hold_reg_8_9 , masks_hold_reg_8_10 , config0_onehot_decoded_masks_9_0 ,
        config0_onehot_decoded_masks_9_1 , config0_onehot_decoded_masks_9_2 , config0_onehot_decoded_masks_9_3 , config0_onehot_decoded_masks_9_4 ,
        config0_onehot_decoded_masks_9_5 , config0_onehot_decoded_masks_9_6 , config0_onehot_decoded_masks_9_7 , config0_onehot_decoded_masks_9_8 ,
        config0_onehot_decoded_masks_9_9 , config0_onehot_decoded_masks_9_10 , config0_onehot_decoded_masks_9_11 , config0_onehot_decoded_masks_9_12 ,
        config0_onehot_decoded_masks_9_13 , config0_onehot_decoded_masks_9_14 , config0_onehot_decoded_masks_9_15 , config0_onehot_decoded_masks_9_16 ,
        config0_onehot_decoded_masks_9_17 , config0_onehot_decoded_masks_9_18 , config0_onehot_decoded_masks_9_19 , config0_onehot_decoded_masks_9_20 ,
        config0_onehot_decoded_masks_9_21 , config0_onehot_decoded_masks_9_22 , config0_onehot_decoded_masks_9_23 , config0_onehot_decoded_masks_9_24 ,
        config0_onehot_decoded_masks_9_25 , config0_onehot_decoded_masks_9_26 , config0_onehot_decoded_masks_9_27 , config0_onehot_decoded_masks_9_28 ,
        config0_onehot_decoded_masks_9_29 , config0_onehot_decoded_masks_9_30 , config0_onehot_decoded_masks_9_31 , config0_onehot_decoded_masks_9_32 ,
        config0_onehot_decoded_masks_9_33 , config0_onehot_decoded_masks_9_34 , config0_onehot_decoded_masks_9_35 , config0_onehot_decoded_masks_9_36 ,
        config0_onehot_decoded_masks_9_37 , config0_onehot_decoded_masks_9_38 , config0_onehot_decoded_masks_9_39 , config0_onehot_decoded_masks_9_40 ,
        config0_onehot_decoded_masks_9_41 , config0_onehot_decoded_masks_9_42 , config0_onehot_decoded_masks_9_43 , config0_onehot_decoded_masks_9_44 ,
        config0_onehot_decoded_masks_9_45 , config0_onehot_decoded_masks_9_46 , config0_onehot_decoded_masks_9_47 , config0_onehot_decoded_masks_9_48 ,
        config0_onehot_decoded_masks_9_49 , config0_onehot_decoded_masks_9_50 , config0_onehot_decoded_masks_9_51 , config0_onehot_decoded_masks_9_52 ,
        masks_hold_reg_9_0 , masks_hold_reg_9_1 , masks_hold_reg_9_2 , masks_hold_reg_9_3 ,
        masks_hold_reg_9_4 , masks_hold_reg_9_5 , masks_hold_reg_9_6 , masks_hold_reg_9_7 ,
        masks_hold_reg_9_8 , masks_hold_reg_9_9 , masks_hold_reg_9_10 , config0_onehot_decoded_masks_10_0 ,
        config0_onehot_decoded_masks_10_1 , config0_onehot_decoded_masks_10_2 , config0_onehot_decoded_masks_10_3 , config0_onehot_decoded_masks_10_4 ,
        config0_onehot_decoded_masks_10_5 , config0_onehot_decoded_masks_10_6 , config0_onehot_decoded_masks_10_7 , config0_onehot_decoded_masks_10_8 ,
        config0_onehot_decoded_masks_10_9 , config0_onehot_decoded_masks_10_10 , config0_onehot_decoded_masks_10_11 , config0_onehot_decoded_masks_10_12 ,
        config0_onehot_decoded_masks_10_13 , config0_onehot_decoded_masks_10_14 , config0_onehot_decoded_masks_10_15 , config0_onehot_decoded_masks_10_16 ,
        config0_onehot_decoded_masks_10_17 , config0_onehot_decoded_masks_10_18 , config0_onehot_decoded_masks_10_19 , config0_onehot_decoded_masks_10_20 ,
        config0_onehot_decoded_masks_10_21 , config0_onehot_decoded_masks_10_22 , config0_onehot_decoded_masks_10_23 , config0_onehot_decoded_masks_10_24 ,
        config0_onehot_decoded_masks_10_25 , config0_onehot_decoded_masks_10_26 , config0_onehot_decoded_masks_10_27 , config0_onehot_decoded_masks_10_28 ,
        config0_onehot_decoded_masks_10_29 , config0_onehot_decoded_masks_10_30 , config0_onehot_decoded_masks_10_31 , config0_onehot_decoded_masks_10_32 ,
        config0_onehot_decoded_masks_10_33 , config0_onehot_decoded_masks_10_34 , config0_onehot_decoded_masks_10_35 , config0_onehot_decoded_masks_10_36 ,
        config0_onehot_decoded_masks_10_37 , config0_onehot_decoded_masks_10_38 , config0_onehot_decoded_masks_10_39 , config0_onehot_decoded_masks_10_40 ,
        config0_onehot_decoded_masks_10_41 , config0_onehot_decoded_masks_10_42 , config0_onehot_decoded_masks_10_43 , config0_onehot_decoded_masks_10_44 ,
        config0_onehot_decoded_masks_10_45 , config0_onehot_decoded_masks_10_46 , config0_onehot_decoded_masks_10_47 , config0_onehot_decoded_masks_10_48 ,
        config0_onehot_decoded_masks_10_49 , config0_onehot_decoded_masks_10_50 , config0_onehot_decoded_masks_10_51 , config0_onehot_decoded_masks_10_52 ,
        masks_hold_reg_12_0 , masks_hold_reg_12_1 , masks_hold_reg_12_2 , masks_hold_reg_12_3 ,
        masks_hold_reg_12_4 , masks_hold_reg_12_5 , masks_hold_reg_12_6 , masks_hold_reg_12_7 ,
        masks_hold_reg_12_8 , masks_hold_reg_12_9 , masks_hold_reg_12_10 , config0_onehot_decoded_masks_13_0 ,
        config0_onehot_decoded_masks_13_1 , config0_onehot_decoded_masks_13_2 , config0_onehot_decoded_masks_13_3 , config0_onehot_decoded_masks_13_4 ,
        config0_onehot_decoded_masks_13_5 , config0_onehot_decoded_masks_13_6 , config0_onehot_decoded_masks_13_7 , config0_onehot_decoded_masks_13_8 ,
        config0_onehot_decoded_masks_13_9 , config0_onehot_decoded_masks_13_10 , config0_onehot_decoded_masks_13_11 , config0_onehot_decoded_masks_13_12 ,
        config0_onehot_decoded_masks_13_13 , config0_onehot_decoded_masks_13_14 , config0_onehot_decoded_masks_13_15 , config0_onehot_decoded_masks_13_16 ,
        config0_onehot_decoded_masks_13_17 , config0_onehot_decoded_masks_13_18 , config0_onehot_decoded_masks_13_19 , config0_onehot_decoded_masks_13_20 ,
        config0_onehot_decoded_masks_13_21 , config0_onehot_decoded_masks_13_22 , config0_onehot_decoded_masks_13_23 , config0_onehot_decoded_masks_13_24 ,
        config0_onehot_decoded_masks_13_25 , config0_onehot_decoded_masks_13_26 , config0_onehot_decoded_masks_13_27 , config0_onehot_decoded_masks_13_28 ,
        config0_onehot_decoded_masks_13_29 , config0_onehot_decoded_masks_13_30 , config0_onehot_decoded_masks_13_31 , config0_onehot_decoded_masks_13_32 ,
        config0_onehot_decoded_masks_13_33 , config0_onehot_decoded_masks_13_34 , config0_onehot_decoded_masks_13_35 , config0_onehot_decoded_masks_13_36 ,
        config0_onehot_decoded_masks_13_37 , config0_onehot_decoded_masks_13_38 , config0_onehot_decoded_masks_13_39 , config0_onehot_decoded_masks_13_40 ,
        config0_onehot_decoded_masks_13_41 , config0_onehot_decoded_masks_13_42 , config0_onehot_decoded_masks_13_43 , config0_onehot_decoded_masks_13_44 ,
        config0_onehot_decoded_masks_13_45 , config0_onehot_decoded_masks_13_46 , config0_onehot_decoded_masks_13_47 , config0_onehot_decoded_masks_13_48 ,
        config0_onehot_decoded_masks_13_49 , config0_onehot_decoded_masks_13_50 , config0_onehot_decoded_masks_13_51 , config0_onehot_decoded_masks_13_52 ,
        masks_hold_reg_13_0 , masks_hold_reg_13_1 , masks_hold_reg_13_2 , masks_hold_reg_13_3 ,
        masks_hold_reg_13_4 , masks_hold_reg_13_5 , masks_hold_reg_13_6 , masks_hold_reg_13_7 ,
        config0_onehot_decoded_masks_14_0 , config0_onehot_decoded_masks_14_1 , config0_onehot_decoded_masks_14_2 , config0_onehot_decoded_masks_14_3 ,
        config0_onehot_decoded_masks_14_4 , config0_onehot_decoded_masks_14_5 , config0_onehot_decoded_masks_14_6 , config0_onehot_decoded_masks_14_7 ,
        config0_onehot_decoded_masks_14_8 , config0_onehot_decoded_masks_14_9 , config0_onehot_decoded_masks_14_10 , config0_onehot_decoded_masks_14_11 ,
        config0_onehot_decoded_masks_14_12 , config0_onehot_decoded_masks_14_13 , config0_onehot_decoded_masks_14_14 , config0_onehot_decoded_masks_14_15 ,
        config0_onehot_decoded_masks_14_16 , config0_onehot_decoded_masks_14_17 , config0_onehot_decoded_masks_14_18 , config0_onehot_decoded_masks_14_19 ,
        config0_onehot_decoded_masks_14_20 , config0_onehot_decoded_masks_14_21 , config0_onehot_decoded_masks_14_22 , config0_onehot_decoded_masks_14_23 ,
        config0_onehot_decoded_masks_14_24 , config0_onehot_decoded_masks_14_25 , config0_onehot_decoded_masks_14_26 , config0_onehot_decoded_masks_14_27 ,
        config0_onehot_decoded_masks_14_28 , config0_onehot_decoded_masks_14_29 , config0_onehot_decoded_masks_14_30 , config0_onehot_decoded_masks_14_31 ,
        config0_onehot_decoded_masks_14_32 , config0_onehot_decoded_masks_14_33 , config0_onehot_decoded_masks_14_34 , config0_onehot_decoded_masks_14_35 ,
        config0_onehot_decoded_masks_14_36 , config0_onehot_decoded_masks_14_37 , config0_onehot_decoded_masks_14_38 , config0_onehot_decoded_masks_14_39 ,
        config0_onehot_decoded_masks_14_40 , config0_onehot_decoded_masks_14_41 , config0_onehot_decoded_masks_14_42 , config0_onehot_decoded_masks_14_43 ,
        config0_onehot_decoded_masks_14_44 , config0_onehot_decoded_masks_14_45 , config0_onehot_decoded_masks_14_46 , config0_onehot_decoded_masks_14_47 ,
        config0_onehot_decoded_masks_14_48 , config0_onehot_decoded_masks_14_49 , config0_onehot_decoded_masks_14_50 , config0_onehot_decoded_masks_14_51 ,
        config0_onehot_decoded_masks_14_52 , masks_hold_reg_7_0 , masks_hold_reg_7_1 , masks_hold_reg_7_2 ,
        masks_hold_reg_7_3 , masks_hold_reg_7_4 , masks_hold_reg_7_5 , masks_hold_reg_7_6 ,
        masks_hold_reg_7_7 , masks_hold_reg_7_8 , masks_hold_reg_7_9 , masks_hold_reg_7_10 ,
        masks_hold_reg_6_0 , masks_hold_reg_6_1 , masks_hold_reg_6_2 , masks_hold_reg_6_3 ,
        masks_hold_reg_6_4 , masks_hold_reg_6_5 , masks_hold_reg_6_6 , masks_hold_reg_6_7 ,
        masks_hold_reg_6_8 , masks_hold_reg_6_9 , masks_hold_reg_6_10 , masks_hold_reg_4_0 ,
        masks_hold_reg_4_1 , masks_hold_reg_4_2 , masks_hold_reg_4_3 , masks_hold_reg_4_4 ,
        masks_hold_reg_4_5 , masks_hold_reg_4_6 , masks_hold_reg_4_7 , masks_hold_reg_4_8 ,
        masks_hold_reg_4_9 , masks_hold_reg_4_10 , masks_hold_reg_5_0 , masks_hold_reg_5_1 ,
        masks_hold_reg_5_2 , masks_hold_reg_5_3 , masks_hold_reg_5_4 , masks_hold_reg_5_5 ,
        masks_hold_reg_5_6 , masks_hold_reg_5_7 , masks_hold_reg_5_8 , masks_hold_reg_5_9 ,
        masks_hold_reg_5_10 , masks_hold_reg_2_0 , masks_hold_reg_2_1 , masks_hold_reg_2_2 ,
        masks_hold_reg_2_3 , masks_hold_reg_2_4 , masks_hold_reg_2_5 , masks_hold_reg_2_6 ,
        masks_hold_reg_2_7 , masks_hold_reg_2_8 , masks_hold_reg_2_9 , masks_hold_reg_2_10 ,
        masks_hold_reg_3_0 , masks_hold_reg_3_1 , masks_hold_reg_3_2 , masks_hold_reg_3_3 ,
        masks_hold_reg_3_4 , masks_hold_reg_3_5 , masks_hold_reg_3_6 , masks_hold_reg_3_7 ,
        masks_hold_reg_3_8 , masks_hold_reg_3_9 , masks_hold_reg_3_10 , masks_hold_reg_1_0 ,
        masks_hold_reg_1_1 , masks_hold_reg_1_2 , masks_hold_reg_1_3 , masks_hold_reg_1_4 ,
        masks_hold_reg_1_5 , masks_hold_reg_1_6 , masks_hold_reg_1_7 , masks_hold_reg_1_8 ,
        masks_hold_reg_1_9 , masks_hold_reg_1_10 , masks_hold_reg_0_0 , masks_hold_reg_0_1 ,
        masks_hold_reg_0_2 , masks_hold_reg_0_3 , masks_hold_reg_0_4 , masks_hold_reg_0_5 ,
        masks_hold_reg_0_6 , masks_hold_reg_0_7 , masks_hold_reg_0_8 , masks_hold_reg_0_9 ,
        config1_xor_encoded_masks_0 , config1_xor_encoded_masks_1 , config1_xor_encoded_masks_2 , config1_xor_encoded_masks_3 ,
        config1_xor_encoded_masks_4 , config1_xor_encoded_masks_5 , config1_xor_encoded_masks_6 , config1_xor_encoded_masks_7 ,
        config1_xor_encoded_masks_8 , config1_xor_encoded_masks_9 , config1_xor_encoded_masks_10 , config1_xor_encoded_masks_11 ,
        config1_xor_encoded_masks_12 , config1_xor_encoded_masks_13 , config1_xor_encoded_masks_14 , config1_xor_encoded_masks_15 ,
        config1_xor_encoded_masks_16 , config1_xor_encoded_masks_17 , config1_xor_encoded_masks_18 , config1_xor_encoded_masks_19 ,
        config1_xor_encoded_masks_20 , config1_xor_encoded_masks_21 , config1_xor_encoded_masks_22 , config1_xor_encoded_masks_23 ,
        config1_xor_encoded_masks_24 , config1_xor_encoded_masks_25 , config1_xor_encoded_masks_26 , config1_xor_encoded_masks_27 ,
        config1_xor_encoded_masks_28 , config1_xor_encoded_masks_29 , config1_xor_encoded_masks_30 , config1_xor_encoded_masks_31 ,
        config1_xor_encoded_masks_32 , config1_xor_encoded_masks_33 , config1_xor_encoded_masks_34 , config1_xor_encoded_masks_35 ,
        config1_xor_encoded_masks_36 , config1_xor_encoded_masks_37 , config1_xor_encoded_masks_38 , config1_xor_encoded_masks_39 ,
        config1_xor_encoded_masks_40 , config1_xor_encoded_masks_41 , config1_xor_encoded_masks_42 , config1_xor_encoded_masks_43 ,
        config1_xor_encoded_masks_44 , config1_xor_encoded_masks_45 , config1_xor_encoded_masks_46 , config1_xor_encoded_masks_47 ,
        config1_xor_encoded_masks_48 , config1_xor_encoded_masks_49 , config1_xor_encoded_masks_50 , config1_xor_encoded_masks_51 ,
        config1_xor_encoded_masks_52 , config1_xor_encoded_masks_53 , config1_xor_encoded_masks_54 , config1_xor_encoded_masks_55 ,
        config1_xor_encoded_masks_56 , config1_xor_encoded_masks_57 , config1_xor_encoded_masks_58 , config1_xor_encoded_masks_59 ,
        config1_xor_encoded_masks_60 , config1_xor_encoded_masks_61 , config1_xor_encoded_masks_62 , config1_xor_encoded_masks_63 ,
        config1_xor_encoded_masks_64 , config1_xor_encoded_masks_65 , config1_xor_encoded_masks_66 , config1_xor_encoded_masks_67 ,
        config1_xor_encoded_masks_68 , config1_xor_encoded_masks_69 , config1_xor_encoded_masks_70 , config1_xor_encoded_masks_71 ,
        config1_xor_encoded_masks_72 , config1_xor_encoded_masks_73 , config1_xor_encoded_masks_74 , config1_xor_encoded_masks_75 ,
        config1_xor_encoded_masks_76 , config1_xor_encoded_masks_77 , config1_xor_encoded_masks_78 , config1_xor_encoded_masks_79 ,
        config1_xor_encoded_masks_80 , config1_xor_encoded_masks_81 , config1_xor_encoded_masks_82 , config1_xor_encoded_masks_83 ,
        config1_xor_encoded_masks_84 , config1_xor_encoded_masks_85 , config1_xor_encoded_masks_86 , config1_xor_encoded_masks_87 ,
        config1_xor_encoded_masks_88 , config1_xor_encoded_masks_89 , config1_xor_encoded_masks_90 , config1_xor_encoded_masks_91 ,
        config1_xor_encoded_masks_92 , config1_xor_encoded_masks_93 , config1_xor_encoded_masks_94 , config1_xor_encoded_masks_95 ,
        config1_xor_encoded_masks_96 , config1_xor_encoded_masks_97 , config1_xor_encoded_masks_98 , config1_xor_encoded_masks_99 ,
        config1_xor_encoded_masks_100 , config1_xor_encoded_masks_101 , config1_xor_encoded_masks_102 , config1_xor_encoded_masks_103 ,
        config1_xor_encoded_masks_104 , config1_xor_encoded_masks_105 , config1_xor_encoded_masks_106 , config1_xor_encoded_masks_107 ,
        config1_xor_encoded_masks_108 , config1_xor_encoded_masks_109 , config1_xor_encoded_masks_110 , config1_xor_encoded_masks_111 ,
        config1_xor_encoded_masks_112 , config1_xor_encoded_masks_113 , config1_xor_encoded_masks_114 , config1_xor_encoded_masks_115 ,
        config1_xor_encoded_masks_116 , config1_xor_encoded_masks_117 , config1_xor_encoded_masks_118 , config1_xor_encoded_masks_119 ,
        config1_xor_encoded_masks_120 , config1_xor_encoded_masks_121 , config1_xor_encoded_masks_122 , config1_xor_encoded_masks_123 ,
        config1_xor_encoded_masks_124 , config1_xor_encoded_masks_125 , config1_xor_encoded_masks_126 , config1_xor_encoded_masks_127 ,
        config1_xor_encoded_masks_128 , config1_xor_encoded_masks_129 , config1_xor_encoded_masks_130 , config1_xor_encoded_masks_131 ,
        config1_xor_encoded_masks_132 , config1_xor_encoded_masks_133 , config1_xor_encoded_masks_134 , config1_xor_encoded_masks_135 ,
        config1_xor_encoded_masks_136 , config1_xor_encoded_masks_137 , config1_xor_encoded_masks_138 , config1_xor_encoded_masks_139 ,
        config1_xor_encoded_masks_140 , config1_xor_encoded_masks_141 , config1_xor_encoded_masks_142 , config1_xor_encoded_masks_143 ,
        config1_xor_encoded_masks_144 , config1_xor_encoded_masks_145 , config1_xor_encoded_masks_146 , config1_xor_encoded_masks_147 ,
        config1_xor_encoded_masks_148 , config1_xor_encoded_masks_149 , edt_channels_out_from_constant_shift_control_0 , edt_channels_out_from_constant_shift_control_1 ,
        edt_channels_out_from_constant_shift_control_2 , edt_channels_out_from_constant_shift_control_3 , edt_channels_out_from_constant_shift_control_4 , edt_channels_out_from_constant_shift_control_5 ,
        edt_channels_out_from_constant_shift_control_6 , edt_channels_out_from_constant_shift_control_7 , edt_channels_out_from_constant_shift_control_8 , edt_channels_out_from_constant_shift_control_9 ,
        edt_channels_out_from_constant_shift_control_10 , edt_channels_out_from_constant_shift_control_11 , edt_channels_out_from_constant_shift_control_12 , edt_channels_out_from_constant_shift_control_13 ,
        edt_channels_out_from_constant_shift_control_14 , xor_encoded_masks_0 , xor_encoded_masks_1 , xor_encoded_masks_2 ,
        xor_encoded_masks_3 , xor_encoded_masks_4 , xor_encoded_masks_5 , xor_encoded_masks_6 ,
        xor_encoded_masks_7 , xor_encoded_masks_8 , xor_encoded_masks_9 , xor_encoded_masks_10 ,
        xor_encoded_masks_11 , xor_encoded_masks_12 , xor_encoded_masks_13 , xor_encoded_masks_14 ,
        xor_encoded_masks_15 , xor_encoded_masks_16 , xor_encoded_masks_17 , xor_encoded_masks_18 ,
        xor_encoded_masks_19 , xor_encoded_masks_20 , xor_encoded_masks_21 , xor_encoded_masks_22 ,
        xor_encoded_masks_23 , xor_encoded_masks_24 , xor_encoded_masks_25 , xor_encoded_masks_26 ,
        xor_encoded_masks_27 , xor_encoded_masks_28 , xor_encoded_masks_29 , xor_encoded_masks_30 ,
        xor_encoded_masks_31 , xor_encoded_masks_32 , xor_encoded_masks_33 , xor_encoded_masks_34 ,
        xor_encoded_masks_35 , xor_encoded_masks_36 , xor_encoded_masks_37 , xor_encoded_masks_38 ,
        xor_encoded_masks_39 , xor_encoded_masks_40 , xor_encoded_masks_41 , xor_encoded_masks_42 ,
        xor_encoded_masks_43 , xor_encoded_masks_44 , xor_encoded_masks_45 , xor_encoded_masks_46 ,
        xor_encoded_masks_47 , xor_encoded_masks_48 , xor_encoded_masks_49 , xor_encoded_masks_50 ,
        xor_encoded_masks_51 , xor_encoded_masks_52 , xor_encoded_masks_53 , xor_encoded_masks_54 ,
        xor_encoded_masks_55 , xor_encoded_masks_56 , xor_encoded_masks_57 , xor_encoded_masks_58 ,
        xor_encoded_masks_59 , xor_encoded_masks_60 , xor_encoded_masks_61 , xor_encoded_masks_62 ,
        xor_encoded_masks_63 , xor_encoded_masks_64 , xor_encoded_masks_65 , xor_encoded_masks_66 ,
        xor_encoded_masks_67 , xor_encoded_masks_68 , xor_encoded_masks_69 , xor_encoded_masks_70 ,
        xor_encoded_masks_71 , xor_encoded_masks_72 , xor_encoded_masks_73 , xor_encoded_masks_74 ,
        xor_encoded_masks_75 , xor_encoded_masks_76 , xor_encoded_masks_77 , xor_encoded_masks_78 ,
        xor_encoded_masks_79 , xor_encoded_masks_80 , xor_encoded_masks_81 , xor_encoded_masks_82 ,
        xor_encoded_masks_83 , xor_encoded_masks_84 , xor_encoded_masks_85 , xor_encoded_masks_86 ,
        xor_encoded_masks_87 , xor_encoded_masks_88 , xor_encoded_masks_89 , xor_encoded_masks_90 ,
        xor_encoded_masks_91 , xor_encoded_masks_92 , xor_encoded_masks_93 , xor_encoded_masks_94 ,
        xor_encoded_masks_95 , xor_encoded_masks_96 , xor_encoded_masks_97 , xor_encoded_masks_98 ,
        xor_encoded_masks_99 , xor_encoded_masks_100 , xor_encoded_masks_101 , xor_encoded_masks_102 ,
        xor_encoded_masks_103 , xor_encoded_masks_104 , xor_encoded_masks_105 , xor_encoded_masks_106 ,
        xor_encoded_masks_107 , xor_encoded_masks_108 , xor_encoded_masks_109 , xor_encoded_masks_110 ,
        xor_encoded_masks_111 , xor_encoded_masks_112 , xor_encoded_masks_113 , xor_encoded_masks_114 ,
        xor_encoded_masks_115 , xor_encoded_masks_116 , xor_encoded_masks_117 , xor_encoded_masks_118 ,
        xor_encoded_masks_119 , xor_encoded_masks_120 , xor_encoded_masks_121 , xor_encoded_masks_122 ,
        xor_encoded_masks_123 , xor_encoded_masks_124 , xor_encoded_masks_125 , xor_encoded_masks_126 ,
        xor_encoded_masks_127 , xor_encoded_masks_128 , xor_encoded_masks_129 , xor_encoded_masks_130 ,
        xor_encoded_masks_131 , xor_encoded_masks_132 , xor_encoded_masks_133 , xor_encoded_masks_134 ,
        xor_encoded_masks_135 , xor_encoded_masks_136 , xor_encoded_masks_137 , xor_encoded_masks_138 ,
        xor_encoded_masks_139 , xor_encoded_masks_140 , xor_encoded_masks_141 , xor_encoded_masks_142 ,
        xor_encoded_masks_143 , xor_encoded_masks_144 , xor_encoded_masks_145 , xor_encoded_masks_146 ,
        xor_encoded_masks_147 , xor_encoded_masks_148 , xor_encoded_masks_149 , xor_decoded_masks_0_0 ,
        xor_decoded_masks_0_1 , xor_decoded_masks_0_2 , xor_decoded_masks_0_3 , xor_decoded_masks_0_4 ,
        xor_decoded_masks_0_5 , xor_decoded_masks_0_6 , xor_decoded_masks_0_7 , xor_decoded_masks_0_8 ,
        xor_decoded_masks_0_9 , xor_decoded_masks_0_10 , xor_decoded_masks_0_11 , xor_decoded_masks_0_12 ,
        xor_decoded_masks_0_13 , xor_decoded_masks_0_14 , xor_decoded_masks_0_15 , xor_decoded_masks_0_16 ,
        xor_decoded_masks_0_17 , xor_decoded_masks_0_18 , xor_decoded_masks_0_19 , xor_decoded_masks_0_20 ,
        xor_decoded_masks_0_21 , xor_decoded_masks_0_22 , xor_decoded_masks_0_23 , xor_decoded_masks_0_24 ,
        xor_decoded_masks_0_25 , xor_decoded_masks_0_26 , xor_decoded_masks_0_27 , xor_decoded_masks_0_28 ,
        xor_decoded_masks_0_29 , xor_decoded_masks_0_30 , xor_decoded_masks_0_31 , xor_decoded_masks_0_32 ,
        xor_decoded_masks_0_33 , xor_decoded_masks_0_34 , xor_decoded_masks_0_35 , xor_decoded_masks_0_36 ,
        xor_decoded_masks_0_37 , xor_decoded_masks_0_38 , xor_decoded_masks_0_39 , xor_decoded_masks_0_40 ,
        xor_decoded_masks_0_41 , xor_decoded_masks_0_42 , xor_decoded_masks_0_43 , xor_decoded_masks_0_44 ,
        xor_decoded_masks_0_45 , xor_decoded_masks_0_46 , xor_decoded_masks_0_47 , xor_decoded_masks_0_48 ,
        xor_decoded_masks_0_49 , xor_decoded_masks_0_50 , xor_decoded_masks_0_51 , xor_decoded_masks_0_52 ,
        xor_decoded_masks_0_53 , xor_decoded_masks_1_0 , xor_decoded_masks_1_1 , xor_decoded_masks_1_2 ,
        xor_decoded_masks_1_3 , xor_decoded_masks_1_4 , xor_decoded_masks_1_5 , xor_decoded_masks_1_6 ,
        xor_decoded_masks_1_7 , xor_decoded_masks_1_8 , xor_decoded_masks_1_9 , xor_decoded_masks_1_10 ,
        xor_decoded_masks_1_11 , xor_decoded_masks_1_12 , xor_decoded_masks_1_13 , xor_decoded_masks_1_14 ,
        xor_decoded_masks_1_15 , xor_decoded_masks_1_16 , xor_decoded_masks_1_17 , xor_decoded_masks_1_18 ,
        xor_decoded_masks_1_19 , xor_decoded_masks_1_20 , xor_decoded_masks_1_21 , xor_decoded_masks_1_22 ,
        xor_decoded_masks_1_23 , xor_decoded_masks_1_24 , xor_decoded_masks_1_25 , xor_decoded_masks_1_26 ,
        xor_decoded_masks_1_27 , xor_decoded_masks_1_28 , xor_decoded_masks_1_29 , xor_decoded_masks_1_30 ,
        xor_decoded_masks_1_31 , xor_decoded_masks_1_32 , xor_decoded_masks_1_33 , xor_decoded_masks_1_34 ,
        xor_decoded_masks_1_35 , xor_decoded_masks_1_36 , xor_decoded_masks_1_37 , xor_decoded_masks_1_38 ,
        xor_decoded_masks_1_39 , xor_decoded_masks_1_40 , xor_decoded_masks_1_41 , xor_decoded_masks_1_42 ,
        xor_decoded_masks_1_43 , xor_decoded_masks_1_44 , xor_decoded_masks_1_45 , xor_decoded_masks_1_46 ,
        xor_decoded_masks_1_47 , xor_decoded_masks_1_48 , xor_decoded_masks_1_49 , xor_decoded_masks_1_50 ,
        xor_decoded_masks_1_51 , xor_decoded_masks_1_52 , xor_decoded_masks_2_0 , xor_decoded_masks_2_1 ,
        xor_decoded_masks_2_2 , xor_decoded_masks_2_3 , xor_decoded_masks_2_4 , xor_decoded_masks_2_5 ,
        xor_decoded_masks_2_6 , xor_decoded_masks_2_7 , xor_decoded_masks_2_8 , xor_decoded_masks_2_9 ,
        xor_decoded_masks_2_10 , xor_decoded_masks_2_11 , xor_decoded_masks_2_12 , xor_decoded_masks_2_13 ,
        xor_decoded_masks_2_14 , xor_decoded_masks_2_15 , xor_decoded_masks_2_16 , xor_decoded_masks_2_17 ,
        xor_decoded_masks_2_18 , xor_decoded_masks_2_19 , xor_decoded_masks_2_20 , xor_decoded_masks_2_21 ,
        xor_decoded_masks_2_22 , xor_decoded_masks_2_23 , xor_decoded_masks_2_24 , xor_decoded_masks_2_25 ,
        xor_decoded_masks_2_26 , xor_decoded_masks_2_27 , xor_decoded_masks_2_28 , xor_decoded_masks_2_29 ,
        xor_decoded_masks_2_30 , xor_decoded_masks_2_31 , xor_decoded_masks_2_32 , xor_decoded_masks_2_33 ,
        xor_decoded_masks_2_34 , xor_decoded_masks_2_35 , xor_decoded_masks_2_36 , xor_decoded_masks_2_37 ,
        xor_decoded_masks_2_38 , xor_decoded_masks_2_39 , xor_decoded_masks_2_40 , xor_decoded_masks_2_41 ,
        xor_decoded_masks_2_42 , xor_decoded_masks_2_43 , xor_decoded_masks_2_44 , xor_decoded_masks_2_45 ,
        xor_decoded_masks_2_46 , xor_decoded_masks_2_47 , xor_decoded_masks_2_48 , xor_decoded_masks_2_49 ,
        xor_decoded_masks_2_50 , xor_decoded_masks_2_51 , xor_decoded_masks_2_52 , xor_decoded_masks_3_0 ,
        xor_decoded_masks_3_1 , xor_decoded_masks_3_2 , xor_decoded_masks_3_3 , xor_decoded_masks_3_4 ,
        xor_decoded_masks_3_5 , xor_decoded_masks_3_6 , xor_decoded_masks_3_7 , xor_decoded_masks_3_8 ,
        xor_decoded_masks_3_9 , xor_decoded_masks_3_10 , xor_decoded_masks_3_11 , xor_decoded_masks_3_12 ,
        xor_decoded_masks_3_13 , xor_decoded_masks_3_14 , xor_decoded_masks_3_15 , xor_decoded_masks_3_16 ,
        xor_decoded_masks_3_17 , xor_decoded_masks_3_18 , xor_decoded_masks_3_19 , xor_decoded_masks_3_20 ,
        xor_decoded_masks_3_21 , xor_decoded_masks_3_22 , xor_decoded_masks_3_23 , xor_decoded_masks_3_24 ,
        xor_decoded_masks_3_25 , xor_decoded_masks_3_26 , xor_decoded_masks_3_27 , xor_decoded_masks_3_28 ,
        xor_decoded_masks_3_29 , xor_decoded_masks_3_30 , xor_decoded_masks_3_31 , xor_decoded_masks_3_32 ,
        xor_decoded_masks_3_33 , xor_decoded_masks_3_34 , xor_decoded_masks_3_35 , xor_decoded_masks_3_36 ,
        xor_decoded_masks_3_37 , xor_decoded_masks_3_38 , xor_decoded_masks_3_39 , xor_decoded_masks_3_40 ,
        xor_decoded_masks_3_41 , xor_decoded_masks_3_42 , xor_decoded_masks_3_43 , xor_decoded_masks_3_44 ,
        xor_decoded_masks_3_45 , xor_decoded_masks_3_46 , xor_decoded_masks_3_47 , xor_decoded_masks_3_48 ,
        xor_decoded_masks_3_49 , xor_decoded_masks_3_50 , xor_decoded_masks_3_51 , xor_decoded_masks_3_52 ,
        xor_decoded_masks_4_0 , xor_decoded_masks_4_1 , xor_decoded_masks_4_2 , xor_decoded_masks_4_3 ,
        xor_decoded_masks_4_4 , xor_decoded_masks_4_5 , xor_decoded_masks_4_6 , xor_decoded_masks_4_7 ,
        xor_decoded_masks_4_8 , xor_decoded_masks_4_9 , xor_decoded_masks_4_10 , xor_decoded_masks_4_11 ,
        xor_decoded_masks_4_12 , xor_decoded_masks_4_13 , xor_decoded_masks_4_14 , xor_decoded_masks_4_15 ,
        xor_decoded_masks_4_16 , xor_decoded_masks_4_17 , xor_decoded_masks_4_18 , xor_decoded_masks_4_19 ,
        xor_decoded_masks_4_20 , xor_decoded_masks_4_21 , xor_decoded_masks_4_22 , xor_decoded_masks_4_23 ,
        xor_decoded_masks_4_24 , xor_decoded_masks_4_25 , xor_decoded_masks_4_26 , xor_decoded_masks_4_27 ,
        xor_decoded_masks_4_28 , xor_decoded_masks_4_29 , xor_decoded_masks_4_30 , xor_decoded_masks_4_31 ,
        xor_decoded_masks_4_32 , xor_decoded_masks_4_33 , xor_decoded_masks_4_34 , xor_decoded_masks_4_35 ,
        xor_decoded_masks_4_36 , xor_decoded_masks_4_37 , xor_decoded_masks_4_38 , xor_decoded_masks_4_39 ,
        xor_decoded_masks_4_40 , xor_decoded_masks_4_41 , xor_decoded_masks_4_42 , xor_decoded_masks_4_43 ,
        xor_decoded_masks_4_44 , xor_decoded_masks_4_45 , xor_decoded_masks_4_46 , xor_decoded_masks_4_47 ,
        xor_decoded_masks_4_48 , xor_decoded_masks_4_49 , xor_decoded_masks_4_50 , xor_decoded_masks_4_51 ,
        xor_decoded_masks_4_52 , xor_decoded_masks_5_0 , xor_decoded_masks_5_1 , xor_decoded_masks_5_2 ,
        xor_decoded_masks_5_3 , xor_decoded_masks_5_4 , xor_decoded_masks_5_5 , xor_decoded_masks_5_6 ,
        xor_decoded_masks_5_7 , xor_decoded_masks_5_8 , xor_decoded_masks_5_9 , xor_decoded_masks_5_10 ,
        xor_decoded_masks_5_11 , xor_decoded_masks_5_12 , xor_decoded_masks_5_13 , xor_decoded_masks_5_14 ,
        xor_decoded_masks_5_15 , xor_decoded_masks_5_16 , xor_decoded_masks_5_17 , xor_decoded_masks_5_18 ,
        xor_decoded_masks_5_19 , xor_decoded_masks_5_20 , xor_decoded_masks_5_21 , xor_decoded_masks_5_22 ,
        xor_decoded_masks_5_23 , xor_decoded_masks_5_24 , xor_decoded_masks_5_25 , xor_decoded_masks_5_26 ,
        xor_decoded_masks_5_27 , xor_decoded_masks_5_28 , xor_decoded_masks_5_29 , xor_decoded_masks_5_30 ,
        xor_decoded_masks_5_31 , xor_decoded_masks_5_32 , xor_decoded_masks_5_33 , xor_decoded_masks_5_34 ,
        xor_decoded_masks_5_35 , xor_decoded_masks_5_36 , xor_decoded_masks_5_37 , xor_decoded_masks_5_38 ,
        xor_decoded_masks_5_39 , xor_decoded_masks_5_40 , xor_decoded_masks_5_41 , xor_decoded_masks_5_42 ,
        xor_decoded_masks_5_43 , xor_decoded_masks_5_44 , xor_decoded_masks_5_45 , xor_decoded_masks_5_46 ,
        xor_decoded_masks_5_47 , xor_decoded_masks_5_48 , xor_decoded_masks_5_49 , xor_decoded_masks_5_50 ,
        xor_decoded_masks_5_51 , xor_decoded_masks_5_52 , xor_decoded_masks_6_0 , xor_decoded_masks_6_1 ,
        xor_decoded_masks_6_2 , xor_decoded_masks_6_3 , xor_decoded_masks_6_4 , xor_decoded_masks_6_5 ,
        xor_decoded_masks_6_6 , xor_decoded_masks_6_7 , xor_decoded_masks_6_8 , xor_decoded_masks_6_9 ,
        xor_decoded_masks_6_10 , xor_decoded_masks_6_11 , xor_decoded_masks_6_12 , xor_decoded_masks_6_13 ,
        xor_decoded_masks_6_14 , xor_decoded_masks_6_15 , xor_decoded_masks_6_16 , xor_decoded_masks_6_17 ,
        xor_decoded_masks_6_18 , xor_decoded_masks_6_19 , xor_decoded_masks_6_20 , xor_decoded_masks_6_21 ,
        xor_decoded_masks_6_22 , xor_decoded_masks_6_23 , xor_decoded_masks_6_24 , xor_decoded_masks_6_25 ,
        xor_decoded_masks_6_26 , xor_decoded_masks_6_27 , xor_decoded_masks_6_28 , xor_decoded_masks_6_29 ,
        xor_decoded_masks_6_30 , xor_decoded_masks_6_31 , xor_decoded_masks_6_32 , xor_decoded_masks_6_33 ,
        xor_decoded_masks_6_34 , xor_decoded_masks_6_35 , xor_decoded_masks_6_36 , xor_decoded_masks_6_37 ,
        xor_decoded_masks_6_38 , xor_decoded_masks_6_39 , xor_decoded_masks_6_40 , xor_decoded_masks_6_41 ,
        xor_decoded_masks_6_42 , xor_decoded_masks_6_43 , xor_decoded_masks_6_44 , xor_decoded_masks_6_45 ,
        xor_decoded_masks_6_46 , xor_decoded_masks_6_47 , xor_decoded_masks_6_48 , xor_decoded_masks_6_49 ,
        xor_decoded_masks_6_50 , xor_decoded_masks_6_51 , xor_decoded_masks_6_52 , xor_decoded_masks_7_0 ,
        xor_decoded_masks_7_1 , xor_decoded_masks_7_2 , xor_decoded_masks_7_3 , xor_decoded_masks_7_4 ,
        xor_decoded_masks_7_5 , xor_decoded_masks_7_6 , xor_decoded_masks_7_7 , xor_decoded_masks_7_8 ,
        xor_decoded_masks_7_9 , xor_decoded_masks_7_10 , xor_decoded_masks_7_11 , xor_decoded_masks_7_12 ,
        xor_decoded_masks_7_13 , xor_decoded_masks_7_14 , xor_decoded_masks_7_15 , xor_decoded_masks_7_16 ,
        xor_decoded_masks_7_17 , xor_decoded_masks_7_18 , xor_decoded_masks_7_19 , xor_decoded_masks_7_20 ,
        xor_decoded_masks_7_21 , xor_decoded_masks_7_22 , xor_decoded_masks_7_23 , xor_decoded_masks_7_24 ,
        xor_decoded_masks_7_25 , xor_decoded_masks_7_26 , xor_decoded_masks_7_27 , xor_decoded_masks_7_28 ,
        xor_decoded_masks_7_29 , xor_decoded_masks_7_30 , xor_decoded_masks_7_31 , xor_decoded_masks_7_32 ,
        xor_decoded_masks_7_33 , xor_decoded_masks_7_34 , xor_decoded_masks_7_35 , xor_decoded_masks_7_36 ,
        xor_decoded_masks_7_37 , xor_decoded_masks_7_38 , xor_decoded_masks_7_39 , xor_decoded_masks_7_40 ,
        xor_decoded_masks_7_41 , xor_decoded_masks_7_42 , xor_decoded_masks_7_43 , xor_decoded_masks_7_44 ,
        xor_decoded_masks_7_45 , xor_decoded_masks_7_46 , xor_decoded_masks_7_47 , xor_decoded_masks_7_48 ,
        xor_decoded_masks_7_49 , xor_decoded_masks_7_50 , xor_decoded_masks_7_51 , xor_decoded_masks_7_52 ,
        xor_decoded_masks_8_0 , xor_decoded_masks_8_1 , xor_decoded_masks_8_2 , xor_decoded_masks_8_3 ,
        xor_decoded_masks_8_4 , xor_decoded_masks_8_5 , xor_decoded_masks_8_6 , xor_decoded_masks_8_7 ,
        xor_decoded_masks_8_8 , xor_decoded_masks_8_9 , xor_decoded_masks_8_10 , xor_decoded_masks_8_11 ,
        xor_decoded_masks_8_12 , xor_decoded_masks_8_13 , xor_decoded_masks_8_14 , xor_decoded_masks_8_15 ,
        xor_decoded_masks_8_16 , xor_decoded_masks_8_17 , xor_decoded_masks_8_18 , xor_decoded_masks_8_19 ,
        xor_decoded_masks_8_20 , xor_decoded_masks_8_21 , xor_decoded_masks_8_22 , xor_decoded_masks_8_23 ,
        xor_decoded_masks_8_24 , xor_decoded_masks_8_25 , xor_decoded_masks_8_26 , xor_decoded_masks_8_27 ,
        xor_decoded_masks_8_28 , xor_decoded_masks_8_29 , xor_decoded_masks_8_30 , xor_decoded_masks_8_31 ,
        xor_decoded_masks_8_32 , xor_decoded_masks_8_33 , xor_decoded_masks_8_34 , xor_decoded_masks_8_35 ,
        xor_decoded_masks_8_36 , xor_decoded_masks_8_37 , xor_decoded_masks_8_38 , xor_decoded_masks_8_39 ,
        xor_decoded_masks_8_40 , xor_decoded_masks_8_41 , xor_decoded_masks_8_42 , xor_decoded_masks_8_43 ,
        xor_decoded_masks_8_44 , xor_decoded_masks_8_45 , xor_decoded_masks_8_46 , xor_decoded_masks_8_47 ,
        xor_decoded_masks_8_48 , xor_decoded_masks_8_49 , xor_decoded_masks_8_50 , xor_decoded_masks_8_51 ,
        xor_decoded_masks_8_52 , xor_decoded_masks_9_0 , xor_decoded_masks_9_1 , xor_decoded_masks_9_2 ,
        xor_decoded_masks_9_3 , xor_decoded_masks_9_4 , xor_decoded_masks_9_5 , xor_decoded_masks_9_6 ,
        xor_decoded_masks_9_7 , xor_decoded_masks_9_8 , xor_decoded_masks_9_9 , xor_decoded_masks_9_10 ,
        xor_decoded_masks_9_11 , xor_decoded_masks_9_12 , xor_decoded_masks_9_13 , xor_decoded_masks_9_14 ,
        xor_decoded_masks_9_15 , xor_decoded_masks_9_16 , xor_decoded_masks_9_17 , xor_decoded_masks_9_18 ,
        xor_decoded_masks_9_19 , xor_decoded_masks_9_20 , xor_decoded_masks_9_21 , xor_decoded_masks_9_22 ,
        xor_decoded_masks_9_23 , xor_decoded_masks_9_24 , xor_decoded_masks_9_25 , xor_decoded_masks_9_26 ,
        xor_decoded_masks_9_27 , xor_decoded_masks_9_28 , xor_decoded_masks_9_29 , xor_decoded_masks_9_30 ,
        xor_decoded_masks_9_31 , xor_decoded_masks_9_32 , xor_decoded_masks_9_33 , xor_decoded_masks_9_34 ,
        xor_decoded_masks_9_35 , xor_decoded_masks_9_36 , xor_decoded_masks_9_37 , xor_decoded_masks_9_38 ,
        xor_decoded_masks_9_39 , xor_decoded_masks_9_40 , xor_decoded_masks_9_41 , xor_decoded_masks_9_42 ,
        xor_decoded_masks_9_43 , xor_decoded_masks_9_44 , xor_decoded_masks_9_45 , xor_decoded_masks_9_46 ,
        xor_decoded_masks_9_47 , xor_decoded_masks_9_48 , xor_decoded_masks_9_49 , xor_decoded_masks_9_50 ,
        xor_decoded_masks_9_51 , xor_decoded_masks_9_52 , xor_decoded_masks_10_0 , xor_decoded_masks_10_1 ,
        xor_decoded_masks_10_2 , xor_decoded_masks_10_3 , xor_decoded_masks_10_4 , xor_decoded_masks_10_5 ,
        xor_decoded_masks_10_6 , xor_decoded_masks_10_7 , xor_decoded_masks_10_8 , xor_decoded_masks_10_9 ,
        xor_decoded_masks_10_10 , xor_decoded_masks_10_11 , xor_decoded_masks_10_12 , xor_decoded_masks_10_13 ,
        xor_decoded_masks_10_14 , xor_decoded_masks_10_15 , xor_decoded_masks_10_16 , xor_decoded_masks_10_17 ,
        xor_decoded_masks_10_18 , xor_decoded_masks_10_19 , xor_decoded_masks_10_20 , xor_decoded_masks_10_21 ,
        xor_decoded_masks_10_22 , xor_decoded_masks_10_23 , xor_decoded_masks_10_24 , xor_decoded_masks_10_25 ,
        xor_decoded_masks_10_26 , xor_decoded_masks_10_27 , xor_decoded_masks_10_28 , xor_decoded_masks_10_29 ,
        xor_decoded_masks_10_30 , xor_decoded_masks_10_31 , xor_decoded_masks_10_32 , xor_decoded_masks_10_33 ,
        xor_decoded_masks_10_34 , xor_decoded_masks_10_35 , xor_decoded_masks_10_36 , xor_decoded_masks_10_37 ,
        xor_decoded_masks_10_38 , xor_decoded_masks_10_39 , xor_decoded_masks_10_40 , xor_decoded_masks_10_41 ,
        xor_decoded_masks_10_42 , xor_decoded_masks_10_43 , xor_decoded_masks_10_44 , xor_decoded_masks_10_45 ,
        xor_decoded_masks_10_46 , xor_decoded_masks_10_47 , xor_decoded_masks_10_48 , xor_decoded_masks_10_49 ,
        xor_decoded_masks_10_50 , xor_decoded_masks_10_51 , xor_decoded_masks_10_52 , xor_decoded_masks_11_0 ,
        xor_decoded_masks_11_1 , xor_decoded_masks_11_2 , xor_decoded_masks_11_3 , xor_decoded_masks_11_4 ,
        xor_decoded_masks_11_5 , xor_decoded_masks_11_6 , xor_decoded_masks_11_7 , xor_decoded_masks_11_8 ,
        xor_decoded_masks_11_9 , xor_decoded_masks_11_10 , xor_decoded_masks_11_11 , xor_decoded_masks_11_12 ,
        xor_decoded_masks_11_13 , xor_decoded_masks_11_14 , xor_decoded_masks_11_15 , xor_decoded_masks_11_16 ,
        xor_decoded_masks_11_17 , xor_decoded_masks_11_18 , xor_decoded_masks_11_19 , xor_decoded_masks_11_20 ,
        xor_decoded_masks_11_21 , xor_decoded_masks_11_22 , xor_decoded_masks_11_23 , xor_decoded_masks_11_24 ,
        xor_decoded_masks_11_25 , xor_decoded_masks_11_26 , xor_decoded_masks_11_27 , xor_decoded_masks_11_28 ,
        xor_decoded_masks_11_29 , xor_decoded_masks_11_30 , xor_decoded_masks_11_31 , xor_decoded_masks_11_32 ,
        xor_decoded_masks_11_33 , xor_decoded_masks_11_34 , xor_decoded_masks_11_35 , xor_decoded_masks_11_36 ,
        xor_decoded_masks_11_37 , xor_decoded_masks_11_38 , xor_decoded_masks_11_39 , xor_decoded_masks_11_40 ,
        xor_decoded_masks_11_41 , xor_decoded_masks_11_42 , xor_decoded_masks_11_43 , xor_decoded_masks_11_44 ,
        xor_decoded_masks_11_45 , xor_decoded_masks_11_46 , xor_decoded_masks_11_47 , xor_decoded_masks_11_48 ,
        xor_decoded_masks_11_49 , xor_decoded_masks_11_50 , xor_decoded_masks_11_51 , xor_decoded_masks_11_52 ,
        xor_decoded_masks_12_0 , xor_decoded_masks_12_1 , xor_decoded_masks_12_2 , xor_decoded_masks_12_3 ,
        xor_decoded_masks_12_4 , xor_decoded_masks_12_5 , xor_decoded_masks_12_6 , xor_decoded_masks_12_7 ,
        xor_decoded_masks_12_8 , xor_decoded_masks_12_9 , xor_decoded_masks_12_10 , xor_decoded_masks_12_11 ,
        xor_decoded_masks_12_12 , xor_decoded_masks_12_13 , xor_decoded_masks_12_14 , xor_decoded_masks_12_15 ,
        xor_decoded_masks_12_16 , xor_decoded_masks_12_17 , xor_decoded_masks_12_18 , xor_decoded_masks_12_19 ,
        xor_decoded_masks_12_20 , xor_decoded_masks_12_21 , xor_decoded_masks_12_22 , xor_decoded_masks_12_23 ,
        xor_decoded_masks_12_24 , xor_decoded_masks_12_25 , xor_decoded_masks_12_26 , xor_decoded_masks_12_27 ,
        xor_decoded_masks_12_28 , xor_decoded_masks_12_29 , xor_decoded_masks_12_30 , xor_decoded_masks_12_31 ,
        xor_decoded_masks_12_32 , xor_decoded_masks_12_33 , xor_decoded_masks_12_34 , xor_decoded_masks_12_35 ,
        xor_decoded_masks_12_36 , xor_decoded_masks_12_37 , xor_decoded_masks_12_38 , xor_decoded_masks_12_39 ,
        xor_decoded_masks_12_40 , xor_decoded_masks_12_41 , xor_decoded_masks_12_42 , xor_decoded_masks_12_43 ,
        xor_decoded_masks_12_44 , xor_decoded_masks_12_45 , xor_decoded_masks_12_46 , xor_decoded_masks_12_47 ,
        xor_decoded_masks_12_48 , xor_decoded_masks_12_49 , xor_decoded_masks_12_50 , xor_decoded_masks_12_51 ,
        xor_decoded_masks_12_52 , xor_decoded_masks_13_0 , xor_decoded_masks_13_1 , xor_decoded_masks_13_2 ,
        xor_decoded_masks_13_3 , xor_decoded_masks_13_4 , xor_decoded_masks_13_5 , xor_decoded_masks_13_6 ,
        xor_decoded_masks_13_7 , xor_decoded_masks_13_8 , xor_decoded_masks_13_9 , xor_decoded_masks_13_10 ,
        xor_decoded_masks_13_11 , xor_decoded_masks_13_12 , xor_decoded_masks_13_13 , xor_decoded_masks_13_14 ,
        xor_decoded_masks_13_15 , xor_decoded_masks_13_16 , xor_decoded_masks_13_17 , xor_decoded_masks_13_18 ,
        xor_decoded_masks_13_19 , xor_decoded_masks_13_20 , xor_decoded_masks_13_21 , xor_decoded_masks_13_22 ,
        xor_decoded_masks_13_23 , xor_decoded_masks_13_24 , xor_decoded_masks_13_25 , xor_decoded_masks_13_26 ,
        xor_decoded_masks_13_27 , xor_decoded_masks_13_28 , xor_decoded_masks_13_29 , xor_decoded_masks_13_30 ,
        xor_decoded_masks_13_31 , xor_decoded_masks_13_32 , xor_decoded_masks_13_33 , xor_decoded_masks_13_34 ,
        xor_decoded_masks_13_35 , xor_decoded_masks_13_36 , xor_decoded_masks_13_37 , xor_decoded_masks_13_38 ,
        xor_decoded_masks_13_39 , xor_decoded_masks_13_40 , xor_decoded_masks_13_41 , xor_decoded_masks_13_42 ,
        xor_decoded_masks_13_43 , xor_decoded_masks_13_44 , xor_decoded_masks_13_45 , xor_decoded_masks_13_46 ,
        xor_decoded_masks_13_47 , xor_decoded_masks_13_48 , xor_decoded_masks_13_49 , xor_decoded_masks_13_50 ,
        xor_decoded_masks_13_51 , xor_decoded_masks_13_52 , xor_decoded_masks_14_0 , xor_decoded_masks_14_1 ,
        xor_decoded_masks_14_2 , xor_decoded_masks_14_3 , xor_decoded_masks_14_4 , xor_decoded_masks_14_5 ,
        xor_decoded_masks_14_6 , xor_decoded_masks_14_7 , xor_decoded_masks_14_8 , xor_decoded_masks_14_9 ,
        xor_decoded_masks_14_10 , xor_decoded_masks_14_11 , xor_decoded_masks_14_12 , xor_decoded_masks_14_13 ,
        xor_decoded_masks_14_14 , xor_decoded_masks_14_15 , xor_decoded_masks_14_16 , xor_decoded_masks_14_17 ,
        xor_decoded_masks_14_18 , xor_decoded_masks_14_19 , xor_decoded_masks_14_20 , xor_decoded_masks_14_21 ,
        xor_decoded_masks_14_22 , xor_decoded_masks_14_23 , xor_decoded_masks_14_24 , xor_decoded_masks_14_25 ,
        xor_decoded_masks_14_26 , xor_decoded_masks_14_27 , xor_decoded_masks_14_28 , xor_decoded_masks_14_29 ,
        xor_decoded_masks_14_30 , xor_decoded_masks_14_31 , xor_decoded_masks_14_32 , xor_decoded_masks_14_33 ,
        xor_decoded_masks_14_34 , xor_decoded_masks_14_35 , xor_decoded_masks_14_36 , xor_decoded_masks_14_37 ,
        xor_decoded_masks_14_38 , xor_decoded_masks_14_39 , xor_decoded_masks_14_40 , xor_decoded_masks_14_41 ,
        xor_decoded_masks_14_42 , xor_decoded_masks_14_43 , xor_decoded_masks_14_44 , xor_decoded_masks_14_45 ,
        xor_decoded_masks_14_46 , xor_decoded_masks_14_47 , xor_decoded_masks_14_48 , xor_decoded_masks_14_49 ,
        xor_decoded_masks_14_50 , xor_decoded_masks_14_51 , xor_decoded_masks_14_52 , config0_onehot_decoded_masks_8_0 ,
        config0_onehot_decoded_masks_8_1 , config0_onehot_decoded_masks_8_2 , config0_onehot_decoded_masks_8_3 , config0_onehot_decoded_masks_8_4 ,
        config0_onehot_decoded_masks_8_5 , config0_onehot_decoded_masks_8_6 , config0_onehot_decoded_masks_8_7 , config0_onehot_decoded_masks_8_8 ,
        config0_onehot_decoded_masks_8_9 , config0_onehot_decoded_masks_8_10 , config0_onehot_decoded_masks_8_11 , config0_onehot_decoded_masks_8_12 ,
        config0_onehot_decoded_masks_8_13 , config0_onehot_decoded_masks_8_14 , config0_onehot_decoded_masks_8_15 , config0_onehot_decoded_masks_8_16 ,
        config0_onehot_decoded_masks_8_17 , config0_onehot_decoded_masks_8_18 , config0_onehot_decoded_masks_8_19 , config0_onehot_decoded_masks_8_20 ,
        config0_onehot_decoded_masks_8_21 , config0_onehot_decoded_masks_8_22 , config0_onehot_decoded_masks_8_23 , config0_onehot_decoded_masks_8_24 ,
        config0_onehot_decoded_masks_8_25 , config0_onehot_decoded_masks_8_26 , config0_onehot_decoded_masks_8_27 , config0_onehot_decoded_masks_8_28 ,
        config0_onehot_decoded_masks_8_29 , config0_onehot_decoded_masks_8_30 , config0_onehot_decoded_masks_8_31 , config0_onehot_decoded_masks_8_32 ,
        config0_onehot_decoded_masks_8_33 , config0_onehot_decoded_masks_8_34 , config0_onehot_decoded_masks_8_35 , config0_onehot_decoded_masks_8_36 ,
        config0_onehot_decoded_masks_8_37 , config0_onehot_decoded_masks_8_38 , config0_onehot_decoded_masks_8_39 , config0_onehot_decoded_masks_8_40 ,
        config0_onehot_decoded_masks_8_41 , config0_onehot_decoded_masks_8_42 , config0_onehot_decoded_masks_8_43 , config0_onehot_decoded_masks_8_44 ,
        config0_onehot_decoded_masks_8_45 , config0_onehot_decoded_masks_8_46 , config0_onehot_decoded_masks_8_47 , config0_onehot_decoded_masks_8_48 ,
        config0_onehot_decoded_masks_8_49 , config0_onehot_decoded_masks_8_50 , config0_onehot_decoded_masks_8_51 , config0_onehot_decoded_masks_8_52 ,
        config0_onehot_decoded_masks_7_0 , config0_onehot_decoded_masks_7_1 , config0_onehot_decoded_masks_7_2 , config0_onehot_decoded_masks_7_3 ,
        config0_onehot_decoded_masks_7_4 , config0_onehot_decoded_masks_7_5 , config0_onehot_decoded_masks_7_6 , config0_onehot_decoded_masks_7_7 ,
        config0_onehot_decoded_masks_7_8 , config0_onehot_decoded_masks_7_9 , config0_onehot_decoded_masks_7_10 , config0_onehot_decoded_masks_7_11 ,
        config0_onehot_decoded_masks_7_12 , config0_onehot_decoded_masks_7_13 , config0_onehot_decoded_masks_7_14 , config0_onehot_decoded_masks_7_15 ,
        config0_onehot_decoded_masks_7_16 , config0_onehot_decoded_masks_7_17 , config0_onehot_decoded_masks_7_18 , config0_onehot_decoded_masks_7_19 ,
        config0_onehot_decoded_masks_7_20 , config0_onehot_decoded_masks_7_21 , config0_onehot_decoded_masks_7_22 , config0_onehot_decoded_masks_7_23 ,
        config0_onehot_decoded_masks_7_24 , config0_onehot_decoded_masks_7_25 , config0_onehot_decoded_masks_7_26 , config0_onehot_decoded_masks_7_27 ,
        config0_onehot_decoded_masks_7_28 , config0_onehot_decoded_masks_7_29 , config0_onehot_decoded_masks_7_30 , config0_onehot_decoded_masks_7_31 ,
        config0_onehot_decoded_masks_7_32 , config0_onehot_decoded_masks_7_33 , config0_onehot_decoded_masks_7_34 , config0_onehot_decoded_masks_7_35 ,
        config0_onehot_decoded_masks_7_36 , config0_onehot_decoded_masks_7_37 , config0_onehot_decoded_masks_7_38 , config0_onehot_decoded_masks_7_39 ,
        config0_onehot_decoded_masks_7_40 , config0_onehot_decoded_masks_7_41 , config0_onehot_decoded_masks_7_42 , config0_onehot_decoded_masks_7_43 ,
        config0_onehot_decoded_masks_7_44 , config0_onehot_decoded_masks_7_45 , config0_onehot_decoded_masks_7_46 , config0_onehot_decoded_masks_7_47 ,
        config0_onehot_decoded_masks_7_48 , config0_onehot_decoded_masks_7_49 , config0_onehot_decoded_masks_7_50 , config0_onehot_decoded_masks_7_51 ,
        config0_onehot_decoded_masks_7_52 , config0_onehot_decoded_masks_2_0 , config0_onehot_decoded_masks_2_1 , config0_onehot_decoded_masks_2_2 ,
        config0_onehot_decoded_masks_2_3 , config0_onehot_decoded_masks_2_4 , config0_onehot_decoded_masks_2_5 , config0_onehot_decoded_masks_2_6 ,
        config0_onehot_decoded_masks_2_7 , config0_onehot_decoded_masks_2_8 , config0_onehot_decoded_masks_2_9 , config0_onehot_decoded_masks_2_10 ,
        config0_onehot_decoded_masks_2_11 , config0_onehot_decoded_masks_2_12 , config0_onehot_decoded_masks_2_13 , config0_onehot_decoded_masks_2_14 ,
        config0_onehot_decoded_masks_2_15 , config0_onehot_decoded_masks_2_16 , config0_onehot_decoded_masks_2_17 , config0_onehot_decoded_masks_2_18 ,
        config0_onehot_decoded_masks_2_19 , config0_onehot_decoded_masks_2_20 , config0_onehot_decoded_masks_2_21 , config0_onehot_decoded_masks_2_22 ,
        config0_onehot_decoded_masks_2_23 , config0_onehot_decoded_masks_2_24 , config0_onehot_decoded_masks_2_25 , config0_onehot_decoded_masks_2_26 ,
        config0_onehot_decoded_masks_2_27 , config0_onehot_decoded_masks_2_28 , config0_onehot_decoded_masks_2_29 , config0_onehot_decoded_masks_2_30 ,
        config0_onehot_decoded_masks_2_31 , config0_onehot_decoded_masks_2_32 , config0_onehot_decoded_masks_2_33 , config0_onehot_decoded_masks_2_34 ,
        config0_onehot_decoded_masks_2_35 , config0_onehot_decoded_masks_2_36 , config0_onehot_decoded_masks_2_37 , config0_onehot_decoded_masks_2_38 ,
        config0_onehot_decoded_masks_2_39 , config0_onehot_decoded_masks_2_40 , config0_onehot_decoded_masks_2_41 , config0_onehot_decoded_masks_2_42 ,
        config0_onehot_decoded_masks_2_43 , config0_onehot_decoded_masks_2_44 , config0_onehot_decoded_masks_2_45 , config0_onehot_decoded_masks_2_46 ,
        config0_onehot_decoded_masks_2_47 , config0_onehot_decoded_masks_2_48 , config0_onehot_decoded_masks_2_49 , config0_onehot_decoded_masks_2_50 ,
        config0_onehot_decoded_masks_2_51 , config0_onehot_decoded_masks_2_52 , config0_onehot_decoded_masks_1_0 , config0_onehot_decoded_masks_1_1 ,
        config0_onehot_decoded_masks_1_2 , config0_onehot_decoded_masks_1_3 , config0_onehot_decoded_masks_1_4 , config0_onehot_decoded_masks_1_5 ,
        config0_onehot_decoded_masks_1_6 , config0_onehot_decoded_masks_1_7 , config0_onehot_decoded_masks_1_8 , config0_onehot_decoded_masks_1_9 ,
        config0_onehot_decoded_masks_1_10 , config0_onehot_decoded_masks_1_11 , config0_onehot_decoded_masks_1_12 , config0_onehot_decoded_masks_1_13 ,
        config0_onehot_decoded_masks_1_14 , config0_onehot_decoded_masks_1_15 , config0_onehot_decoded_masks_1_16 , config0_onehot_decoded_masks_1_17 ,
        config0_onehot_decoded_masks_1_18 , config0_onehot_decoded_masks_1_19 , config0_onehot_decoded_masks_1_20 , config0_onehot_decoded_masks_1_21 ,
        config0_onehot_decoded_masks_1_22 , config0_onehot_decoded_masks_1_23 , config0_onehot_decoded_masks_1_24 , config0_onehot_decoded_masks_1_25 ,
        config0_onehot_decoded_masks_1_26 , config0_onehot_decoded_masks_1_27 , config0_onehot_decoded_masks_1_28 , config0_onehot_decoded_masks_1_29 ,
        config0_onehot_decoded_masks_1_30 , config0_onehot_decoded_masks_1_31 , config0_onehot_decoded_masks_1_32 , config0_onehot_decoded_masks_1_33 ,
        config0_onehot_decoded_masks_1_34 , config0_onehot_decoded_masks_1_35 , config0_onehot_decoded_masks_1_36 , config0_onehot_decoded_masks_1_37 ,
        config0_onehot_decoded_masks_1_38 , config0_onehot_decoded_masks_1_39 , config0_onehot_decoded_masks_1_40 , config0_onehot_decoded_masks_1_41 ,
        config0_onehot_decoded_masks_1_42 , config0_onehot_decoded_masks_1_43 , config0_onehot_decoded_masks_1_44 , config0_onehot_decoded_masks_1_45 ,
        config0_onehot_decoded_masks_1_46 , config0_onehot_decoded_masks_1_47 , config0_onehot_decoded_masks_1_48 , config0_onehot_decoded_masks_1_49 ,
        config0_onehot_decoded_masks_1_50 , config0_onehot_decoded_masks_1_51 , config0_onehot_decoded_masks_1_52 , config0_onehot_decoded_masks_0_0 ,
        config0_onehot_decoded_masks_0_1 , config0_onehot_decoded_masks_0_2 , config0_onehot_decoded_masks_0_3 , config0_onehot_decoded_masks_0_4 ,
        config0_onehot_decoded_masks_0_5 , config0_onehot_decoded_masks_0_6 , config0_onehot_decoded_masks_0_7 , config0_onehot_decoded_masks_0_8 ,
        config0_onehot_decoded_masks_0_9 , config0_onehot_decoded_masks_0_10 , config0_onehot_decoded_masks_0_11 , config0_onehot_decoded_masks_0_12 ,
        config0_onehot_decoded_masks_0_13 , config0_onehot_decoded_masks_0_14 , config0_onehot_decoded_masks_0_15 , config0_onehot_decoded_masks_0_16 ,
        config0_onehot_decoded_masks_0_17 , config0_onehot_decoded_masks_0_18 , config0_onehot_decoded_masks_0_19 , config0_onehot_decoded_masks_0_20 ,
        config0_onehot_decoded_masks_0_21 , config0_onehot_decoded_masks_0_22 , config0_onehot_decoded_masks_0_23 , config0_onehot_decoded_masks_0_24 ,
        config0_onehot_decoded_masks_0_25 , config0_onehot_decoded_masks_0_26 , config0_onehot_decoded_masks_0_27 , config0_onehot_decoded_masks_0_28 ,
        config0_onehot_decoded_masks_0_29 , config0_onehot_decoded_masks_0_30 , config0_onehot_decoded_masks_0_31 , config0_onehot_decoded_masks_0_32 ,
        config0_onehot_decoded_masks_0_33 , config0_onehot_decoded_masks_0_34 , config0_onehot_decoded_masks_0_35 , config0_onehot_decoded_masks_0_36 ,
        config0_onehot_decoded_masks_0_37 , config0_onehot_decoded_masks_0_38 , config0_onehot_decoded_masks_0_39 , config0_onehot_decoded_masks_0_40 ,
        config0_onehot_decoded_masks_0_41 , config0_onehot_decoded_masks_0_42 , config0_onehot_decoded_masks_0_43 , config0_onehot_decoded_masks_0_44 ,
        config0_onehot_decoded_masks_0_45 , config0_onehot_decoded_masks_0_46 , config0_onehot_decoded_masks_0_47 , config0_onehot_decoded_masks_0_48 ,
        config0_onehot_decoded_masks_0_49 , config0_onehot_decoded_masks_0_50 , config0_onehot_decoded_masks_0_51 , config0_onehot_decoded_masks_0_52 ,
        config0_onehot_decoded_masks_0_53 , config0_onehot_decoded_masks_6_0 , config0_onehot_decoded_masks_6_1 , config0_onehot_decoded_masks_6_2 ,
        config0_onehot_decoded_masks_6_3 , config0_onehot_decoded_masks_6_4 , config0_onehot_decoded_masks_6_5 , config0_onehot_decoded_masks_6_6 ,
        config0_onehot_decoded_masks_6_7 , config0_onehot_decoded_masks_6_8 , config0_onehot_decoded_masks_6_9 , config0_onehot_decoded_masks_6_10 ,
        config0_onehot_decoded_masks_6_11 , config0_onehot_decoded_masks_6_12 , config0_onehot_decoded_masks_6_13 , config0_onehot_decoded_masks_6_14 ,
        config0_onehot_decoded_masks_6_15 , config0_onehot_decoded_masks_6_16 , config0_onehot_decoded_masks_6_17 , config0_onehot_decoded_masks_6_18 ,
        config0_onehot_decoded_masks_6_19 , config0_onehot_decoded_masks_6_20 , config0_onehot_decoded_masks_6_21 , config0_onehot_decoded_masks_6_22 ,
        config0_onehot_decoded_masks_6_23 , config0_onehot_decoded_masks_6_24 , config0_onehot_decoded_masks_6_25 , config0_onehot_decoded_masks_6_26 ,
        config0_onehot_decoded_masks_6_27 , config0_onehot_decoded_masks_6_28 , config0_onehot_decoded_masks_6_29 , config0_onehot_decoded_masks_6_30 ,
        config0_onehot_decoded_masks_6_31 , config0_onehot_decoded_masks_6_32 , config0_onehot_decoded_masks_6_33 , config0_onehot_decoded_masks_6_34 ,
        config0_onehot_decoded_masks_6_35 , config0_onehot_decoded_masks_6_36 , config0_onehot_decoded_masks_6_37 , config0_onehot_decoded_masks_6_38 ,
        config0_onehot_decoded_masks_6_39 , config0_onehot_decoded_masks_6_40 , config0_onehot_decoded_masks_6_41 , config0_onehot_decoded_masks_6_42 ,
        config0_onehot_decoded_masks_6_43 , config0_onehot_decoded_masks_6_44 , config0_onehot_decoded_masks_6_45 , config0_onehot_decoded_masks_6_46 ,
        config0_onehot_decoded_masks_6_47 , config0_onehot_decoded_masks_6_48 , config0_onehot_decoded_masks_6_49 , config0_onehot_decoded_masks_6_50 ,
        config0_onehot_decoded_masks_6_51 , config0_onehot_decoded_masks_6_52 , config0_onehot_decoded_masks_5_0 , config0_onehot_decoded_masks_5_1 ,
        config0_onehot_decoded_masks_5_2 , config0_onehot_decoded_masks_5_3 , config0_onehot_decoded_masks_5_4 , config0_onehot_decoded_masks_5_5 ,
        config0_onehot_decoded_masks_5_6 , config0_onehot_decoded_masks_5_7 , config0_onehot_decoded_masks_5_8 , config0_onehot_decoded_masks_5_9 ,
        config0_onehot_decoded_masks_5_10 , config0_onehot_decoded_masks_5_11 , config0_onehot_decoded_masks_5_12 , config0_onehot_decoded_masks_5_13 ,
        config0_onehot_decoded_masks_5_14 , config0_onehot_decoded_masks_5_15 , config0_onehot_decoded_masks_5_16 , config0_onehot_decoded_masks_5_17 ,
        config0_onehot_decoded_masks_5_18 , config0_onehot_decoded_masks_5_19 , config0_onehot_decoded_masks_5_20 , config0_onehot_decoded_masks_5_21 ,
        config0_onehot_decoded_masks_5_22 , config0_onehot_decoded_masks_5_23 , config0_onehot_decoded_masks_5_24 , config0_onehot_decoded_masks_5_25 ,
        config0_onehot_decoded_masks_5_26 , config0_onehot_decoded_masks_5_27 , config0_onehot_decoded_masks_5_28 , config0_onehot_decoded_masks_5_29 ,
        config0_onehot_decoded_masks_5_30 , config0_onehot_decoded_masks_5_31 , config0_onehot_decoded_masks_5_32 , config0_onehot_decoded_masks_5_33 ,
        config0_onehot_decoded_masks_5_34 , config0_onehot_decoded_masks_5_35 , config0_onehot_decoded_masks_5_36 , config0_onehot_decoded_masks_5_37 ,
        config0_onehot_decoded_masks_5_38 , config0_onehot_decoded_masks_5_39 , config0_onehot_decoded_masks_5_40 , config0_onehot_decoded_masks_5_41 ,
        config0_onehot_decoded_masks_5_42 , config0_onehot_decoded_masks_5_43 , config0_onehot_decoded_masks_5_44 , config0_onehot_decoded_masks_5_45 ,
        config0_onehot_decoded_masks_5_46 , config0_onehot_decoded_masks_5_47 , config0_onehot_decoded_masks_5_48 , config0_onehot_decoded_masks_5_49 ,
        config0_onehot_decoded_masks_5_50 , config0_onehot_decoded_masks_5_51 , config0_onehot_decoded_masks_5_52 , config0_onehot_decoded_masks_4_0 ,
        config0_onehot_decoded_masks_4_1 , config0_onehot_decoded_masks_4_2 , config0_onehot_decoded_masks_4_3 , config0_onehot_decoded_masks_4_4 ,
        config0_onehot_decoded_masks_4_5 , config0_onehot_decoded_masks_4_6 , config0_onehot_decoded_masks_4_7 , config0_onehot_decoded_masks_4_8 ,
        config0_onehot_decoded_masks_4_9 , config0_onehot_decoded_masks_4_10 , config0_onehot_decoded_masks_4_11 , config0_onehot_decoded_masks_4_12 ,
        config0_onehot_decoded_masks_4_13 , config0_onehot_decoded_masks_4_14 , config0_onehot_decoded_masks_4_15 , config0_onehot_decoded_masks_4_16 ,
        config0_onehot_decoded_masks_4_17 , config0_onehot_decoded_masks_4_18 , config0_onehot_decoded_masks_4_19 , config0_onehot_decoded_masks_4_20 ,
        config0_onehot_decoded_masks_4_21 , config0_onehot_decoded_masks_4_22 , config0_onehot_decoded_masks_4_23 , config0_onehot_decoded_masks_4_24 ,
        config0_onehot_decoded_masks_4_25 , config0_onehot_decoded_masks_4_26 , config0_onehot_decoded_masks_4_27 , config0_onehot_decoded_masks_4_28 ,
        config0_onehot_decoded_masks_4_29 , config0_onehot_decoded_masks_4_30 , config0_onehot_decoded_masks_4_31 , config0_onehot_decoded_masks_4_32 ,
        config0_onehot_decoded_masks_4_33 , config0_onehot_decoded_masks_4_34 , config0_onehot_decoded_masks_4_35 , config0_onehot_decoded_masks_4_36 ,
        config0_onehot_decoded_masks_4_37 , config0_onehot_decoded_masks_4_38 , config0_onehot_decoded_masks_4_39 , config0_onehot_decoded_masks_4_40 ,
        config0_onehot_decoded_masks_4_41 , config0_onehot_decoded_masks_4_42 , config0_onehot_decoded_masks_4_43 , config0_onehot_decoded_masks_4_44 ,
        config0_onehot_decoded_masks_4_45 , config0_onehot_decoded_masks_4_46 , config0_onehot_decoded_masks_4_47 , config0_onehot_decoded_masks_4_48 ,
        config0_onehot_decoded_masks_4_49 , config0_onehot_decoded_masks_4_50 , config0_onehot_decoded_masks_4_51 , config0_onehot_decoded_masks_4_52 ,
        config0_onehot_decoded_masks_3_0 , config0_onehot_decoded_masks_3_1 , config0_onehot_decoded_masks_3_2 , config0_onehot_decoded_masks_3_3 ,
        config0_onehot_decoded_masks_3_4 , config0_onehot_decoded_masks_3_5 , config0_onehot_decoded_masks_3_6 , config0_onehot_decoded_masks_3_7 ,
        config0_onehot_decoded_masks_3_8 , config0_onehot_decoded_masks_3_9 , config0_onehot_decoded_masks_3_10 , config0_onehot_decoded_masks_3_11 ,
        config0_onehot_decoded_masks_3_12 , config0_onehot_decoded_masks_3_13 , config0_onehot_decoded_masks_3_14 , config0_onehot_decoded_masks_3_15 ,
        config0_onehot_decoded_masks_3_16 , config0_onehot_decoded_masks_3_17 , config0_onehot_decoded_masks_3_18 , config0_onehot_decoded_masks_3_19 ,
        config0_onehot_decoded_masks_3_20 , config0_onehot_decoded_masks_3_21 , config0_onehot_decoded_masks_3_22 , config0_onehot_decoded_masks_3_23 ,
        config0_onehot_decoded_masks_3_24 , config0_onehot_decoded_masks_3_25 , config0_onehot_decoded_masks_3_26 , config0_onehot_decoded_masks_3_27 ,
        config0_onehot_decoded_masks_3_28 , config0_onehot_decoded_masks_3_29 , config0_onehot_decoded_masks_3_30 , config0_onehot_decoded_masks_3_31 ,
        config0_onehot_decoded_masks_3_32 , config0_onehot_decoded_masks_3_33 , config0_onehot_decoded_masks_3_34 , config0_onehot_decoded_masks_3_35 ,
        config0_onehot_decoded_masks_3_36 , config0_onehot_decoded_masks_3_37 , config0_onehot_decoded_masks_3_38 , config0_onehot_decoded_masks_3_39 ,
        config0_onehot_decoded_masks_3_40 , config0_onehot_decoded_masks_3_41 , config0_onehot_decoded_masks_3_42 , config0_onehot_decoded_masks_3_43 ,
        config0_onehot_decoded_masks_3_44 , config0_onehot_decoded_masks_3_45 , config0_onehot_decoded_masks_3_46 , config0_onehot_decoded_masks_3_47 ,
        config0_onehot_decoded_masks_3_48 , config0_onehot_decoded_masks_3_49 , config0_onehot_decoded_masks_3_50 , config0_onehot_decoded_masks_3_51 ,
        config0_onehot_decoded_masks_3_52 , config1_onehot_decoded_masks_1_0 , config1_onehot_decoded_masks_1_1 , config1_onehot_decoded_masks_1_2 ,
        config1_onehot_decoded_masks_1_3 , config1_onehot_decoded_masks_1_4 , config1_onehot_decoded_masks_1_5 , config1_onehot_decoded_masks_1_6 ,
        config1_onehot_decoded_masks_1_7 , config1_onehot_decoded_masks_1_8 , config1_onehot_decoded_masks_1_9 , config1_onehot_decoded_masks_1_10 ,
        config1_onehot_decoded_masks_1_11 , config1_onehot_decoded_masks_1_12 , config1_onehot_decoded_masks_1_13 , config1_onehot_decoded_masks_1_14 ,
        config1_onehot_decoded_masks_1_15 , config1_onehot_decoded_masks_1_16 , config1_onehot_decoded_masks_1_17 , config1_onehot_decoded_masks_1_18 ,
        config1_onehot_decoded_masks_1_19 , config1_onehot_decoded_masks_1_20 , config1_onehot_decoded_masks_1_21 , config1_onehot_decoded_masks_1_22 ,
        config1_onehot_decoded_masks_1_23 , config1_onehot_decoded_masks_1_24 , config1_onehot_decoded_masks_1_25 , config1_onehot_decoded_masks_1_26 ,
        config1_onehot_decoded_masks_1_27 , config1_onehot_decoded_masks_1_28 , config1_onehot_decoded_masks_1_29 , config1_onehot_decoded_masks_1_30 ,
        config1_onehot_decoded_masks_1_31 , config1_onehot_decoded_masks_1_32 , config1_onehot_decoded_masks_1_33 , config1_onehot_decoded_masks_1_34 ,
        config1_onehot_decoded_masks_1_35 , config1_onehot_decoded_masks_1_36 , config1_onehot_decoded_masks_1_37 , config1_onehot_decoded_masks_1_38 ,
        config1_onehot_decoded_masks_1_39 , config1_onehot_decoded_masks_1_40 , config1_onehot_decoded_masks_1_41 , config1_onehot_decoded_masks_1_42 ,
        config1_onehot_decoded_masks_1_43 , config1_onehot_decoded_masks_1_44 , config1_onehot_decoded_masks_1_45 , config1_onehot_decoded_masks_1_46 ,
        config1_onehot_decoded_masks_1_47 , config1_onehot_decoded_masks_1_48 , config1_onehot_decoded_masks_1_49 , config1_onehot_decoded_masks_1_50 ,
        config1_onehot_decoded_masks_1_51 , config1_onehot_decoded_masks_1_52 , config1_onehot_decoded_masks_1_53 , config1_onehot_decoded_masks_1_54 ,
        config1_onehot_decoded_masks_1_55 , config1_onehot_decoded_masks_1_56 , config1_onehot_decoded_masks_1_57 , config1_onehot_decoded_masks_1_58 ,
        config1_onehot_decoded_masks_1_59 , config1_onehot_decoded_masks_1_60 , config1_onehot_decoded_masks_1_61 , config1_onehot_decoded_masks_1_62 ,
        config1_onehot_decoded_masks_1_63 , config1_onehot_decoded_masks_1_64 , config1_onehot_decoded_masks_1_65 , config1_onehot_decoded_masks_1_66 ,
        config1_onehot_decoded_masks_1_67 , config1_onehot_decoded_masks_1_68 , config1_onehot_decoded_masks_1_69 , config1_onehot_decoded_masks_1_70 ,
        config1_onehot_decoded_masks_1_71 , config1_onehot_decoded_masks_1_72 , config1_onehot_decoded_masks_1_73 , config1_onehot_decoded_masks_1_74 ,
        config1_onehot_decoded_masks_1_75 , config1_onehot_decoded_masks_1_76 , config1_onehot_decoded_masks_1_77 , config1_onehot_decoded_masks_1_78 ,
        config1_onehot_decoded_masks_1_79 , config1_onehot_decoded_masks_1_80 , config1_onehot_decoded_masks_1_81 , config1_onehot_decoded_masks_1_82 ,
        config1_onehot_decoded_masks_1_83 , config1_onehot_decoded_masks_1_84 , config1_onehot_decoded_masks_1_85 , config1_onehot_decoded_masks_1_86 ,
        config1_onehot_decoded_masks_1_87 , config1_onehot_decoded_masks_1_88 , config1_onehot_decoded_masks_1_89 , config1_onehot_decoded_masks_1_90 ,
        config1_onehot_decoded_masks_1_91 , config1_onehot_decoded_masks_1_92 , config1_onehot_decoded_masks_1_93 , config1_onehot_decoded_masks_1_94 ,
        config1_onehot_decoded_masks_1_95 , config1_onehot_decoded_masks_1_96 , config1_onehot_decoded_masks_1_97 , config1_onehot_decoded_masks_1_98 ,
        config1_onehot_decoded_masks_1_99 , config1_onehot_decoded_masks_1_100 , config1_onehot_decoded_masks_1_101 , config1_onehot_decoded_masks_1_102 ,
        config1_onehot_decoded_masks_1_103 , config1_onehot_decoded_masks_1_104 , config1_onehot_decoded_masks_1_105 , config1_onehot_decoded_masks_2_0 ,
        config1_onehot_decoded_masks_2_1 , config1_onehot_decoded_masks_2_2 , config1_onehot_decoded_masks_2_3 , config1_onehot_decoded_masks_2_4 ,
        config1_onehot_decoded_masks_2_5 , config1_onehot_decoded_masks_2_6 , config1_onehot_decoded_masks_2_7 , config1_onehot_decoded_masks_2_8 ,
        config1_onehot_decoded_masks_2_9 , config1_onehot_decoded_masks_2_10 , config1_onehot_decoded_masks_2_11 , config1_onehot_decoded_masks_2_12 ,
        config1_onehot_decoded_masks_2_13 , config1_onehot_decoded_masks_2_14 , config1_onehot_decoded_masks_2_15 , config1_onehot_decoded_masks_2_16 ,
        config1_onehot_decoded_masks_2_17 , config1_onehot_decoded_masks_2_18 , config1_onehot_decoded_masks_2_19 , config1_onehot_decoded_masks_2_20 ,
        config1_onehot_decoded_masks_2_21 , config1_onehot_decoded_masks_2_22 , config1_onehot_decoded_masks_2_23 , config1_onehot_decoded_masks_2_24 ,
        config1_onehot_decoded_masks_2_25 , config1_onehot_decoded_masks_2_26 , config1_onehot_decoded_masks_2_27 , config1_onehot_decoded_masks_2_28 ,
        config1_onehot_decoded_masks_2_29 , config1_onehot_decoded_masks_2_30 , config1_onehot_decoded_masks_2_31 , config1_onehot_decoded_masks_2_32 ,
        config1_onehot_decoded_masks_2_33 , config1_onehot_decoded_masks_2_34 , config1_onehot_decoded_masks_2_35 , config1_onehot_decoded_masks_2_36 ,
        config1_onehot_decoded_masks_2_37 , config1_onehot_decoded_masks_2_38 , config1_onehot_decoded_masks_2_39 , config1_onehot_decoded_masks_2_40 ,
        config1_onehot_decoded_masks_2_41 , config1_onehot_decoded_masks_2_42 , config1_onehot_decoded_masks_2_43 , config1_onehot_decoded_masks_2_44 ,
        config1_onehot_decoded_masks_2_45 , config1_onehot_decoded_masks_2_46 , config1_onehot_decoded_masks_2_47 , config1_onehot_decoded_masks_2_48 ,
        config1_onehot_decoded_masks_2_49 , config1_onehot_decoded_masks_2_50 , config1_onehot_decoded_masks_2_51 , config1_onehot_decoded_masks_2_52 ,
        config1_onehot_decoded_masks_2_53 , config1_onehot_decoded_masks_2_54 , config1_onehot_decoded_masks_2_55 , config1_onehot_decoded_masks_2_56 ,
        config1_onehot_decoded_masks_2_57 , config1_onehot_decoded_masks_2_58 , config1_onehot_decoded_masks_2_59 , config1_onehot_decoded_masks_2_60 ,
        config1_onehot_decoded_masks_2_61 , config1_onehot_decoded_masks_2_62 , config1_onehot_decoded_masks_2_63 , config1_onehot_decoded_masks_2_64 ,
        config1_onehot_decoded_masks_2_65 , config1_onehot_decoded_masks_2_66 , config1_onehot_decoded_masks_2_67 , config1_onehot_decoded_masks_2_68 ,
        config1_onehot_decoded_masks_2_69 , config1_onehot_decoded_masks_2_70 , config1_onehot_decoded_masks_2_71 , config1_onehot_decoded_masks_2_72 ,
        config1_onehot_decoded_masks_2_73 , config1_onehot_decoded_masks_2_74 , config1_onehot_decoded_masks_2_75 , config1_onehot_decoded_masks_2_76 ,
        config1_onehot_decoded_masks_2_77 , config1_onehot_decoded_masks_2_78 , config1_onehot_decoded_masks_2_79 , config1_onehot_decoded_masks_2_80 ,
        config1_onehot_decoded_masks_2_81 , config1_onehot_decoded_masks_2_82 , config1_onehot_decoded_masks_2_83 , config1_onehot_decoded_masks_2_84 ,
        config1_onehot_decoded_masks_2_85 , config1_onehot_decoded_masks_2_86 , config1_onehot_decoded_masks_2_87 , config1_onehot_decoded_masks_2_88 ,
        config1_onehot_decoded_masks_2_89 , config1_onehot_decoded_masks_2_90 , config1_onehot_decoded_masks_2_91 , config1_onehot_decoded_masks_2_92 ,
        config1_onehot_decoded_masks_2_93 , config1_onehot_decoded_masks_2_94 , config1_onehot_decoded_masks_2_95 , config1_onehot_decoded_masks_2_96 ,
        config1_onehot_decoded_masks_2_97 , config1_onehot_decoded_masks_2_98 , config1_onehot_decoded_masks_2_99 , config1_onehot_decoded_masks_2_100 ,
        config1_onehot_decoded_masks_2_101 , config1_onehot_decoded_masks_2_102 , config1_onehot_decoded_masks_2_103 , config1_onehot_decoded_masks_2_104 ,
        config1_onehot_decoded_masks_2_105 , config1_onehot_decoded_masks_0_0 , config1_onehot_decoded_masks_0_1 , config1_onehot_decoded_masks_0_2 ,
        config1_onehot_decoded_masks_0_3 , config1_onehot_decoded_masks_0_4 , config1_onehot_decoded_masks_0_5 , config1_onehot_decoded_masks_0_6 ,
        config1_onehot_decoded_masks_0_7 , config1_onehot_decoded_masks_0_8 , config1_onehot_decoded_masks_0_9 , config1_onehot_decoded_masks_0_10 ,
        config1_onehot_decoded_masks_0_11 , config1_onehot_decoded_masks_0_12 , config1_onehot_decoded_masks_0_13 , config1_onehot_decoded_masks_0_14 ,
        config1_onehot_decoded_masks_0_15 , config1_onehot_decoded_masks_0_16 , config1_onehot_decoded_masks_0_17 , config1_onehot_decoded_masks_0_18 ,
        config1_onehot_decoded_masks_0_19 , config1_onehot_decoded_masks_0_20 , config1_onehot_decoded_masks_0_21 , config1_onehot_decoded_masks_0_22 ,
        config1_onehot_decoded_masks_0_23 , config1_onehot_decoded_masks_0_24 , config1_onehot_decoded_masks_0_25 , config1_onehot_decoded_masks_0_26 ,
        config1_onehot_decoded_masks_0_27 , config1_onehot_decoded_masks_0_28 , config1_onehot_decoded_masks_0_29 , config1_onehot_decoded_masks_0_30 ,
        config1_onehot_decoded_masks_0_31 , config1_onehot_decoded_masks_0_32 , config1_onehot_decoded_masks_0_33 , config1_onehot_decoded_masks_0_34 ,
        config1_onehot_decoded_masks_0_35 , config1_onehot_decoded_masks_0_36 , config1_onehot_decoded_masks_0_37 , config1_onehot_decoded_masks_0_38 ,
        config1_onehot_decoded_masks_0_39 , config1_onehot_decoded_masks_0_40 , config1_onehot_decoded_masks_0_41 , config1_onehot_decoded_masks_0_42 ,
        config1_onehot_decoded_masks_0_43 , config1_onehot_decoded_masks_0_44 , config1_onehot_decoded_masks_0_45 , config1_onehot_decoded_masks_0_46 ,
        config1_onehot_decoded_masks_0_47 , config1_onehot_decoded_masks_0_48 , config1_onehot_decoded_masks_0_49 , config1_onehot_decoded_masks_0_50 ,
        config1_onehot_decoded_masks_0_51 , config1_onehot_decoded_masks_0_52 , config1_onehot_decoded_masks_0_53 , config1_onehot_decoded_masks_0_54 ,
        config1_onehot_decoded_masks_0_55 , config1_onehot_decoded_masks_0_56 , config1_onehot_decoded_masks_0_57 , config1_onehot_decoded_masks_0_58 ,
        config1_onehot_decoded_masks_0_59 , config1_onehot_decoded_masks_0_60 , config1_onehot_decoded_masks_0_61 , config1_onehot_decoded_masks_0_62 ,
        config1_onehot_decoded_masks_0_63 , config1_onehot_decoded_masks_0_64 , config1_onehot_decoded_masks_0_65 , config1_onehot_decoded_masks_0_66 ,
        config1_onehot_decoded_masks_0_67 , config1_onehot_decoded_masks_0_68 , config1_onehot_decoded_masks_0_69 , config1_onehot_decoded_masks_0_70 ,
        config1_onehot_decoded_masks_0_71 , config1_onehot_decoded_masks_0_72 , config1_onehot_decoded_masks_0_73 , config1_onehot_decoded_masks_0_74 ,
        config1_onehot_decoded_masks_0_75 , config1_onehot_decoded_masks_0_76 , config1_onehot_decoded_masks_0_77 , config1_onehot_decoded_masks_0_78 ,
        config1_onehot_decoded_masks_0_79 , config1_onehot_decoded_masks_0_80 , config1_onehot_decoded_masks_0_81 , config1_onehot_decoded_masks_0_82 ,
        config1_onehot_decoded_masks_0_83 , config1_onehot_decoded_masks_0_84 , config1_onehot_decoded_masks_0_85 , config1_onehot_decoded_masks_0_86 ,
        config1_onehot_decoded_masks_0_87 , config1_onehot_decoded_masks_0_88 , config1_onehot_decoded_masks_0_89 , config1_onehot_decoded_masks_0_90 ,
        config1_onehot_decoded_masks_0_91 , config1_onehot_decoded_masks_0_92 , config1_onehot_decoded_masks_0_93 , config1_onehot_decoded_masks_0_94 ,
        config1_onehot_decoded_masks_0_95 , config1_onehot_decoded_masks_0_96 , config1_onehot_decoded_masks_0_97 , config1_onehot_decoded_masks_0_98 ,
        config1_onehot_decoded_masks_0_99 , config1_onehot_decoded_masks_0_100 , config1_onehot_decoded_masks_0_101 , config1_onehot_decoded_masks_0_102 ,
        config1_onehot_decoded_masks_0_103 , config1_onehot_decoded_masks_0_104 , config1_onehot_decoded_masks_0_105 , config1_onehot_decoded_masks_0_106 ,
        config1_onehot_decoded_masks_0_107 , config1_onehot_decoded_masks_0_108 , config1_onehot_decoded_masks_0_109 , config1_onehot_decoded_masks_0_110 ,
        config1_onehot_decoded_masks_0_111 , config1_onehot_decoded_masks_0_112 , config1_onehot_decoded_masks_0_113 , config1_onehot_decoded_masks_0_114 ,
        config1_onehot_decoded_masks_0_115 , config1_onehot_decoded_masks_0_116 , config1_onehot_decoded_masks_0_117 , config1_onehot_decoded_masks_0_118 ,
        config1_onehot_decoded_masks_0_119 , config1_onehot_decoded_masks_0_120 , config1_onehot_decoded_masks_0_121 , config1_onehot_decoded_masks_0_122 ,
        config1_onehot_decoded_masks_0_123 , config1_onehot_decoded_masks_0_124 , config1_onehot_decoded_masks_0_125 , config1_onehot_decoded_masks_0_126 ,
        config1_onehot_decoded_masks_0_127 , config1_onehot_decoded_masks_0_128 , config1_onehot_decoded_masks_0_129 , config1_onehot_decoded_masks_0_130 ,
        config1_onehot_decoded_masks_0_131 , config1_onehot_decoded_masks_0_132 , config1_onehot_decoded_masks_0_133 , config1_onehot_decoded_masks_0_134 ,
        config1_onehot_decoded_masks_0_135 , config1_onehot_decoded_masks_0_136 , config1_onehot_decoded_masks_0_137 , config1_onehot_decoded_masks_0_138 ,
        config1_onehot_decoded_masks_0_139 , config1_onehot_decoded_masks_0_140 , config1_onehot_decoded_masks_0_141 , config1_onehot_decoded_masks_0_142 ,
        config1_onehot_decoded_masks_0_143 , config1_onehot_decoded_masks_0_144 , config1_onehot_decoded_masks_0_145 , config1_onehot_decoded_masks_0_146 ,
        config1_onehot_decoded_masks_0_147 , config1_onehot_decoded_masks_0_148 , config1_onehot_decoded_masks_0_149 , config1_onehot_decoded_masks_0_150 ,
        config1_onehot_decoded_masks_0_151 , config1_onehot_decoded_masks_0_152 , config1_onehot_decoded_masks_0_153 , config1_onehot_decoded_masks_0_154 ,
        config1_onehot_decoded_masks_0_155 , config1_onehot_decoded_masks_0_156 , config1_onehot_decoded_masks_0_157 , config1_onehot_decoded_masks_0_158 ,
        config1_onehot_decoded_masks_0_159 , config1_onehot_decoded_masks_5_0 , config1_onehot_decoded_masks_5_1 , config1_onehot_decoded_masks_5_2 ,
        config1_onehot_decoded_masks_5_3 , config1_onehot_decoded_masks_5_4 , config1_onehot_decoded_masks_5_5 , config1_onehot_decoded_masks_5_6 ,
        config1_onehot_decoded_masks_5_7 , config1_onehot_decoded_masks_5_8 , config1_onehot_decoded_masks_5_9 , config1_onehot_decoded_masks_5_10 ,
        config1_onehot_decoded_masks_5_11 , config1_onehot_decoded_masks_5_12 , config1_onehot_decoded_masks_5_13 , config1_onehot_decoded_masks_5_14 ,
        config1_onehot_decoded_masks_5_15 , config1_onehot_decoded_masks_5_16 , config1_onehot_decoded_masks_5_17 , config1_onehot_decoded_masks_5_18 ,
        config1_onehot_decoded_masks_5_19 , config1_onehot_decoded_masks_5_20 , config1_onehot_decoded_masks_5_21 , config1_onehot_decoded_masks_5_22 ,
        config1_onehot_decoded_masks_5_23 , config1_onehot_decoded_masks_5_24 , config1_onehot_decoded_masks_5_25 , config1_onehot_decoded_masks_5_26 ,
        config1_onehot_decoded_masks_5_27 , config1_onehot_decoded_masks_5_28 , config1_onehot_decoded_masks_5_29 , config1_onehot_decoded_masks_5_30 ,
        config1_onehot_decoded_masks_5_31 , config1_onehot_decoded_masks_5_32 , config1_onehot_decoded_masks_5_33 , config1_onehot_decoded_masks_5_34 ,
        config1_onehot_decoded_masks_5_35 , config1_onehot_decoded_masks_5_36 , config1_onehot_decoded_masks_5_37 , config1_onehot_decoded_masks_5_38 ,
        config1_onehot_decoded_masks_5_39 , config1_onehot_decoded_masks_5_40 , config1_onehot_decoded_masks_5_41 , config1_onehot_decoded_masks_5_42 ,
        config1_onehot_decoded_masks_5_43 , config1_onehot_decoded_masks_5_44 , config1_onehot_decoded_masks_5_45 , config1_onehot_decoded_masks_5_46 ,
        config1_onehot_decoded_masks_5_47 , config1_onehot_decoded_masks_5_48 , config1_onehot_decoded_masks_5_49 , config1_onehot_decoded_masks_5_50 ,
        config1_onehot_decoded_masks_5_51 , config1_onehot_decoded_masks_5_52 , config1_onehot_decoded_masks_5_53 , config1_onehot_decoded_masks_5_54 ,
        config1_onehot_decoded_masks_5_55 , config1_onehot_decoded_masks_5_56 , config1_onehot_decoded_masks_5_57 , config1_onehot_decoded_masks_5_58 ,
        config1_onehot_decoded_masks_5_59 , config1_onehot_decoded_masks_5_60 , config1_onehot_decoded_masks_5_61 , config1_onehot_decoded_masks_5_62 ,
        config1_onehot_decoded_masks_5_63 , config1_onehot_decoded_masks_5_64 , config1_onehot_decoded_masks_5_65 , config1_onehot_decoded_masks_5_66 ,
        config1_onehot_decoded_masks_5_67 , config1_onehot_decoded_masks_5_68 , config1_onehot_decoded_masks_5_69 , config1_onehot_decoded_masks_5_70 ,
        config1_onehot_decoded_masks_5_71 , config1_onehot_decoded_masks_5_72 , config1_onehot_decoded_masks_5_73 , config1_onehot_decoded_masks_5_74 ,
        config1_onehot_decoded_masks_5_75 , config1_onehot_decoded_masks_5_76 , config1_onehot_decoded_masks_5_77 , config1_onehot_decoded_masks_5_78 ,
        config1_onehot_decoded_masks_5_79 , config1_onehot_decoded_masks_5_80 , config1_onehot_decoded_masks_5_81 , config1_onehot_decoded_masks_5_82 ,
        config1_onehot_decoded_masks_5_83 , config1_onehot_decoded_masks_5_84 , config1_onehot_decoded_masks_5_85 , config1_onehot_decoded_masks_5_86 ,
        config1_onehot_decoded_masks_5_87 , config1_onehot_decoded_masks_5_88 , config1_onehot_decoded_masks_5_89 , config1_onehot_decoded_masks_5_90 ,
        config1_onehot_decoded_masks_5_91 , config1_onehot_decoded_masks_5_92 , config1_onehot_decoded_masks_5_93 , config1_onehot_decoded_masks_5_94 ,
        config1_onehot_decoded_masks_5_95 , config1_onehot_decoded_masks_5_96 , config1_onehot_decoded_masks_5_97 , config1_onehot_decoded_masks_5_98 ,
        config1_onehot_decoded_masks_5_99 , config1_onehot_decoded_masks_5_100 , config1_onehot_decoded_masks_5_101 , config1_onehot_decoded_masks_5_102 ,
        config1_onehot_decoded_masks_5_103 , config1_onehot_decoded_masks_5_104 , config1_onehot_decoded_masks_5_105 , config1_onehot_decoded_masks_6_0 ,
        config1_onehot_decoded_masks_6_1 , config1_onehot_decoded_masks_6_2 , config1_onehot_decoded_masks_6_3 , config1_onehot_decoded_masks_6_4 ,
        config1_onehot_decoded_masks_6_5 , config1_onehot_decoded_masks_6_6 , config1_onehot_decoded_masks_6_7 , config1_onehot_decoded_masks_6_8 ,
        config1_onehot_decoded_masks_6_9 , config1_onehot_decoded_masks_6_10 , config1_onehot_decoded_masks_6_11 , config1_onehot_decoded_masks_6_12 ,
        config1_onehot_decoded_masks_6_13 , config1_onehot_decoded_masks_6_14 , config1_onehot_decoded_masks_6_15 , config1_onehot_decoded_masks_6_16 ,
        config1_onehot_decoded_masks_6_17 , config1_onehot_decoded_masks_6_18 , config1_onehot_decoded_masks_6_19 , config1_onehot_decoded_masks_6_20 ,
        config1_onehot_decoded_masks_6_21 , config1_onehot_decoded_masks_6_22 , config1_onehot_decoded_masks_6_23 , config1_onehot_decoded_masks_6_24 ,
        config1_onehot_decoded_masks_6_25 , config1_onehot_decoded_masks_6_26 , config1_onehot_decoded_masks_6_27 , config1_onehot_decoded_masks_6_28 ,
        config1_onehot_decoded_masks_6_29 , config1_onehot_decoded_masks_6_30 , config1_onehot_decoded_masks_6_31 , config1_onehot_decoded_masks_6_32 ,
        config1_onehot_decoded_masks_6_33 , config1_onehot_decoded_masks_6_34 , config1_onehot_decoded_masks_6_35 , config1_onehot_decoded_masks_6_36 ,
        config1_onehot_decoded_masks_6_37 , config1_onehot_decoded_masks_6_38 , config1_onehot_decoded_masks_6_39 , config1_onehot_decoded_masks_6_40 ,
        config1_onehot_decoded_masks_6_41 , config1_onehot_decoded_masks_6_42 , config1_onehot_decoded_masks_6_43 , config1_onehot_decoded_masks_6_44 ,
        config1_onehot_decoded_masks_6_45 , config1_onehot_decoded_masks_6_46 , config1_onehot_decoded_masks_6_47 , config1_onehot_decoded_masks_6_48 ,
        config1_onehot_decoded_masks_6_49 , config1_onehot_decoded_masks_6_50 , config1_onehot_decoded_masks_6_51 , config1_onehot_decoded_masks_6_52 ,
        config1_onehot_decoded_masks_6_53 , config1_onehot_decoded_masks_6_54 , config1_onehot_decoded_masks_6_55 , config1_onehot_decoded_masks_6_56 ,
        config1_onehot_decoded_masks_6_57 , config1_onehot_decoded_masks_6_58 , config1_onehot_decoded_masks_6_59 , config1_onehot_decoded_masks_6_60 ,
        config1_onehot_decoded_masks_6_61 , config1_onehot_decoded_masks_6_62 , config1_onehot_decoded_masks_6_63 , config1_onehot_decoded_masks_6_64 ,
        config1_onehot_decoded_masks_6_65 , config1_onehot_decoded_masks_6_66 , config1_onehot_decoded_masks_6_67 , config1_onehot_decoded_masks_6_68 ,
        config1_onehot_decoded_masks_6_69 , config1_onehot_decoded_masks_6_70 , config1_onehot_decoded_masks_6_71 , config1_onehot_decoded_masks_6_72 ,
        config1_onehot_decoded_masks_6_73 , config1_onehot_decoded_masks_6_74 , config1_onehot_decoded_masks_6_75 , config1_onehot_decoded_masks_6_76 ,
        config1_onehot_decoded_masks_6_77 , config1_onehot_decoded_masks_6_78 , config1_onehot_decoded_masks_6_79 , config1_onehot_decoded_masks_6_80 ,
        config1_onehot_decoded_masks_6_81 , config1_onehot_decoded_masks_6_82 , config1_onehot_decoded_masks_6_83 , config1_onehot_decoded_masks_6_84 ,
        config1_onehot_decoded_masks_6_85 , config1_onehot_decoded_masks_6_86 , config1_onehot_decoded_masks_6_87 , config1_onehot_decoded_masks_6_88 ,
        config1_onehot_decoded_masks_6_89 , config1_onehot_decoded_masks_6_90 , config1_onehot_decoded_masks_6_91 , config1_onehot_decoded_masks_6_92 ,
        config1_onehot_decoded_masks_6_93 , config1_onehot_decoded_masks_6_94 , config1_onehot_decoded_masks_6_95 , config1_onehot_decoded_masks_6_96 ,
        config1_onehot_decoded_masks_6_97 , config1_onehot_decoded_masks_6_98 , config1_onehot_decoded_masks_6_99 , config1_onehot_decoded_masks_6_100 ,
        config1_onehot_decoded_masks_6_101 , config1_onehot_decoded_masks_6_102 , config1_onehot_decoded_masks_6_103 , config1_onehot_decoded_masks_6_104 ,
        config1_onehot_decoded_masks_6_105 , config1_onehot_decoded_masks_3_0 , config1_onehot_decoded_masks_3_1 , config1_onehot_decoded_masks_3_2 ,
        config1_onehot_decoded_masks_3_3 , config1_onehot_decoded_masks_3_4 , config1_onehot_decoded_masks_3_5 , config1_onehot_decoded_masks_3_6 ,
        config1_onehot_decoded_masks_3_7 , config1_onehot_decoded_masks_3_8 , config1_onehot_decoded_masks_3_9 , config1_onehot_decoded_masks_3_10 ,
        config1_onehot_decoded_masks_3_11 , config1_onehot_decoded_masks_3_12 , config1_onehot_decoded_masks_3_13 , config1_onehot_decoded_masks_3_14 ,
        config1_onehot_decoded_masks_3_15 , config1_onehot_decoded_masks_3_16 , config1_onehot_decoded_masks_3_17 , config1_onehot_decoded_masks_3_18 ,
        config1_onehot_decoded_masks_3_19 , config1_onehot_decoded_masks_3_20 , config1_onehot_decoded_masks_3_21 , config1_onehot_decoded_masks_3_22 ,
        config1_onehot_decoded_masks_3_23 , config1_onehot_decoded_masks_3_24 , config1_onehot_decoded_masks_3_25 , config1_onehot_decoded_masks_3_26 ,
        config1_onehot_decoded_masks_3_27 , config1_onehot_decoded_masks_3_28 , config1_onehot_decoded_masks_3_29 , config1_onehot_decoded_masks_3_30 ,
        config1_onehot_decoded_masks_3_31 , config1_onehot_decoded_masks_3_32 , config1_onehot_decoded_masks_3_33 , config1_onehot_decoded_masks_3_34 ,
        config1_onehot_decoded_masks_3_35 , config1_onehot_decoded_masks_3_36 , config1_onehot_decoded_masks_3_37 , config1_onehot_decoded_masks_3_38 ,
        config1_onehot_decoded_masks_3_39 , config1_onehot_decoded_masks_3_40 , config1_onehot_decoded_masks_3_41 , config1_onehot_decoded_masks_3_42 ,
        config1_onehot_decoded_masks_3_43 , config1_onehot_decoded_masks_3_44 , config1_onehot_decoded_masks_3_45 , config1_onehot_decoded_masks_3_46 ,
        config1_onehot_decoded_masks_3_47 , config1_onehot_decoded_masks_3_48 , config1_onehot_decoded_masks_3_49 , config1_onehot_decoded_masks_3_50 ,
        config1_onehot_decoded_masks_3_51 , config1_onehot_decoded_masks_3_52 , config1_onehot_decoded_masks_3_53 , config1_onehot_decoded_masks_3_54 ,
        config1_onehot_decoded_masks_3_55 , config1_onehot_decoded_masks_3_56 , config1_onehot_decoded_masks_3_57 , config1_onehot_decoded_masks_3_58 ,
        config1_onehot_decoded_masks_3_59 , config1_onehot_decoded_masks_3_60 , config1_onehot_decoded_masks_3_61 , config1_onehot_decoded_masks_3_62 ,
        config1_onehot_decoded_masks_3_63 , config1_onehot_decoded_masks_3_64 , config1_onehot_decoded_masks_3_65 , config1_onehot_decoded_masks_3_66 ,
        config1_onehot_decoded_masks_3_67 , config1_onehot_decoded_masks_3_68 , config1_onehot_decoded_masks_3_69 , config1_onehot_decoded_masks_3_70 ,
        config1_onehot_decoded_masks_3_71 , config1_onehot_decoded_masks_3_72 , config1_onehot_decoded_masks_3_73 , config1_onehot_decoded_masks_3_74 ,
        config1_onehot_decoded_masks_3_75 , config1_onehot_decoded_masks_3_76 , config1_onehot_decoded_masks_3_77 , config1_onehot_decoded_masks_3_78 ,
        config1_onehot_decoded_masks_3_79 , config1_onehot_decoded_masks_3_80 , config1_onehot_decoded_masks_3_81 , config1_onehot_decoded_masks_3_82 ,
        config1_onehot_decoded_masks_3_83 , config1_onehot_decoded_masks_3_84 , config1_onehot_decoded_masks_3_85 , config1_onehot_decoded_masks_3_86 ,
        config1_onehot_decoded_masks_3_87 , config1_onehot_decoded_masks_3_88 , config1_onehot_decoded_masks_3_89 , config1_onehot_decoded_masks_3_90 ,
        config1_onehot_decoded_masks_3_91 , config1_onehot_decoded_masks_3_92 , config1_onehot_decoded_masks_3_93 , config1_onehot_decoded_masks_3_94 ,
        config1_onehot_decoded_masks_3_95 , config1_onehot_decoded_masks_3_96 , config1_onehot_decoded_masks_3_97 , config1_onehot_decoded_masks_3_98 ,
        config1_onehot_decoded_masks_3_99 , config1_onehot_decoded_masks_3_100 , config1_onehot_decoded_masks_3_101 , config1_onehot_decoded_masks_3_102 ,
        config1_onehot_decoded_masks_3_103 , config1_onehot_decoded_masks_3_104 , config1_onehot_decoded_masks_3_105 , config1_onehot_decoded_masks_4_0 ,
        config1_onehot_decoded_masks_4_1 , config1_onehot_decoded_masks_4_2 , config1_onehot_decoded_masks_4_3 , config1_onehot_decoded_masks_4_4 ,
        config1_onehot_decoded_masks_4_5 , config1_onehot_decoded_masks_4_6 , config1_onehot_decoded_masks_4_7 , config1_onehot_decoded_masks_4_8 ,
        config1_onehot_decoded_masks_4_9 , config1_onehot_decoded_masks_4_10 , config1_onehot_decoded_masks_4_11 , config1_onehot_decoded_masks_4_12 ,
        config1_onehot_decoded_masks_4_13 , config1_onehot_decoded_masks_4_14 , config1_onehot_decoded_masks_4_15 , config1_onehot_decoded_masks_4_16 ,
        config1_onehot_decoded_masks_4_17 , config1_onehot_decoded_masks_4_18 , config1_onehot_decoded_masks_4_19 , config1_onehot_decoded_masks_4_20 ,
        config1_onehot_decoded_masks_4_21 , config1_onehot_decoded_masks_4_22 , config1_onehot_decoded_masks_4_23 , config1_onehot_decoded_masks_4_24 ,
        config1_onehot_decoded_masks_4_25 , config1_onehot_decoded_masks_4_26 , config1_onehot_decoded_masks_4_27 , config1_onehot_decoded_masks_4_28 ,
        config1_onehot_decoded_masks_4_29 , config1_onehot_decoded_masks_4_30 , config1_onehot_decoded_masks_4_31 , config1_onehot_decoded_masks_4_32 ,
        config1_onehot_decoded_masks_4_33 , config1_onehot_decoded_masks_4_34 , config1_onehot_decoded_masks_4_35 , config1_onehot_decoded_masks_4_36 ,
        config1_onehot_decoded_masks_4_37 , config1_onehot_decoded_masks_4_38 , config1_onehot_decoded_masks_4_39 , config1_onehot_decoded_masks_4_40 ,
        config1_onehot_decoded_masks_4_41 , config1_onehot_decoded_masks_4_42 , config1_onehot_decoded_masks_4_43 , config1_onehot_decoded_masks_4_44 ,
        config1_onehot_decoded_masks_4_45 , config1_onehot_decoded_masks_4_46 , config1_onehot_decoded_masks_4_47 , config1_onehot_decoded_masks_4_48 ,
        config1_onehot_decoded_masks_4_49 , config1_onehot_decoded_masks_4_50 , config1_onehot_decoded_masks_4_51 , config1_onehot_decoded_masks_4_52 ,
        config1_onehot_decoded_masks_4_53 , config1_onehot_decoded_masks_4_54 , config1_onehot_decoded_masks_4_55 , config1_onehot_decoded_masks_4_56 ,
        config1_onehot_decoded_masks_4_57 , config1_onehot_decoded_masks_4_58 , config1_onehot_decoded_masks_4_59 , config1_onehot_decoded_masks_4_60 ,
        config1_onehot_decoded_masks_4_61 , config1_onehot_decoded_masks_4_62 , config1_onehot_decoded_masks_4_63 , config1_onehot_decoded_masks_4_64 ,
        config1_onehot_decoded_masks_4_65 , config1_onehot_decoded_masks_4_66 , config1_onehot_decoded_masks_4_67 , config1_onehot_decoded_masks_4_68 ,
        config1_onehot_decoded_masks_4_69 , config1_onehot_decoded_masks_4_70 , config1_onehot_decoded_masks_4_71 , config1_onehot_decoded_masks_4_72 ,
        config1_onehot_decoded_masks_4_73 , config1_onehot_decoded_masks_4_74 , config1_onehot_decoded_masks_4_75 , config1_onehot_decoded_masks_4_76 ,
        config1_onehot_decoded_masks_4_77 , config1_onehot_decoded_masks_4_78 , config1_onehot_decoded_masks_4_79 , config1_onehot_decoded_masks_4_80 ,
        config1_onehot_decoded_masks_4_81 , config1_onehot_decoded_masks_4_82 , config1_onehot_decoded_masks_4_83 , config1_onehot_decoded_masks_4_84 ,
        config1_onehot_decoded_masks_4_85 , config1_onehot_decoded_masks_4_86 , config1_onehot_decoded_masks_4_87 , config1_onehot_decoded_masks_4_88 ,
        config1_onehot_decoded_masks_4_89 , config1_onehot_decoded_masks_4_90 , config1_onehot_decoded_masks_4_91 , config1_onehot_decoded_masks_4_92 ,
        config1_onehot_decoded_masks_4_93 , config1_onehot_decoded_masks_4_94 , config1_onehot_decoded_masks_4_95 , config1_onehot_decoded_masks_4_96 ,
        config1_onehot_decoded_masks_4_97 , config1_onehot_decoded_masks_4_98 , config1_onehot_decoded_masks_4_99 , config1_onehot_decoded_masks_4_100 ,
        config1_onehot_decoded_masks_4_101 , config1_onehot_decoded_masks_4_102 , config1_onehot_decoded_masks_4_103 , config1_onehot_decoded_masks_4_104 ,
        config1_onehot_decoded_masks_4_105 , masks_shift_reg_7_0 , masks_shift_reg_7_1 , masks_shift_reg_7_2 ,
        masks_shift_reg_7_3 , masks_shift_reg_7_4 , masks_shift_reg_7_5 , masks_shift_reg_7_6 ,
        masks_shift_reg_7_7 , masks_shift_reg_7_8 , masks_shift_reg_7_9 , masks_shift_reg_7_10 ,
        masks_shift_reg_4_0 , masks_shift_reg_4_1 , masks_shift_reg_4_2 , masks_shift_reg_4_3 ,
        masks_shift_reg_4_4 , masks_shift_reg_4_5 , masks_shift_reg_4_6 , masks_shift_reg_4_7 ,
        masks_shift_reg_4_8 , masks_shift_reg_4_9 , masks_shift_reg_4_10 , masks_shift_reg_2_0 ,
        masks_shift_reg_2_1 , masks_shift_reg_2_2 , masks_shift_reg_2_3 , masks_shift_reg_2_4 ,
        masks_shift_reg_2_5 , masks_shift_reg_2_6 , masks_shift_reg_2_7 , masks_shift_reg_2_8 ,
        masks_shift_reg_2_9 , masks_shift_reg_2_10 , masks_shift_reg_9_0 , masks_shift_reg_9_1 ,
        masks_shift_reg_9_2 , masks_shift_reg_9_3 , masks_shift_reg_9_4 , masks_shift_reg_9_5 ,
        masks_shift_reg_9_6 , masks_shift_reg_9_7 , masks_shift_reg_9_8 , masks_shift_reg_9_9 ,
        masks_shift_reg_9_10 , masks_shift_reg_3_0 , masks_shift_reg_3_1 , masks_shift_reg_3_2 ,
        masks_shift_reg_3_3 , masks_shift_reg_3_4 , masks_shift_reg_3_5 , masks_shift_reg_3_6 ,
        masks_shift_reg_3_7 , masks_shift_reg_3_8 , masks_shift_reg_3_9 , masks_shift_reg_3_10 ,
        masks_shift_reg_10_0 , masks_shift_reg_10_1 , masks_shift_reg_10_2 , masks_shift_reg_10_3 ,
        masks_shift_reg_10_4 , masks_shift_reg_10_5 , masks_shift_reg_10_6 , masks_shift_reg_10_7 ,
        masks_shift_reg_10_8 , masks_shift_reg_10_9 , masks_shift_reg_10_10 , masks_shift_reg_8_0 ,
        masks_shift_reg_8_1 , masks_shift_reg_8_2 , masks_shift_reg_8_3 , masks_shift_reg_8_4 ,
        masks_shift_reg_8_5 , masks_shift_reg_8_6 , masks_shift_reg_8_7 , masks_shift_reg_8_8 ,
        masks_shift_reg_8_9 , masks_shift_reg_8_10 , masks_shift_reg_5_0 , masks_shift_reg_5_1 ,
        masks_shift_reg_5_2 , masks_shift_reg_5_3 , masks_shift_reg_5_4 , masks_shift_reg_5_5 ,
        masks_shift_reg_5_6 , masks_shift_reg_5_7 , masks_shift_reg_5_8 , masks_shift_reg_5_9 ,
        masks_shift_reg_5_10 , masks_shift_reg_1_0 , masks_shift_reg_1_1 , masks_shift_reg_1_2 ,
        masks_shift_reg_1_3 , masks_shift_reg_1_4 , masks_shift_reg_1_5 , masks_shift_reg_1_6 ,
        masks_shift_reg_1_7 , masks_shift_reg_1_8 , masks_shift_reg_1_9 , masks_shift_reg_1_10 ,
        masks_shift_reg_12_0 , masks_shift_reg_12_1 , masks_shift_reg_12_2 , masks_shift_reg_12_3 ,
        masks_shift_reg_12_4 , masks_shift_reg_12_5 , masks_shift_reg_12_6 , masks_shift_reg_12_7 ,
        masks_shift_reg_12_8 , masks_shift_reg_12_9 , masks_shift_reg_12_10 , masks_shift_reg_6_0 ,
        masks_shift_reg_6_1 , masks_shift_reg_6_2 , masks_shift_reg_6_3 , masks_shift_reg_6_4 ,
        masks_shift_reg_6_5 , masks_shift_reg_6_6 , masks_shift_reg_6_7 , masks_shift_reg_6_8 ,
        masks_shift_reg_6_9 , masks_shift_reg_6_10 , masks_shift_reg_0_0 , masks_shift_reg_0_1 ,
        masks_shift_reg_0_2 , masks_shift_reg_0_3 , masks_shift_reg_0_4 , masks_shift_reg_0_5 ,
        masks_shift_reg_0_6 , masks_shift_reg_0_7 , masks_shift_reg_0_8 , masks_shift_reg_0_9 ,
        masks_shift_reg_0_10 , masks_shift_reg_13_0 , masks_shift_reg_13_1 , masks_shift_reg_13_2 ,
        masks_shift_reg_13_3 , masks_shift_reg_13_4 , masks_shift_reg_13_5 , masks_shift_reg_13_6 ,
        masks_shift_reg_13_7 , masks_shift_reg_11_0 , masks_shift_reg_11_1 , masks_shift_reg_11_2 ,
        masks_shift_reg_11_3 , masks_shift_reg_11_4 , masks_shift_reg_11_5 , masks_shift_reg_11_6 ,
        masks_shift_reg_11_7 , masks_shift_reg_11_8 , masks_shift_reg_11_9 , masks_shift_reg_11_10 ,
        constant_shift_controller_i.control_hold_reg_14_0 , constant_shift_controller_i.control_hold_reg_14_1 , constant_shift_controller_i.control_hold_reg_14_2 , constant_shift_controller_i.control_hold_reg_14_3 ,
        constant_shift_controller_i.control_hold_reg_14_4 , constant_shift_controller_i.control_hold_reg_14_5 , constant_shift_controller_i.control_hold_reg_14_6 , constant_shift_controller_i.control_hold_reg_13_0 ,
        constant_shift_controller_i.control_hold_reg_13_1 , constant_shift_controller_i.control_hold_reg_13_2 , constant_shift_controller_i.control_hold_reg_13_3 , constant_shift_controller_i.control_hold_reg_13_4 ,
        constant_shift_controller_i.control_hold_reg_13_5 , constant_shift_controller_i.control_hold_reg_13_6 , constant_shift_controller_i.control_hold_reg_13_7 , constant_shift_controller_i.control_hold_reg_12_0 ,
        constant_shift_controller_i.control_hold_reg_12_1 , constant_shift_controller_i.control_hold_reg_12_2 , constant_shift_controller_i.control_hold_reg_12_3 , constant_shift_controller_i.control_hold_reg_12_4 ,
        constant_shift_controller_i.control_hold_reg_12_5 , constant_shift_controller_i.control_hold_reg_12_6 , constant_shift_controller_i.control_hold_reg_12_7 , constant_shift_controller_i.control_hold_reg_11_0 ,
        constant_shift_controller_i.control_hold_reg_11_1 , constant_shift_controller_i.control_hold_reg_11_2 , constant_shift_controller_i.control_hold_reg_11_3 , constant_shift_controller_i.control_hold_reg_11_4 ,
        constant_shift_controller_i.control_hold_reg_11_5 , constant_shift_controller_i.control_hold_reg_11_6 , constant_shift_controller_i.control_hold_reg_11_7 , constant_shift_controller_i.control_hold_reg_10_0 ,
        constant_shift_controller_i.control_hold_reg_10_1 , constant_shift_controller_i.control_hold_reg_10_2 , constant_shift_controller_i.control_hold_reg_10_3 , constant_shift_controller_i.control_hold_reg_10_4 ,
        constant_shift_controller_i.control_hold_reg_10_5 , constant_shift_controller_i.control_hold_reg_10_6 , constant_shift_controller_i.control_hold_reg_10_7 , constant_shift_controller_i.control_hold_reg_9_0 ,
        constant_shift_controller_i.control_hold_reg_9_1 , constant_shift_controller_i.control_hold_reg_9_2 , constant_shift_controller_i.control_hold_reg_9_3 , constant_shift_controller_i.control_hold_reg_9_4 ,
        constant_shift_controller_i.control_hold_reg_9_5 , constant_shift_controller_i.control_hold_reg_9_6 , constant_shift_controller_i.control_hold_reg_9_7 , constant_shift_controller_i.control_hold_reg_8_0 ,
        constant_shift_controller_i.control_hold_reg_8_1 , constant_shift_controller_i.control_hold_reg_8_2 , constant_shift_controller_i.control_hold_reg_8_3 , constant_shift_controller_i.control_hold_reg_8_4 ,
        constant_shift_controller_i.control_hold_reg_8_5 , constant_shift_controller_i.control_hold_reg_8_6 , constant_shift_controller_i.control_hold_reg_8_7 , constant_shift_controller_i.control_hold_reg_7_0 ,
        constant_shift_controller_i.control_hold_reg_7_1 , constant_shift_controller_i.control_hold_reg_7_2 , constant_shift_controller_i.control_hold_reg_7_3 , constant_shift_controller_i.control_hold_reg_7_4 ,
        constant_shift_controller_i.control_hold_reg_7_5 , constant_shift_controller_i.control_hold_reg_7_6 , constant_shift_controller_i.control_hold_reg_7_7 , constant_shift_controller_i.control_hold_reg_6_0 ,
        constant_shift_controller_i.control_hold_reg_6_1 , constant_shift_controller_i.control_hold_reg_6_2 , constant_shift_controller_i.control_hold_reg_6_3 , constant_shift_controller_i.control_hold_reg_6_4 ,
        constant_shift_controller_i.control_hold_reg_6_5 , constant_shift_controller_i.control_hold_reg_6_6 , constant_shift_controller_i.control_hold_reg_6_7 , constant_shift_controller_i.control_hold_reg_5_0 ,
        constant_shift_controller_i.control_hold_reg_5_1 , constant_shift_controller_i.control_hold_reg_5_2 , constant_shift_controller_i.control_hold_reg_5_3 , constant_shift_controller_i.control_hold_reg_5_4 ,
        constant_shift_controller_i.control_hold_reg_5_5 , constant_shift_controller_i.control_hold_reg_5_6 , constant_shift_controller_i.control_hold_reg_5_7 , constant_shift_controller_i.control_hold_reg_4_0 ,
        constant_shift_controller_i.control_hold_reg_4_1 , constant_shift_controller_i.control_hold_reg_4_2 , constant_shift_controller_i.control_hold_reg_4_3 , constant_shift_controller_i.control_hold_reg_4_4 ,
        constant_shift_controller_i.control_hold_reg_4_5 , constant_shift_controller_i.control_hold_reg_4_6 , constant_shift_controller_i.control_hold_reg_4_7 , constant_shift_controller_i.control_hold_reg_3_0 ,
        constant_shift_controller_i.control_hold_reg_3_1 , constant_shift_controller_i.control_hold_reg_3_2 , constant_shift_controller_i.control_hold_reg_3_3 , constant_shift_controller_i.control_hold_reg_3_4 ,
        constant_shift_controller_i.control_hold_reg_3_5 , constant_shift_controller_i.control_hold_reg_3_6 , constant_shift_controller_i.control_hold_reg_3_7 , constant_shift_controller_i.control_hold_reg_2_0 ,
        constant_shift_controller_i.control_hold_reg_2_1 , constant_shift_controller_i.control_hold_reg_2_2 , constant_shift_controller_i.control_hold_reg_2_3 , constant_shift_controller_i.control_hold_reg_2_4 ,
        constant_shift_controller_i.control_hold_reg_2_5 , constant_shift_controller_i.control_hold_reg_2_6 , constant_shift_controller_i.control_hold_reg_2_7 , constant_shift_controller_i.control_hold_reg_1_0 ,
        constant_shift_controller_i.control_hold_reg_1_1 , constant_shift_controller_i.control_hold_reg_1_2 , constant_shift_controller_i.control_hold_reg_1_3 , constant_shift_controller_i.control_hold_reg_1_4 ,
        constant_shift_controller_i.control_hold_reg_1_5 , constant_shift_controller_i.control_hold_reg_1_6 , constant_shift_controller_i.control_hold_reg_1_7 , constant_shift_controller_i.control_hold_reg_0_0 ,
        constant_shift_controller_i.control_hold_reg_0_1 , constant_shift_controller_i.control_hold_reg_0_2 , constant_shift_controller_i.control_hold_reg_0_3 , constant_shift_controller_i.control_hold_reg_0_4 ,
        constant_shift_controller_i.control_hold_reg_0_5 , constant_shift_controller_i.control_hold_reg_0_6 , constant_shift_controller_i.control_hold_reg_0_7 , constant_shift_controller_i.bias_inputs_0 ,
        constant_shift_controller_i.bias_inputs_1 , constant_shift_controller_i.bias_inputs_2 , constant_shift_controller_i.bias_inputs_3 , constant_shift_controller_i.bias_inputs_4 ,
        constant_shift_controller_i.bias_inputs_5 , constant_shift_controller_i.bias_inputs_6 , constant_shift_controller_i.bias_inputs_7 , constant_shift_controller_i.bias_inputs_8 ,
        constant_shift_controller_i.bias_inputs_9 , constant_shift_controller_i.bias_inputs_10 , constant_shift_controller_i.bias_inputs_11 , constant_shift_controller_i.bias_inputs_12 ,
        constant_shift_controller_i.bias_inputs_13 , constant_shift_controller_i.bias_inputs_14 , constant_shift_controller_i.bias_inputs_15 , constant_shift_controller_i.bias_inputs_16 ,
        constant_shift_controller_i.bias_inputs_17 , constant_shift_controller_i.bias_inputs_18 , constant_shift_controller_i.bias_inputs_19 , constant_shift_controller_i.bias_inputs_20 ,
        constant_shift_controller_i.bias_inputs_21 , constant_shift_controller_i.bias_inputs_22 , constant_shift_controller_i.bias_inputs_23 , constant_shift_controller_i.bias_inputs_24 ,
        constant_shift_controller_i.bias_inputs_25 , constant_shift_controller_i.bias_inputs_26 , constant_shift_controller_i.bias_inputs_27 , constant_shift_controller_i.bias_inputs_28 ,
        constant_shift_controller_i.bias_inputs_29 , constant_shift_controller_i.bias_inputs_30 , constant_shift_controller_i.bias_inputs_31 , constant_shift_controller_i.bias_inputs_32 ,
        constant_shift_controller_i.bias_inputs_33 , constant_shift_controller_i.bias_inputs_34 , constant_shift_controller_i.bias_inputs_35 , constant_shift_controller_i.bias_inputs_36 ,
        constant_shift_controller_i.bias_inputs_37 , constant_shift_controller_i.bias_inputs_38 , constant_shift_controller_i.bias_inputs_39 , constant_shift_controller_i.bias_inputs_40 ,
        constant_shift_controller_i.bias_inputs_41 , constant_shift_controller_i.bias_inputs_42 , constant_shift_controller_i.bias_inputs_43 , constant_shift_controller_i.bias_inputs_44 ,
        constant_shift_controller_i.bias_inputs_45 , constant_shift_controller_i.bias_inputs_46 , constant_shift_controller_i.bias_inputs_47 , constant_shift_controller_i.bias_inputs_48 ,
        constant_shift_controller_i.bias_inputs_49 , constant_shift_controller_i.bias_inputs_50 , constant_shift_controller_i.bias_inputs_51 , constant_shift_controller_i.bias_inputs_52 ,
        constant_shift_controller_i.bias_inputs_53 , constant_shift_controller_i.bias_inputs_54 , constant_shift_controller_i.bias_inputs_55 , constant_shift_controller_i.bias_inputs_56 ,
        constant_shift_controller_i.bias_inputs_57 , constant_shift_controller_i.bias_inputs_58 , constant_shift_controller_i.bias_inputs_59 , constant_shift_controller_i.bias_inputs_60 ,
        constant_shift_controller_i.bias_inputs_61 , constant_shift_controller_i.bias_inputs_62 , constant_shift_controller_i.bias_inputs_63 , constant_shift_controller_i.bias_inputs_64 ,
        constant_shift_controller_i.bias_inputs_65 , constant_shift_controller_i.bias_inputs_66 , constant_shift_controller_i.bias_inputs_67 , constant_shift_controller_i.bias_inputs_68 ,
        constant_shift_controller_i.bias_inputs_69 , constant_shift_controller_i.bias_inputs_70 , constant_shift_controller_i.bias_inputs_71 , constant_shift_controller_i.bias_inputs_72 ,
        constant_shift_controller_i.bias_inputs_73 , constant_shift_controller_i.bias_inputs_74 , constant_shift_controller_i.bias_inputs_75 , constant_shift_controller_i.bias_inputs_76 ,
        constant_shift_controller_i.bias_inputs_77 , constant_shift_controller_i.bias_inputs_78 , constant_shift_controller_i.bias_inputs_79 , constant_shift_controller_i.bias_inputs_80 ,
        constant_shift_controller_i.bias_inputs_81 , constant_shift_controller_i.bias_inputs_82 , constant_shift_controller_i.bias_inputs_83 , constant_shift_controller_i.bias_inputs_84 ,
        constant_shift_controller_i.bias_inputs_85 , constant_shift_controller_i.bias_inputs_86 , constant_shift_controller_i.bias_inputs_87 , constant_shift_controller_i.bias_inputs_88 ,
        constant_shift_controller_i.bias_inputs_89 , constant_shift_controller_i.bias_inputs_90 , constant_shift_controller_i.bias_inputs_91 , constant_shift_controller_i.bias_inputs_92 ,
        constant_shift_controller_i.bias_inputs_93 , constant_shift_controller_i.bias_inputs_94 , constant_shift_controller_i.bias_inputs_95 , constant_shift_controller_i.bias_inputs_96 ,
        constant_shift_controller_i.bias_inputs_97 , constant_shift_controller_i.bias_inputs_98 , constant_shift_controller_i.bias_inputs_99 , constant_shift_controller_i.bias_inputs_100 ,
        constant_shift_controller_i.bias_inputs_101 , constant_shift_controller_i.bias_inputs_102 , constant_shift_controller_i.bias_inputs_103 , constant_shift_controller_i.bias_inputs_104 ,
        constant_shift_controller_i.bias_inputs_105 , constant_shift_controller_i.bias_inputs_106 , constant_shift_controller_i.bias_inputs_107 , constant_shift_controller_i.bias_inputs_108 ,
        constant_shift_controller_i.bias_inputs_109 , constant_shift_controller_i.bias_inputs_110 , constant_shift_controller_i.bias_inputs_111 , constant_shift_controller_i.bias_inputs_112 ,
        constant_shift_controller_i.bias_inputs_113 , constant_shift_controller_i.bias_inputs_114 , constant_shift_controller_i.bias_inputs_115 , constant_shift_controller_i.bias_inputs_116 ,
        constant_shift_controller_i.bias_inputs_117 , constant_shift_controller_i.bias_inputs_118 , constant_shift_controller_i.bias_inputs_119 , constant_shift_controller_i.bias_inputs_120 ,
        constant_shift_controller_i.bias_inputs_121 , constant_shift_controller_i.bias_inputs_122 , constant_shift_controller_i.bias_inputs_123 , constant_shift_controller_i.bias_inputs_124 ,
        constant_shift_controller_i.bias_inputs_125 , constant_shift_controller_i.bias_inputs_126 , constant_shift_controller_i.bias_inputs_127 , constant_shift_controller_i.bias_inputs_128 ,
        constant_shift_controller_i.bias_inputs_129 , constant_shift_controller_i.bias_inputs_130 , constant_shift_controller_i.bias_inputs_131 , constant_shift_controller_i.bias_inputs_132 ,
        constant_shift_controller_i.bias_inputs_133 , constant_shift_controller_i.bias_inputs_134 , constant_shift_controller_i.bias_inputs_135 , constant_shift_controller_i.bias_inputs_136 ,
        constant_shift_controller_i.bias_inputs_137 , constant_shift_controller_i.bias_inputs_138 , constant_shift_controller_i.bias_inputs_139 , constant_shift_controller_i.bias_inputs_140 ,
        constant_shift_controller_i.bias_inputs_141 , constant_shift_controller_i.bias_inputs_142 , constant_shift_controller_i.bias_inputs_143 , constant_shift_controller_i.bias_inputs_144 ,
        constant_shift_controller_i.bias_inputs_145 , constant_shift_controller_i.bias_inputs_146 , constant_shift_controller_i.bias_inputs_147 , constant_shift_controller_i.bias_inputs_148 ,
        constant_shift_controller_i.bias_inputs_149 , constant_shift_controller_i.bias_inputs_150 , constant_shift_controller_i.bias_inputs_151 , constant_shift_controller_i.bias_inputs_152 ,
        constant_shift_controller_i.bias_inputs_153 , constant_shift_controller_i.bias_inputs_154 , constant_shift_controller_i.bias_inputs_155 , constant_shift_controller_i.bias_inputs_156 ,
        constant_shift_controller_i.bias_inputs_157 , constant_shift_controller_i.bias_inputs_158 , constant_shift_controller_i.bias_inputs_159 , constant_shift_controller_i.bias_inputs_160 ,
        constant_shift_controller_i.bias_inputs_161 , constant_shift_controller_i.bias_inputs_162 , constant_shift_controller_i.bias_inputs_163 , constant_shift_controller_i.bias_inputs_164 ,
        constant_shift_controller_i.bias_inputs_165 , constant_shift_controller_i.bias_inputs_166 , constant_shift_controller_i.bias_inputs_167 , constant_shift_controller_i.bias_inputs_168 ,
        constant_shift_controller_i.bias_inputs_169 , constant_shift_controller_i.bias_inputs_170 , constant_shift_controller_i.bias_inputs_171 , constant_shift_controller_i.bias_inputs_172 ,
        constant_shift_controller_i.bias_inputs_173 , constant_shift_controller_i.bias_inputs_174 , constant_shift_controller_i.bias_inputs_175 , constant_shift_controller_i.bias_inputs_176 ,
        constant_shift_controller_i.bias_inputs_177 , constant_shift_controller_i.bias_inputs_178 , constant_shift_controller_i.bias_inputs_179 , constant_shift_controller_i.bias_inputs_180 ,
        constant_shift_controller_i.bias_inputs_181 , constant_shift_controller_i.bias_inputs_182 , constant_shift_controller_i.bias_inputs_183 , constant_shift_controller_i.bias_inputs_184 ,
        constant_shift_controller_i.bias_inputs_185 , constant_shift_controller_i.bias_inputs_186 , constant_shift_controller_i.bias_inputs_187 , constant_shift_controller_i.bias_inputs_188 ,
        constant_shift_controller_i.bias_inputs_189 , constant_shift_controller_i.bias_inputs_190 , constant_shift_controller_i.bias_inputs_191 , constant_shift_controller_i.bias_inputs_192 ,
        constant_shift_controller_i.bias_inputs_193 , constant_shift_controller_i.bias_inputs_194 , constant_shift_controller_i.bias_inputs_195 , constant_shift_controller_i.bias_inputs_196 ,
        constant_shift_controller_i.bias_inputs_197 , constant_shift_controller_i.bias_inputs_198 , constant_shift_controller_i.bias_inputs_199 , constant_shift_controller_i.bias_inputs_200 ,
        constant_shift_controller_i.bias_inputs_201 , constant_shift_controller_i.bias_inputs_202 , constant_shift_controller_i.bias_inputs_203 , constant_shift_controller_i.bias_inputs_204 ,
        constant_shift_controller_i.bias_inputs_205 , constant_shift_controller_i.bias_inputs_206 , constant_shift_controller_i.bias_inputs_207 , constant_shift_controller_i.bias_inputs_208 ,
        constant_shift_controller_i.bias_inputs_209 , constant_shift_controller_i.bias_inputs_210 , constant_shift_controller_i.bias_inputs_211 , constant_shift_controller_i.bias_inputs_212 ,
        constant_shift_controller_i.bias_inputs_213 , constant_shift_controller_i.bias_inputs_214 , constant_shift_controller_i.bias_inputs_215 , constant_shift_controller_i.bias_inputs_216 ,
        constant_shift_controller_i.bias_inputs_217 , constant_shift_controller_i.bias_inputs_218 , constant_shift_controller_i.bias_inputs_219 , constant_shift_controller_i.bias_inputs_220 ,
        constant_shift_controller_i.bias_inputs_221 , constant_shift_controller_i.bias_inputs_222 , constant_shift_controller_i.bias_inputs_223 , constant_shift_controller_i.bias_inputs_224 ,
        constant_shift_controller_i.bias_inputs_225 , constant_shift_controller_i.bias_inputs_226 , constant_shift_controller_i.bias_inputs_227 , constant_shift_controller_i.bias_inputs_228 ,
        constant_shift_controller_i.bias_inputs_229 , constant_shift_controller_i.bias_inputs_230 , constant_shift_controller_i.bias_inputs_231 , constant_shift_controller_i.bias_inputs_232 ,
        constant_shift_controller_i.bias_inputs_233 , constant_shift_controller_i.bias_inputs_234 , constant_shift_controller_i.bias_inputs_235 , constant_shift_controller_i.bias_inputs_236 ,
        constant_shift_controller_i.bias_inputs_237 , constant_shift_controller_i.bias_inputs_238 , constant_shift_controller_i.bias_inputs_239 , constant_shift_controller_i.bias_inputs_240 ,
        constant_shift_controller_i.bias_inputs_241 , constant_shift_controller_i.bias_inputs_242 , constant_shift_controller_i.bias_inputs_243 , constant_shift_controller_i.bias_inputs_244 ,
        constant_shift_controller_i.bias_inputs_245 , constant_shift_controller_i.bias_inputs_246 , constant_shift_controller_i.bias_inputs_247 , constant_shift_controller_i.bias_inputs_248 ,
        constant_shift_controller_i.bias_inputs_249 , constant_shift_controller_i.bias_inputs_250 , constant_shift_controller_i.bias_inputs_251 , constant_shift_controller_i.bias_inputs_252 ,
        constant_shift_controller_i.bias_inputs_253 , constant_shift_controller_i.bias_inputs_254 , constant_shift_controller_i.bias_inputs_255 , constant_shift_controller_i.bias_inputs_256 ,
        constant_shift_controller_i.bias_inputs_257 , constant_shift_controller_i.bias_inputs_258 , constant_shift_controller_i.bias_inputs_259 , constant_shift_controller_i.bias_inputs_260 ,
        constant_shift_controller_i.bias_inputs_261 , constant_shift_controller_i.bias_inputs_262 , constant_shift_controller_i.bias_inputs_263 , constant_shift_controller_i.bias_inputs_264 ,
        constant_shift_controller_i.bias_inputs_265 , constant_shift_controller_i.bias_inputs_266 , constant_shift_controller_i.bias_inputs_267 , constant_shift_controller_i.bias_inputs_268 ,
        constant_shift_controller_i.bias_inputs_269 , constant_shift_controller_i.bias_inputs_270 , constant_shift_controller_i.bias_inputs_271 , constant_shift_controller_i.bias_inputs_272 ,
        constant_shift_controller_i.bias_inputs_273 , constant_shift_controller_i.bias_inputs_274 , constant_shift_controller_i.bias_inputs_275 , constant_shift_controller_i.bias_inputs_276 ,
        constant_shift_controller_i.bias_inputs_277 , constant_shift_controller_i.bias_inputs_278 , constant_shift_controller_i.bias_inputs_279 , constant_shift_controller_i.bias_inputs_280 ,
        constant_shift_controller_i.bias_inputs_281 , constant_shift_controller_i.bias_inputs_282 , constant_shift_controller_i.bias_inputs_283 , constant_shift_controller_i.bias_inputs_284 ,
        constant_shift_controller_i.bias_inputs_285 , constant_shift_controller_i.bias_inputs_286 , constant_shift_controller_i.bias_inputs_287 , constant_shift_controller_i.bias_inputs_288 ,
        constant_shift_controller_i.bias_inputs_289 , constant_shift_controller_i.bias_inputs_290 , constant_shift_controller_i.bias_inputs_291 , constant_shift_controller_i.bias_inputs_292 ,
        constant_shift_controller_i.bias_inputs_293 , constant_shift_controller_i.bias_inputs_294 , constant_shift_controller_i.bias_inputs_295 , constant_shift_controller_i.bias_inputs_296 ,
        constant_shift_controller_i.bias_inputs_297 , constant_shift_controller_i.bias_inputs_298 , constant_shift_controller_i.bias_inputs_299 , constant_shift_controller_i.bias_inputs_300 ,
        constant_shift_controller_i.bias_inputs_301 , constant_shift_controller_i.bias_inputs_302 , constant_shift_controller_i.bias_inputs_303 , constant_shift_controller_i.bias_inputs_304 ,
        constant_shift_controller_i.bias_inputs_305 , constant_shift_controller_i.bias_inputs_306 , constant_shift_controller_i.bias_inputs_307 , constant_shift_controller_i.bias_inputs_308 ,
        constant_shift_controller_i.bias_inputs_309 , constant_shift_controller_i.bias_inputs_310 , constant_shift_controller_i.bias_inputs_311 , constant_shift_controller_i.bias_inputs_312 ,
        constant_shift_controller_i.bias_inputs_313 , constant_shift_controller_i.bias_inputs_314 , constant_shift_controller_i.bias_inputs_315 , constant_shift_controller_i.bias_inputs_316 ,
        constant_shift_controller_i.bias_inputs_317 , constant_shift_controller_i.bias_inputs_318 , constant_shift_controller_i.bias_inputs_319 , constant_shift_controller_i.bias_inputs_320 ,
        constant_shift_controller_i.bias_inputs_321 , constant_shift_controller_i.bias_inputs_322 , constant_shift_controller_i.bias_inputs_323 , constant_shift_controller_i.bias_inputs_324 ,
        constant_shift_controller_i.bias_inputs_325 , constant_shift_controller_i.bias_inputs_326 , constant_shift_controller_i.bias_inputs_327 , constant_shift_controller_i.bias_inputs_328 ,
        constant_shift_controller_i.bias_inputs_329 , constant_shift_controller_i.bias_inputs_330 , constant_shift_controller_i.bias_inputs_331 , constant_shift_controller_i.bias_inputs_332 ,
        constant_shift_controller_i.bias_inputs_333 , constant_shift_controller_i.bias_inputs_334 , constant_shift_controller_i.bias_inputs_335 , constant_shift_controller_i.bias_inputs_336 ,
        constant_shift_controller_i.bias_inputs_337 , constant_shift_controller_i.bias_inputs_338 , constant_shift_controller_i.bias_inputs_339 , constant_shift_controller_i.bias_inputs_340 ,
        constant_shift_controller_i.bias_inputs_341 , constant_shift_controller_i.bias_inputs_342 , constant_shift_controller_i.bias_inputs_343 , constant_shift_controller_i.bias_inputs_344 ,
        constant_shift_controller_i.bias_inputs_345 , constant_shift_controller_i.bias_inputs_346 , constant_shift_controller_i.bias_inputs_347 , constant_shift_controller_i.bias_inputs_348 ,
        constant_shift_controller_i.bias_inputs_349 , constant_shift_controller_i.bias_inputs_350 , constant_shift_controller_i.bias_inputs_351 , constant_shift_controller_i.bias_inputs_352 ,
        constant_shift_controller_i.bias_inputs_353 , constant_shift_controller_i.bias_inputs_354 , constant_shift_controller_i.bias_inputs_355 , constant_shift_controller_i.bias_inputs_356 ,
        constant_shift_controller_i.bias_inputs_357 , constant_shift_controller_i.bias_inputs_358 , constant_shift_controller_i.bias_inputs_359 , constant_shift_controller_i.bias_inputs_360 ,
        constant_shift_controller_i.bias_inputs_361 , constant_shift_controller_i.bias_inputs_362 , constant_shift_controller_i.bias_inputs_363 , constant_shift_controller_i.bias_inputs_364 ,
        constant_shift_controller_i.bias_inputs_365 , constant_shift_controller_i.bias_inputs_366 , constant_shift_controller_i.bias_inputs_367 , constant_shift_controller_i.bias_inputs_368 ,
        constant_shift_controller_i.bias_inputs_369 , constant_shift_controller_i.bias_inputs_370 , constant_shift_controller_i.bias_inputs_371 , constant_shift_controller_i.bias_inputs_372 ,
        constant_shift_controller_i.bias_inputs_373 , constant_shift_controller_i.bias_inputs_374 , constant_shift_controller_i.bias_inputs_375 , constant_shift_controller_i.bias_inputs_376 ,
        constant_shift_controller_i.bias_inputs_377 , constant_shift_controller_i.bias_inputs_378 , constant_shift_controller_i.bias_inputs_379 , constant_shift_controller_i.bias_inputs_380 ,
        constant_shift_controller_i.bias_inputs_381 , constant_shift_controller_i.bias_inputs_382 , constant_shift_controller_i.bias_inputs_383 , constant_shift_controller_i.bias_inputs_384 ,
        constant_shift_controller_i.bias_inputs_385 , constant_shift_controller_i.bias_inputs_386 , constant_shift_controller_i.bias_inputs_387 , constant_shift_controller_i.bias_inputs_388 ,
        constant_shift_controller_i.bias_inputs_389 , constant_shift_controller_i.bias_inputs_390 , constant_shift_controller_i.bias_inputs_391 , constant_shift_controller_i.bias_inputs_392 ,
        constant_shift_controller_i.bias_inputs_393 , constant_shift_controller_i.bias_inputs_394 , constant_shift_controller_i.bias_inputs_395 , constant_shift_controller_i.bias_inputs_396 ,
        constant_shift_controller_i.bias_inputs_397 , constant_shift_controller_i.bias_inputs_398 , constant_shift_controller_i.bias_inputs_399 , constant_shift_controller_i.bias_inputs_400 ,
        constant_shift_controller_i.bias_inputs_401 , constant_shift_controller_i.bias_inputs_402 , constant_shift_controller_i.bias_inputs_403 , constant_shift_controller_i.bias_inputs_404 ,
        constant_shift_controller_i.bias_inputs_405 , constant_shift_controller_i.bias_inputs_406 , constant_shift_controller_i.bias_inputs_407 , constant_shift_controller_i.bias_inputs_408 ,
        constant_shift_controller_i.bias_inputs_409 , constant_shift_controller_i.bias_inputs_410 , constant_shift_controller_i.bias_inputs_411 , constant_shift_controller_i.bias_inputs_412 ,
        constant_shift_controller_i.bias_inputs_413 , constant_shift_controller_i.bias_inputs_414 , constant_shift_controller_i.bias_inputs_415 , constant_shift_controller_i.bias_inputs_416 ,
        constant_shift_controller_i.bias_inputs_417 , constant_shift_controller_i.bias_inputs_418 , constant_shift_controller_i.bias_inputs_419 , constant_shift_controller_i.bias_inputs_420 ,
        constant_shift_controller_i.bias_inputs_421 , constant_shift_controller_i.bias_inputs_422 , constant_shift_controller_i.bias_inputs_423 , constant_shift_controller_i.bias_inputs_424 ,
        constant_shift_controller_i.bias_inputs_425 , constant_shift_controller_i.bias_inputs_426 , constant_shift_controller_i.bias_inputs_427 , constant_shift_controller_i.bias_inputs_428 ,
        constant_shift_controller_i.bias_inputs_429 , constant_shift_controller_i.bias_inputs_430 , constant_shift_controller_i.bias_inputs_431 , constant_shift_controller_i.bias_inputs_432 ,
        constant_shift_controller_i.bias_inputs_433 , constant_shift_controller_i.bias_inputs_434 , constant_shift_controller_i.bias_inputs_435 , constant_shift_controller_i.bias_inputs_436 ,
        constant_shift_controller_i.bias_inputs_437 , constant_shift_controller_i.bias_inputs_438 , constant_shift_controller_i.bias_inputs_439 , constant_shift_controller_i.bias_inputs_440 ,
        constant_shift_controller_i.bias_inputs_441 , constant_shift_controller_i.bias_inputs_442 , constant_shift_controller_i.bias_inputs_443 , constant_shift_controller_i.bias_inputs_444 ,
        constant_shift_controller_i.bias_inputs_445 , constant_shift_controller_i.bias_inputs_446 , constant_shift_controller_i.bias_inputs_447 , constant_shift_controller_i.bias_inputs_448 ,
        constant_shift_controller_i.bias_inputs_449 , constant_shift_controller_i.bias_inputs_450 , constant_shift_controller_i.bias_inputs_451 , constant_shift_controller_i.bias_inputs_452 ,
        constant_shift_controller_i.bias_inputs_453 , constant_shift_controller_i.bias_inputs_454 , constant_shift_controller_i.bias_inputs_455 , constant_shift_controller_i.bias_inputs_456 ,
        constant_shift_controller_i.bias_inputs_457 , constant_shift_controller_i.bias_inputs_458 , constant_shift_controller_i.bias_inputs_459 , constant_shift_controller_i.bias_inputs_460 ,
        constant_shift_controller_i.bias_inputs_461 , constant_shift_controller_i.bias_inputs_462 , constant_shift_controller_i.bias_inputs_463 , constant_shift_controller_i.bias_inputs_464 ,
        constant_shift_controller_i.bias_inputs_465 , constant_shift_controller_i.bias_inputs_466 , constant_shift_controller_i.bias_inputs_467 , constant_shift_controller_i.bias_inputs_468 ,
        constant_shift_controller_i.bias_inputs_469 , constant_shift_controller_i.bias_inputs_470 , constant_shift_controller_i.bias_inputs_471 , constant_shift_controller_i.bias_inputs_472 ,
        constant_shift_controller_i.bias_inputs_473 , constant_shift_controller_i.bias_inputs_474 , constant_shift_controller_i.bias_inputs_475 , constant_shift_controller_i.bias_inputs_476 ,
        constant_shift_controller_i.bias_inputs_477 , constant_shift_controller_i.bias_inputs_478 , constant_shift_controller_i.bias_inputs_479 , constant_shift_controller_i.bias_inputs_480 ,
        constant_shift_controller_i.bias_inputs_481 , constant_shift_controller_i.bias_inputs_482 , constant_shift_controller_i.bias_inputs_483 , constant_shift_controller_i.bias_inputs_484 ,
        constant_shift_controller_i.bias_inputs_485 , constant_shift_controller_i.bias_inputs_486 , constant_shift_controller_i.bias_inputs_487 , constant_shift_controller_i.bias_inputs_488 ,
        constant_shift_controller_i.bias_inputs_489 , constant_shift_controller_i.bias_inputs_490 , constant_shift_controller_i.bias_inputs_491 , constant_shift_controller_i.bias_inputs_492 ,
        constant_shift_controller_i.bias_inputs_493 , constant_shift_controller_i.bias_inputs_494 , constant_shift_controller_i.bias_inputs_495 , constant_shift_controller_i.bias_inputs_496 ,
        constant_shift_controller_i.bias_inputs_497 , constant_shift_controller_i.bias_inputs_498 , constant_shift_controller_i.bias_inputs_499 , constant_shift_controller_i.bias_inputs_500 ,
        constant_shift_controller_i.bias_inputs_501 , constant_shift_controller_i.bias_inputs_502 , constant_shift_controller_i.bias_inputs_503 , constant_shift_controller_i.bias_inputs_504 ,
        constant_shift_controller_i.bias_inputs_505 , constant_shift_controller_i.bias_inputs_506 , constant_shift_controller_i.bias_inputs_507 , constant_shift_controller_i.bias_inputs_508 ,
        constant_shift_controller_i.bias_inputs_509 , constant_shift_controller_i.bias_inputs_510 , constant_shift_controller_i.bias_inputs_511 , constant_shift_controller_i.bias_inputs_512 ,
        constant_shift_controller_i.bias_inputs_513 , constant_shift_controller_i.bias_inputs_514 , constant_shift_controller_i.bias_inputs_515 , constant_shift_controller_i.bias_inputs_516 ,
        constant_shift_controller_i.bias_inputs_517 , constant_shift_controller_i.bias_inputs_518 , constant_shift_controller_i.bias_inputs_519 , constant_shift_controller_i.bias_inputs_520 ,
        constant_shift_controller_i.bias_inputs_521 , constant_shift_controller_i.bias_inputs_522 , constant_shift_controller_i.bias_inputs_523 , constant_shift_controller_i.bias_inputs_524 ,
        constant_shift_controller_i.bias_inputs_525 , constant_shift_controller_i.bias_inputs_526 , constant_shift_controller_i.bias_inputs_527 , constant_shift_controller_i.bias_inputs_528 ,
        constant_shift_controller_i.bias_inputs_529 , constant_shift_controller_i.bias_inputs_530 , constant_shift_controller_i.bias_inputs_531 , constant_shift_controller_i.bias_inputs_532 ,
        constant_shift_controller_i.bias_inputs_533 , constant_shift_controller_i.bias_inputs_534 , constant_shift_controller_i.bias_inputs_535 , constant_shift_controller_i.bias_inputs_536 ,
        constant_shift_controller_i.bias_inputs_537 , constant_shift_controller_i.bias_inputs_538 , constant_shift_controller_i.bias_inputs_539 , constant_shift_controller_i.bias_inputs_540 ,
        constant_shift_controller_i.bias_inputs_541 , constant_shift_controller_i.bias_inputs_542 , constant_shift_controller_i.bias_inputs_543 , constant_shift_controller_i.bias_inputs_544 ,
        constant_shift_controller_i.bias_inputs_545 , constant_shift_controller_i.bias_inputs_546 , constant_shift_controller_i.bias_inputs_547 , constant_shift_controller_i.bias_inputs_548 ,
        constant_shift_controller_i.bias_inputs_549 , constant_shift_controller_i.bias_inputs_550 , constant_shift_controller_i.bias_inputs_551 , constant_shift_controller_i.bias_inputs_552 ,
        constant_shift_controller_i.bias_inputs_553 , constant_shift_controller_i.bias_inputs_554 , constant_shift_controller_i.bias_inputs_555 , constant_shift_controller_i.bias_inputs_556 ,
        constant_shift_controller_i.bias_inputs_557 , constant_shift_controller_i.bias_inputs_558 , constant_shift_controller_i.bias_inputs_559 , constant_shift_controller_i.bias_inputs_560 ,
        constant_shift_controller_i.bias_inputs_561 , constant_shift_controller_i.bias_inputs_562 , constant_shift_controller_i.bias_inputs_563 , constant_shift_controller_i.bias_inputs_564 ,
        constant_shift_controller_i.bias_inputs_565 , constant_shift_controller_i.bias_inputs_566 , constant_shift_controller_i.bias_inputs_567 , constant_shift_controller_i.bias_inputs_568 ,
        constant_shift_controller_i.bias_inputs_569 , constant_shift_controller_i.bias_inputs_570 , constant_shift_controller_i.bias_inputs_571 , constant_shift_controller_i.bias_inputs_572 ,
        constant_shift_controller_i.bias_inputs_573 , constant_shift_controller_i.bias_inputs_574 , constant_shift_controller_i.bias_inputs_575 , constant_shift_controller_i.bias_inputs_576 ,
        constant_shift_controller_i.bias_inputs_577 , constant_shift_controller_i.bias_inputs_578 , constant_shift_controller_i.bias_inputs_579 , constant_shift_controller_i.bias_inputs_580 ,
        constant_shift_controller_i.bias_inputs_581 , constant_shift_controller_i.bias_inputs_582 , constant_shift_controller_i.bias_inputs_583 , constant_shift_controller_i.bias_inputs_584 ,
        constant_shift_controller_i.bias_inputs_585 , constant_shift_controller_i.bias_inputs_586 , constant_shift_controller_i.bias_inputs_587 , constant_shift_controller_i.bias_inputs_588 ,
        constant_shift_controller_i.bias_inputs_589 , constant_shift_controller_i.bias_inputs_590 , constant_shift_controller_i.bias_inputs_591 , constant_shift_controller_i.bias_inputs_592 ,
        constant_shift_controller_i.bias_inputs_593 , constant_shift_controller_i.bias_inputs_594 , constant_shift_controller_i.bias_inputs_595 , constant_shift_controller_i.bias_inputs_596 ,
        constant_shift_controller_i.bias_inputs_597 , constant_shift_controller_i.bias_inputs_598 , constant_shift_controller_i.bias_inputs_599 , constant_shift_controller_i.bias_inputs_600 ,
        constant_shift_controller_i.bias_inputs_601 , constant_shift_controller_i.bias_inputs_602 , constant_shift_controller_i.bias_inputs_603 , constant_shift_controller_i.bias_inputs_604 ,
        constant_shift_controller_i.bias_inputs_605 , constant_shift_controller_i.bias_inputs_606 , constant_shift_controller_i.bias_inputs_607 , constant_shift_controller_i.bias_inputs_608 ,
        constant_shift_controller_i.bias_inputs_609 , constant_shift_controller_i.bias_inputs_610 , constant_shift_controller_i.bias_inputs_611 , constant_shift_controller_i.bias_inputs_612 ,
        constant_shift_controller_i.bias_inputs_613 , constant_shift_controller_i.bias_inputs_614 , constant_shift_controller_i.bias_inputs_615 , constant_shift_controller_i.bias_inputs_616 ,
        constant_shift_controller_i.bias_inputs_617 , constant_shift_controller_i.bias_inputs_618 , constant_shift_controller_i.bias_inputs_619 , constant_shift_controller_i.bias_inputs_620 ,
        constant_shift_controller_i.bias_inputs_621 , constant_shift_controller_i.bias_inputs_622 , constant_shift_controller_i.bias_inputs_623 , constant_shift_controller_i.bias_inputs_624 ,
        constant_shift_controller_i.bias_inputs_625 , constant_shift_controller_i.bias_inputs_626 , constant_shift_controller_i.bias_inputs_627 , constant_shift_controller_i.bias_inputs_628 ,
        constant_shift_controller_i.bias_inputs_629 , constant_shift_controller_i.bias_inputs_630 , constant_shift_controller_i.bias_inputs_631 , constant_shift_controller_i.bias_inputs_632 ,
        constant_shift_controller_i.bias_inputs_633 , constant_shift_controller_i.bias_inputs_634 , constant_shift_controller_i.bias_inputs_635 , constant_shift_controller_i.bias_inputs_636 ,
        constant_shift_controller_i.bias_inputs_637 , constant_shift_controller_i.bias_inputs_638 , constant_shift_controller_i.bias_inputs_639 , constant_shift_controller_i.bias_inputs_640 ,
        constant_shift_controller_i.bias_inputs_641 , constant_shift_controller_i.bias_inputs_642 , constant_shift_controller_i.bias_inputs_643 , constant_shift_controller_i.bias_inputs_644 ,
        constant_shift_controller_i.bias_inputs_645 , constant_shift_controller_i.bias_inputs_646 , constant_shift_controller_i.bias_inputs_647 , constant_shift_controller_i.bias_inputs_648 ,
        constant_shift_controller_i.bias_inputs_649 , constant_shift_controller_i.bias_inputs_650 , constant_shift_controller_i.bias_inputs_651 , constant_shift_controller_i.bias_inputs_652 ,
        constant_shift_controller_i.bias_inputs_653 , constant_shift_controller_i.bias_inputs_654 , constant_shift_controller_i.bias_inputs_655 , constant_shift_controller_i.bias_inputs_656 ,
        constant_shift_controller_i.bias_inputs_657 , constant_shift_controller_i.bias_inputs_658 , constant_shift_controller_i.bias_inputs_659 , constant_shift_controller_i.bias_inputs_660 ,
        constant_shift_controller_i.bias_inputs_661 , constant_shift_controller_i.bias_inputs_662 , constant_shift_controller_i.bias_inputs_663 , constant_shift_controller_i.bias_inputs_664 ,
        constant_shift_controller_i.bias_inputs_665 , constant_shift_controller_i.bias_inputs_666 , constant_shift_controller_i.bias_inputs_667 , constant_shift_controller_i.bias_inputs_668 ,
        constant_shift_controller_i.bias_inputs_669 , constant_shift_controller_i.bias_inputs_670 , constant_shift_controller_i.bias_inputs_671 , constant_shift_controller_i.bias_inputs_672 ,
        constant_shift_controller_i.bias_inputs_673 , constant_shift_controller_i.bias_inputs_674 , constant_shift_controller_i.bias_inputs_675 , constant_shift_controller_i.bias_inputs_676 ,
        constant_shift_controller_i.bias_inputs_677 , constant_shift_controller_i.bias_inputs_678 , constant_shift_controller_i.bias_inputs_679 , constant_shift_controller_i.bias_inputs_680 ,
        constant_shift_controller_i.bias_inputs_681 , constant_shift_controller_i.bias_inputs_682 , constant_shift_controller_i.bias_inputs_683 , constant_shift_controller_i.bias_inputs_684 ,
        constant_shift_controller_i.bias_inputs_685 , constant_shift_controller_i.bias_inputs_686 , constant_shift_controller_i.bias_inputs_687 , constant_shift_controller_i.bias_inputs_688 ,
        constant_shift_controller_i.bias_inputs_689 , constant_shift_controller_i.bias_inputs_690 , constant_shift_controller_i.bias_inputs_691 , constant_shift_controller_i.bias_inputs_692 ,
        constant_shift_controller_i.bias_inputs_693 , constant_shift_controller_i.bias_inputs_694 , constant_shift_controller_i.bias_inputs_695 , constant_shift_controller_i.bias_inputs_696 ,
        constant_shift_controller_i.bias_inputs_697 , constant_shift_controller_i.bias_inputs_698 , constant_shift_controller_i.bias_inputs_699 , constant_shift_controller_i.bias_inputs_700 ,
        constant_shift_controller_i.bias_inputs_701 , constant_shift_controller_i.bias_inputs_702 , constant_shift_controller_i.bias_inputs_703 , constant_shift_controller_i.bias_inputs_704 ,
        constant_shift_controller_i.bias_inputs_705 , constant_shift_controller_i.bias_inputs_706 , constant_shift_controller_i.bias_inputs_707 , constant_shift_controller_i.bias_inputs_708 ,
        constant_shift_controller_i.bias_inputs_709 , constant_shift_controller_i.bias_inputs_710 , constant_shift_controller_i.bias_inputs_711 , constant_shift_controller_i.bias_inputs_712 ,
        constant_shift_controller_i.bias_inputs_713 , constant_shift_controller_i.bias_inputs_714 , constant_shift_controller_i.bias_inputs_715 , constant_shift_controller_i.bias_inputs_716 ,
        constant_shift_controller_i.bias_inputs_717 , constant_shift_controller_i.bias_inputs_718 , constant_shift_controller_i.bias_inputs_719 , constant_shift_controller_i.bias_inputs_720 ,
        constant_shift_controller_i.bias_inputs_721 , constant_shift_controller_i.bias_inputs_722 , constant_shift_controller_i.bias_inputs_723 , constant_shift_controller_i.bias_inputs_724 ,
        constant_shift_controller_i.bias_inputs_725 , constant_shift_controller_i.bias_inputs_726 , constant_shift_controller_i.bias_inputs_727 , constant_shift_controller_i.bias_inputs_728 ,
        constant_shift_controller_i.bias_inputs_729 , constant_shift_controller_i.bias_inputs_730 , constant_shift_controller_i.bias_inputs_731 , constant_shift_controller_i.bias_inputs_732 ,
        constant_shift_controller_i.bias_inputs_733 , constant_shift_controller_i.bias_inputs_734 , constant_shift_controller_i.bias_inputs_735 , constant_shift_controller_i.bias_inputs_736 ,
        constant_shift_controller_i.bias_inputs_737 , constant_shift_controller_i.bias_inputs_738 , constant_shift_controller_i.bias_inputs_739 , constant_shift_controller_i.bias_inputs_740 ,
        constant_shift_controller_i.bias_inputs_741 , constant_shift_controller_i.bias_inputs_742 , constant_shift_controller_i.bias_inputs_743 , constant_shift_controller_i.bias_inputs_744 ,
        constant_shift_controller_i.bias_inputs_745 , constant_shift_controller_i.bias_inputs_746 , constant_shift_controller_i.bias_inputs_747 , constant_shift_controller_i.bias_inputs_748 ,
        constant_shift_controller_i.bias_inputs_749 , constant_shift_controller_i.bias_inputs_750 , constant_shift_controller_i.bias_inputs_751 , constant_shift_controller_i.bias_inputs_752 ,
        constant_shift_controller_i.bias_inputs_753 , constant_shift_controller_i.bias_inputs_754 , constant_shift_controller_i.bias_inputs_755 , constant_shift_controller_i.bias_inputs_756 ,
        constant_shift_controller_i.bias_inputs_757 , constant_shift_controller_i.bias_inputs_758 , constant_shift_controller_i.bias_inputs_759 , constant_shift_controller_i.bias_inputs_760 ,
        constant_shift_controller_i.bias_inputs_761 , constant_shift_controller_i.bias_inputs_762 , constant_shift_controller_i.bias_inputs_763 , constant_shift_controller_i.bias_inputs_764 ,
        constant_shift_controller_i.bias_inputs_765 , constant_shift_controller_i.bias_inputs_766 , constant_shift_controller_i.bias_inputs_767 , constant_shift_controller_i.bias_inputs_768 ,
        constant_shift_controller_i.bias_inputs_769 , constant_shift_controller_i.bias_inputs_770 , constant_shift_controller_i.bias_inputs_771 , constant_shift_controller_i.bias_inputs_772 ,
        constant_shift_controller_i.bias_inputs_773 , constant_shift_controller_i.bias_inputs_774 , constant_shift_controller_i.bias_inputs_775 , constant_shift_controller_i.bias_inputs_776 ,
        constant_shift_controller_i.bias_inputs_777 , constant_shift_controller_i.bias_inputs_778 , constant_shift_controller_i.bias_inputs_779 , constant_shift_controller_i.bias_inputs_780 ,
        constant_shift_controller_i.bias_inputs_781 , constant_shift_controller_i.bias_inputs_782 , constant_shift_controller_i.bias_inputs_783 , constant_shift_controller_i.bias_inputs_784 ,
        constant_shift_controller_i.bias_inputs_785 , constant_shift_controller_i.bias_inputs_786 , constant_shift_controller_i.bias_inputs_787 , constant_shift_controller_i.bias_inputs_788 ,
        constant_shift_controller_i.bias_inputs_789 , constant_shift_controller_i.bias_inputs_790 , constant_shift_controller_i.bias_inputs_791 , constant_shift_controller_i.bias_inputs_792 ,
        constant_shift_controller_i.bias_inputs_793 , constant_shift_controller_i.bias_inputs_794 , constant_shift_controller_i.bias_inputs_795 , constant_shift_controller_i.control_shift_reg_8_0 ,
        constant_shift_controller_i.control_shift_reg_8_1 , constant_shift_controller_i.control_shift_reg_8_2 , constant_shift_controller_i.control_shift_reg_8_3 , constant_shift_controller_i.control_shift_reg_8_4 ,
        constant_shift_controller_i.control_shift_reg_8_5 , constant_shift_controller_i.control_shift_reg_8_6 , constant_shift_controller_i.control_shift_reg_8_7 , constant_shift_controller_i.control_shift_reg_5_0 ,
        constant_shift_controller_i.control_shift_reg_5_1 , constant_shift_controller_i.control_shift_reg_5_2 , constant_shift_controller_i.control_shift_reg_5_3 , constant_shift_controller_i.control_shift_reg_5_4 ,
        constant_shift_controller_i.control_shift_reg_5_5 , constant_shift_controller_i.control_shift_reg_5_6 , constant_shift_controller_i.control_shift_reg_5_7 , constant_shift_controller_i.control_shift_reg_4_0 ,
        constant_shift_controller_i.control_shift_reg_4_1 , constant_shift_controller_i.control_shift_reg_4_2 , constant_shift_controller_i.control_shift_reg_4_3 , constant_shift_controller_i.control_shift_reg_4_4 ,
        constant_shift_controller_i.control_shift_reg_4_5 , constant_shift_controller_i.control_shift_reg_4_6 , constant_shift_controller_i.control_shift_reg_4_7 , constant_shift_controller_i.control_shift_reg_7_0 ,
        constant_shift_controller_i.control_shift_reg_7_1 , constant_shift_controller_i.control_shift_reg_7_2 , constant_shift_controller_i.control_shift_reg_7_3 , constant_shift_controller_i.control_shift_reg_7_4 ,
        constant_shift_controller_i.control_shift_reg_7_5 , constant_shift_controller_i.control_shift_reg_7_6 , constant_shift_controller_i.control_shift_reg_7_7 , constant_shift_controller_i.control_shift_reg_14_0 ,
        constant_shift_controller_i.control_shift_reg_14_1 , constant_shift_controller_i.control_shift_reg_14_2 , constant_shift_controller_i.control_shift_reg_14_3 , constant_shift_controller_i.control_shift_reg_14_4 ,
        constant_shift_controller_i.control_shift_reg_14_5 , constant_shift_controller_i.control_shift_reg_14_6 , constant_shift_controller_i.control_shift_reg_10_0 , constant_shift_controller_i.control_shift_reg_10_1 ,
        constant_shift_controller_i.control_shift_reg_10_2 , constant_shift_controller_i.control_shift_reg_10_3 , constant_shift_controller_i.control_shift_reg_10_4 , constant_shift_controller_i.control_shift_reg_10_5 ,
        constant_shift_controller_i.control_shift_reg_10_6 , constant_shift_controller_i.control_shift_reg_10_7 , constant_shift_controller_i.control_shift_reg_2_0 , constant_shift_controller_i.control_shift_reg_2_1 ,
        constant_shift_controller_i.control_shift_reg_2_2 , constant_shift_controller_i.control_shift_reg_2_3 , constant_shift_controller_i.control_shift_reg_2_4 , constant_shift_controller_i.control_shift_reg_2_5 ,
        constant_shift_controller_i.control_shift_reg_2_6 , constant_shift_controller_i.control_shift_reg_2_7 , constant_shift_controller_i.control_shift_reg_13_0 , constant_shift_controller_i.control_shift_reg_13_1 ,
        constant_shift_controller_i.control_shift_reg_13_2 , constant_shift_controller_i.control_shift_reg_13_3 , constant_shift_controller_i.control_shift_reg_13_4 , constant_shift_controller_i.control_shift_reg_13_5 ,
        constant_shift_controller_i.control_shift_reg_13_6 , constant_shift_controller_i.control_shift_reg_13_7 , constant_shift_controller_i.control_shift_reg_0_0 , constant_shift_controller_i.control_shift_reg_0_1 ,
        constant_shift_controller_i.control_shift_reg_0_2 , constant_shift_controller_i.control_shift_reg_0_3 , constant_shift_controller_i.control_shift_reg_0_4 , constant_shift_controller_i.control_shift_reg_0_5 ,
        constant_shift_controller_i.control_shift_reg_0_6 , constant_shift_controller_i.control_shift_reg_0_7 , constant_shift_controller_i.control_shift_reg_9_0 , constant_shift_controller_i.control_shift_reg_9_1 ,
        constant_shift_controller_i.control_shift_reg_9_2 , constant_shift_controller_i.control_shift_reg_9_3 , constant_shift_controller_i.control_shift_reg_9_4 , constant_shift_controller_i.control_shift_reg_9_5 ,
        constant_shift_controller_i.control_shift_reg_9_6 , constant_shift_controller_i.control_shift_reg_9_7 , constant_shift_controller_i.control_shift_reg_3_0 , constant_shift_controller_i.control_shift_reg_3_1 ,
        constant_shift_controller_i.control_shift_reg_3_2 , constant_shift_controller_i.control_shift_reg_3_3 , constant_shift_controller_i.control_shift_reg_3_4 , constant_shift_controller_i.control_shift_reg_3_5 ,
        constant_shift_controller_i.control_shift_reg_3_6 , constant_shift_controller_i.control_shift_reg_3_7 , constant_shift_controller_i.control_shift_reg_6_0 , constant_shift_controller_i.control_shift_reg_6_1 ,
        constant_shift_controller_i.control_shift_reg_6_2 , constant_shift_controller_i.control_shift_reg_6_3 , constant_shift_controller_i.control_shift_reg_6_4 , constant_shift_controller_i.control_shift_reg_6_5 ,
        constant_shift_controller_i.control_shift_reg_6_6 , constant_shift_controller_i.control_shift_reg_6_7 , constant_shift_controller_i.control_shift_reg_12_0 , constant_shift_controller_i.control_shift_reg_12_1 ,
        constant_shift_controller_i.control_shift_reg_12_2 , constant_shift_controller_i.control_shift_reg_12_3 , constant_shift_controller_i.control_shift_reg_12_4 , constant_shift_controller_i.control_shift_reg_12_5 ,
        constant_shift_controller_i.control_shift_reg_12_6 , constant_shift_controller_i.control_shift_reg_12_7 , constant_shift_controller_i.control_shift_reg_1_0 , constant_shift_controller_i.control_shift_reg_1_1 ,
        constant_shift_controller_i.control_shift_reg_1_2 , constant_shift_controller_i.control_shift_reg_1_3 , constant_shift_controller_i.control_shift_reg_1_4 , constant_shift_controller_i.control_shift_reg_1_5 ,
        constant_shift_controller_i.control_shift_reg_1_6 , constant_shift_controller_i.control_shift_reg_1_7 , constant_shift_controller_i.control_shift_reg_11_0 , constant_shift_controller_i.control_shift_reg_11_1 ,
        constant_shift_controller_i.control_shift_reg_11_2 , constant_shift_controller_i.control_shift_reg_11_3 , constant_shift_controller_i.control_shift_reg_11_4 , constant_shift_controller_i.control_shift_reg_11_5 ,
        constant_shift_controller_i.control_shift_reg_11_6 , constant_shift_controller_i.control_shift_reg_11_7 ;
or ( 
    .Z ( config0_decoder12.U28.AB ) ,
    .I0 ( config0_decoder12.n40 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
and ( 
    .Z ( config0_decoder12.U28.ZN ) ,
    .I0 ( config0_decoder12.U28.AB ) ,
    .I1 ( config0_decoder12.n52 ) ) ;
not ( 
    .O1 ( config0_decoder12.n1 ) ,
    .IN ( config0_decoder12.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U77.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n47 ) ) ;
and ( 
    .Z ( config0_decoder12.U77.ZN ) ,
    .I0 ( config0_decoder12.U77.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_11 ) ,
    .IN ( config0_decoder12.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U67.AB ) ,
    .I0 ( config0_decoder12.n60 ) ,
    .I1 ( config0_decoder12.n59 ) ) ;
and ( 
    .Z ( config0_decoder12.U67.ZN ) ,
    .I0 ( config0_decoder12.U67.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_8 ) ,
    .IN ( config0_decoder12.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U10.AB ) ,
    .I0 ( config0_decoder12.n53 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U10.ZN ) ,
    .I0 ( config0_decoder12.U10.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_31 ) ,
    .IN ( config0_decoder12.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n50 ) ,
    .I0 ( config0_decoder12.n40 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
or ( 
    .Z ( config0_decoder12.U26.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n54 ) ) ;
and ( 
    .Z ( config0_decoder12.U26.ZN ) ,
    .I0 ( config0_decoder12.U26.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_2 ) ,
    .IN ( config0_decoder12.U26.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n62 ) ,
    .I0 ( config0_decoder12.n35 ) ,
    .I1 ( config0_decoder12.n51 ) ) ;
or ( 
    .Z ( config0_decoder12.U86.AB ) ,
    .I0 ( config0_decoder12.n57 ) ,
    .I1 ( config0_decoder12.n56 ) ) ;
and ( 
    .Z ( config0_decoder12.U86.ZN ) ,
    .I0 ( config0_decoder12.U86.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_52 ) ,
    .IN ( config0_decoder12.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U58.AB ) ,
    .I0 ( config0_decoder12.n56 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U58.ZN ) ,
    .I0 ( config0_decoder12.U58.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_36 ) ,
    .IN ( config0_decoder12.U58.ZN ) ) ;
not ( 
    .O1 ( config0_decoder12.n36 ) ,
    .IN ( masks_hold_reg_10_8 ) ) ;
or ( 
    .Z ( config0_decoder12.U74.AB ) ,
    .I0 ( config0_decoder12.n54 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U74.ZN ) ,
    .I0 ( config0_decoder12.U74.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_17 ) ,
    .IN ( config0_decoder12.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U66.AB ) ,
    .I0 ( config0_decoder12.n58 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U66.ZN ) ,
    .I0 ( config0_decoder12.U66.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_22 ) ,
    .IN ( config0_decoder12.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U11.AB ) ,
    .I0 ( config0_decoder12.n57 ) ,
    .I1 ( config0_decoder12.n53 ) ) ;
and ( 
    .Z ( config0_decoder12.U11.ZN ) ,
    .I0 ( config0_decoder12.U11.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_48 ) ,
    .IN ( config0_decoder12.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder12.n37 ) ,
    .I0 ( config0_decoder12.n36 ) ,
    .I1 ( masks_hold_reg_10_9 ) ) ;
nand ( 
    .Z ( config0_decoder12.n44 ) ,
    .I0 ( config0_decoder12.n37 ) ,
    .I1 ( masks_hold_reg_10_4 ) ) ;
nand ( 
    .Z ( config0_decoder12.n43 ) ,
    .I0 ( config0_decoder12.n37 ) ,
    .I1 ( config0_decoder12.n51 ) ) ;
or ( 
    .Z ( config0_decoder12.U81.AB ) ,
    .I0 ( config0_decoder12.n60 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U81.ZN ) ,
    .I0 ( config0_decoder12.U81.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_39 ) ,
    .IN ( config0_decoder12.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U59.AB ) ,
    .I0 ( config0_decoder12.n56 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U59.ZN ) ,
    .I0 ( config0_decoder12.U59.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_20 ) ,
    .IN ( config0_decoder12.U59.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U49.AB ) ,
    .I0 ( config0_decoder12.n55 ) ,
    .I1 ( config0_decoder12.n53 ) ) ;
and ( 
    .Z ( config0_decoder12.U49.ZN ) ,
    .I0 ( config0_decoder12.U49.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_47 ) ,
    .IN ( config0_decoder12.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U75.AB ) ,
    .I0 ( config0_decoder12.n58 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U75.ZN ) ,
    .I0 ( config0_decoder12.U75.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_21 ) ,
    .IN ( config0_decoder12.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U65.AB ) ,
    .I0 ( config0_decoder12.n58 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U65.ZN ) ,
    .I0 ( config0_decoder12.U65.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_38 ) ,
    .IN ( config0_decoder12.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U12.AB ) ,
    .I0 ( config0_decoder12.n47 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U12.ZN ) ,
    .I0 ( config0_decoder12.U12.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_28 ) ,
    .IN ( config0_decoder12.U12.ZN ) ) ;
not ( 
    .O1 ( config0_decoder12.n45 ) ,
    .IN ( masks_hold_reg_10_9 ) ) ;
nand ( 
    .Z ( config0_decoder12.n54 ) ,
    .I0 ( config0_decoder12.n38 ) ,
    .I1 ( masks_hold_reg_10_5 ) ) ;
nand ( 
    .Z ( config0_decoder12.n56 ) ,
    .I0 ( config0_decoder12.n41 ) ,
    .I1 ( config0_decoder12.n39 ) ,
    .I2 ( masks_hold_reg_10_6 ) ) ;
or ( 
    .Z ( config0_decoder12.U80.AB ) ,
    .I0 ( config0_decoder12.n56 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U80.ZN ) ,
    .I0 ( config0_decoder12.U80.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_35 ) ,
    .IN ( config0_decoder12.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U48.AB ) ,
    .I0 ( config0_decoder12.n53 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U48.ZN ) ,
    .I0 ( config0_decoder12.U48.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_32 ) ,
    .IN ( config0_decoder12.U48.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U64.AB ) ,
    .I0 ( config0_decoder12.n54 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U64.ZN ) ,
    .I0 ( config0_decoder12.U64.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_34 ) ,
    .IN ( config0_decoder12.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U13.AB ) ,
    .I0 ( config0_decoder12.n50 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U13.ZN ) ,
    .I0 ( config0_decoder12.U13.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_30 ) ,
    .IN ( config0_decoder12.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n49 ) ,
    .I0 ( config0_decoder12.n46 ) ,
    .I1 ( masks_hold_reg_10_4 ) ) ;
or ( 
    .Z ( config0_decoder12.U83.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n62 ) ) ;
and ( 
    .Z ( config0_decoder12.U83.ZN ) ,
    .I0 ( config0_decoder12.U83.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_9 ) ,
    .IN ( config0_decoder12.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U50.AB ) ,
    .I0 ( config0_decoder12.n49 ) ,
    .I1 ( config0_decoder12.n47 ) ) ;
and ( 
    .Z ( config0_decoder12.U50.ZN ) ,
    .I0 ( config0_decoder12.U50.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_44 ) ,
    .IN ( config0_decoder12.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n47 ) ,
    .I0 ( masks_hold_reg_10_7 ) ,
    .I1 ( config0_decoder12.n41 ) ,
    .I2 ( masks_hold_reg_10_6 ) ) ;
or ( 
    .Z ( config0_decoder12.U82.AB ) ,
    .I0 ( config0_decoder12.n60 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U82.ZN ) ,
    .I0 ( config0_decoder12.U82.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_23 ) ,
    .IN ( config0_decoder12.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U51.AB ) ,
    .I0 ( config0_decoder12.n56 ) ,
    .I1 ( config0_decoder12.n55 ) ) ;
and ( 
    .Z ( config0_decoder12.U51.ZN ) ,
    .I0 ( config0_decoder12.U51.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_51 ) ,
    .IN ( config0_decoder12.U51.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n57 ) ,
    .I0 ( masks_hold_reg_10_4 ) ,
    .I1 ( config0_decoder12.n52 ) ) ;
or ( 
    .Z ( config0_decoder12.U78.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U78.ZN ) ,
    .I0 ( config0_decoder12.U78.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_41 ) ,
    .IN ( config0_decoder12.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n59 ) ,
    .I0 ( masks_hold_reg_10_4 ) ,
    .I1 ( config0_decoder12.n35 ) ) ;
or ( 
    .Z ( config0_decoder12.U21.AB ) ,
    .I0 ( config0_decoder12.n55 ) ,
    .I1 ( config0_decoder12.n54 ) ) ;
and ( 
    .Z ( config0_decoder12.U21.ZN ) ,
    .I0 ( config0_decoder12.U21.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_49 ) ,
    .IN ( config0_decoder12.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n60 ) ,
    .I0 ( config0_decoder12.n42 ) ,
    .I1 ( config0_decoder12.n41 ) ) ;
and ( 
    .Z ( config0_decoder12.n40 ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( masks_hold_reg_10_5 ) ) ;
nor ( 
    .Z ( config0_decoder12.n38 ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
or ( 
    .Z ( config0_decoder12.U79.AB ) ,
    .I0 ( config0_decoder12.n47 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U79.ZN ) ,
    .I0 ( config0_decoder12.U79.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_27 ) ,
    .IN ( config0_decoder12.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U72.AB ) ,
    .I0 ( config0_decoder12.n54 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U72.ZN ) ,
    .I0 ( config0_decoder12.U72.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_33 ) ,
    .IN ( config0_decoder12.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U69.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U69.ZN ) ,
    .I0 ( config0_decoder12.U69.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_42 ) ,
    .IN ( config0_decoder12.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U20.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n56 ) ) ;
and ( 
    .Z ( config0_decoder12.U20.ZN ) ,
    .I0 ( config0_decoder12.U20.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_3 ) ,
    .IN ( config0_decoder12.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U9.AB ) ,
    .I0 ( config0_decoder12.n53 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U9.ZN ) ,
    .I0 ( config0_decoder12.U9.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_16 ) ,
    .IN ( config0_decoder12.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n53 ) ,
    .I0 ( config0_decoder12.n38 ) ,
    .I1 ( config0_decoder12.n41 ) ) ;
or ( 
    .Z ( config0_decoder12.U53.AB ) ,
    .I0 ( config0_decoder12.n50 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U53.ZN ) ,
    .I0 ( config0_decoder12.U53.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_46 ) ,
    .IN ( config0_decoder12.U53.ZN ) ) ;
nor ( 
    .Z ( config0_decoder12.n46 ) ,
    .I0 ( config0_decoder12.n45 ) ,
    .I1 ( masks_hold_reg_10_8 ) ) ;
or ( 
    .Z ( config0_decoder12.U73.AB ) ,
    .I0 ( config0_decoder12.n58 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U73.ZN ) ,
    .I0 ( config0_decoder12.U73.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_37 ) ,
    .IN ( config0_decoder12.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U68.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n47 ) ) ;
and ( 
    .Z ( config0_decoder12.U68.ZN ) ,
    .I0 ( config0_decoder12.U68.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_12 ) ,
    .IN ( config0_decoder12.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U63.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U63.ZN ) ,
    .I0 ( config0_decoder12.U63.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_26 ) ,
    .IN ( config0_decoder12.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U14.AB ) ,
    .I0 ( config0_decoder12.n54 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U14.ZN ) ,
    .I0 ( config0_decoder12.U14.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_18 ) ,
    .IN ( config0_decoder12.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n55 ) ,
    .I0 ( config0_decoder12.n52 ) ,
    .I1 ( config0_decoder12.n51 ) ) ;
nor ( 
    .Z ( config0_decoder12.n52 ) ,
    .I0 ( config0_decoder12.n45 ) ,
    .I1 ( config0_decoder12.n36 ) ) ;
or ( 
    .Z ( config0_decoder12.U54.AB ) ,
    .I0 ( config0_decoder12.n50 ) ,
    .I1 ( config0_decoder12.n48 ) ) ;
and ( 
    .Z ( config0_decoder12.U54.ZN ) ,
    .I0 ( config0_decoder12.U54.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_45 ) ,
    .IN ( config0_decoder12.U54.ZN ) ) ;
not ( 
    .O1 ( config0_decoder12.n39 ) ,
    .IN ( masks_hold_reg_10_7 ) ) ;
or ( 
    .Z ( config0_decoder12.U70.AB ) ,
    .I0 ( config0_decoder12.n50 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U70.ZN ) ,
    .I0 ( config0_decoder12.U70.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_29 ) ,
    .IN ( config0_decoder12.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U62.AB ) ,
    .I0 ( config0_decoder12.n60 ) ,
    .I1 ( config0_decoder12.n49 ) ) ;
and ( 
    .Z ( config0_decoder12.U62.ZN ) ,
    .I0 ( config0_decoder12.U62.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_40 ) ,
    .IN ( config0_decoder12.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U18.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n58 ) ) ;
and ( 
    .Z ( config0_decoder12.U18.ZN ) ,
    .I0 ( config0_decoder12.U18.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_6 ) ,
    .IN ( config0_decoder12.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U15.AB ) ,
    .I0 ( config0_decoder12.n56 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U15.ZN ) ,
    .I0 ( config0_decoder12.U15.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_19 ) ,
    .IN ( config0_decoder12.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n58 ) ,
    .I0 ( config0_decoder12.n40 ) ,
    .I1 ( config0_decoder12.n39 ) ) ;
or ( 
    .Z ( config0_decoder12.U85.AB ) ,
    .I0 ( config0_decoder12.n48 ) ,
    .I1 ( config0_decoder12.n47 ) ) ;
and ( 
    .Z ( config0_decoder12.U85.ZN ) ,
    .I0 ( config0_decoder12.U85.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_43 ) ,
    .IN ( config0_decoder12.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U55.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n58 ) ) ;
and ( 
    .Z ( config0_decoder12.U55.ZN ) ,
    .I0 ( config0_decoder12.U55.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_5 ) ,
    .IN ( config0_decoder12.U55.ZN ) ) ;
not ( 
    .O1 ( config0_decoder12.n51 ) ,
    .IN ( masks_hold_reg_10_4 ) ) ;
or ( 
    .Z ( config0_decoder12.U71.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U71.ZN ) ,
    .I0 ( config0_decoder12.U71.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_25 ) ,
    .IN ( config0_decoder12.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U61.AB ) ,
    .I0 ( config0_decoder12.n63 ) ,
    .I1 ( config0_decoder12.n59 ) ) ;
and ( 
    .Z ( config0_decoder12.U61.ZN ) ,
    .I0 ( config0_decoder12.U61.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_10 ) ,
    .IN ( config0_decoder12.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U19.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n53 ) ) ;
and ( 
    .Z ( config0_decoder12.U19.ZN ) ,
    .I0 ( config0_decoder12.U19.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_0 ) ,
    .IN ( config0_decoder12.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U16.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n56 ) ) ;
and ( 
    .Z ( config0_decoder12.U16.ZN ) ,
    .I0 ( config0_decoder12.U16.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_4 ) ,
    .IN ( config0_decoder12.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder12.n63 ) ,
    .I0 ( masks_hold_reg_10_5 ) ,
    .I1 ( config0_decoder12.n42 ) ) ;
nand ( 
    .Z ( config0_decoder12.n48 ) ,
    .I0 ( config0_decoder12.n46 ) ,
    .I1 ( config0_decoder12.n51 ) ) ;
or ( 
    .Z ( config0_decoder12.U84.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n50 ) ) ;
and ( 
    .Z ( config0_decoder12.U84.ZN ) ,
    .I0 ( config0_decoder12.U84.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_13 ) ,
    .IN ( config0_decoder12.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U56.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n54 ) ) ;
and ( 
    .Z ( config0_decoder12.U56.ZN ) ,
    .I0 ( config0_decoder12.U56.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_1 ) ,
    .IN ( config0_decoder12.U56.ZN ) ) ;
nor ( 
    .Z ( config0_decoder12.n42 ) ,
    .I0 ( config0_decoder12.n39 ) ,
    .I1 ( masks_hold_reg_10_6 ) ) ;
or ( 
    .Z ( config0_decoder12.U76.AB ) ,
    .I0 ( config0_decoder12.n53 ) ,
    .I1 ( config0_decoder12.n43 ) ) ;
and ( 
    .Z ( config0_decoder12.U76.ZN ) ,
    .I0 ( config0_decoder12.U76.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_15 ) ,
    .IN ( config0_decoder12.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U60.AB ) ,
    .I0 ( config0_decoder12.n59 ) ,
    .I1 ( config0_decoder12.n50 ) ) ;
and ( 
    .Z ( config0_decoder12.U60.ZN ) ,
    .I0 ( config0_decoder12.U60.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_14 ) ,
    .IN ( config0_decoder12.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U17.AB ) ,
    .I0 ( config0_decoder12.n62 ) ,
    .I1 ( config0_decoder12.n60 ) ) ;
and ( 
    .Z ( config0_decoder12.U17.ZN ) ,
    .I0 ( config0_decoder12.U17.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_7 ) ,
    .IN ( config0_decoder12.U17.ZN ) ) ;
nor ( 
    .Z ( config0_decoder12.n35 ) ,
    .I0 ( masks_hold_reg_10_8 ) ,
    .I1 ( masks_hold_reg_10_9 ) ) ;
or ( 
    .Z ( config0_decoder12.U87.AB ) ,
    .I0 ( config0_decoder12.n57 ) ,
    .I1 ( config0_decoder12.n54 ) ) ;
and ( 
    .Z ( config0_decoder12.U87.ZN ) ,
    .I0 ( config0_decoder12.U87.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_50 ) ,
    .IN ( config0_decoder12.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder12.U57.AB ) ,
    .I0 ( config0_decoder12.n60 ) ,
    .I1 ( config0_decoder12.n44 ) ) ;
and ( 
    .Z ( config0_decoder12.U57.ZN ) ,
    .I0 ( config0_decoder12.U57.AB ) ,
    .I1 ( config0_decoder12.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_11_24 ) ,
    .IN ( config0_decoder12.U57.ZN ) ) ;
not ( 
    .O1 ( config0_decoder12.n41 ) ,
    .IN ( masks_hold_reg_10_5 ) ) ;
or ( 
    .Z ( config0_decoder13.U37.AB ) ,
    .I0 ( config0_decoder13.n40 ) ,
    .I1 ( masks_hold_reg_11_8 ) ) ;
and ( 
    .Z ( config0_decoder13.U37.ZN ) ,
    .I0 ( config0_decoder13.U37.AB ) ,
    .I1 ( config0_decoder13.n52 ) ) ;
not ( 
    .O1 ( config0_decoder13.n1 ) ,
    .IN ( config0_decoder13.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U62.AB ) ,
    .I0 ( config0_decoder13.n50 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U62.ZN ) ,
    .I0 ( config0_decoder13.U62.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_46 ) ,
    .IN ( config0_decoder13.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U18.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n54 ) ) ;
and ( 
    .Z ( config0_decoder13.U18.ZN ) ,
    .I0 ( config0_decoder13.U18.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_2 ) ,
    .IN ( config0_decoder13.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U15.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n58 ) ) ;
and ( 
    .Z ( config0_decoder13.U15.ZN ) ,
    .I0 ( config0_decoder13.U15.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_6 ) ,
    .IN ( config0_decoder13.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n53 ) ,
    .I0 ( config0_decoder13.n38 ) ,
    .I1 ( config0_decoder13.n41 ) ) ;
or ( 
    .Z ( config0_decoder13.U85.AB ) ,
    .I0 ( config0_decoder13.n48 ) ,
    .I1 ( config0_decoder13.n47 ) ) ;
and ( 
    .Z ( config0_decoder13.U85.ZN ) ,
    .I0 ( config0_decoder13.U85.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_43 ) ,
    .IN ( config0_decoder13.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U55.AB ) ,
    .I0 ( config0_decoder13.n55 ) ,
    .I1 ( config0_decoder13.n53 ) ) ;
and ( 
    .Z ( config0_decoder13.U55.ZN ) ,
    .I0 ( config0_decoder13.U55.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_47 ) ,
    .IN ( config0_decoder13.U55.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n63 ) ,
    .I0 ( masks_hold_reg_11_6 ) ,
    .I1 ( config0_decoder13.n42 ) ) ;
or ( 
    .Z ( config0_decoder13.U71.AB ) ,
    .I0 ( config0_decoder13.n60 ) ,
    .I1 ( config0_decoder13.n59 ) ) ;
and ( 
    .Z ( config0_decoder13.U71.ZN ) ,
    .I0 ( config0_decoder13.U71.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_8 ) ,
    .IN ( config0_decoder13.U71.ZN ) ) ;
and ( 
    .Z ( config0_decoder13.n40 ) ,
    .I0 ( masks_hold_reg_11_7 ) ,
    .I1 ( masks_hold_reg_11_6 ) ) ;
or ( 
    .Z ( config0_decoder13.U19.AB ) ,
    .I0 ( config0_decoder13.n55 ) ,
    .I1 ( config0_decoder13.n54 ) ) ;
and ( 
    .Z ( config0_decoder13.U19.ZN ) ,
    .I0 ( config0_decoder13.U19.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_49 ) ,
    .IN ( config0_decoder13.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U16.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n53 ) ) ;
and ( 
    .Z ( config0_decoder13.U16.ZN ) ,
    .I0 ( config0_decoder13.U16.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_0 ) ,
    .IN ( config0_decoder13.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U36.AB ) ,
    .I0 ( config0_decoder13.n56 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U36.ZN ) ,
    .I0 ( config0_decoder13.U36.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_35 ) ,
    .IN ( config0_decoder13.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U1.AB ) ,
    .I0 ( config0_decoder13.n53 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U1.ZN ) ,
    .I0 ( config0_decoder13.U1.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_31 ) ,
    .IN ( config0_decoder13.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U84.AB ) ,
    .I0 ( config0_decoder13.n56 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U84.ZN ) ,
    .I0 ( config0_decoder13.U84.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_19 ) ,
    .IN ( config0_decoder13.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U56.AB ) ,
    .I0 ( config0_decoder13.n49 ) ,
    .I1 ( config0_decoder13.n47 ) ) ;
and ( 
    .Z ( config0_decoder13.U56.ZN ) ,
    .I0 ( config0_decoder13.U56.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_44 ) ,
    .IN ( config0_decoder13.U56.ZN ) ) ;
nor ( 
    .Z ( config0_decoder13.n35 ) ,
    .I0 ( masks_hold_reg_11_9 ) ,
    .I1 ( masks_hold_reg_11_10 ) ) ;
or ( 
    .Z ( config0_decoder13.U76.AB ) ,
    .I0 ( config0_decoder13.n53 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U76.ZN ) ,
    .I0 ( config0_decoder13.U76.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_15 ) ,
    .IN ( config0_decoder13.U76.ZN ) ) ;
not ( 
    .O1 ( config0_decoder13.n45 ) ,
    .IN ( masks_hold_reg_11_10 ) ) ;
or ( 
    .Z ( config0_decoder13.U17.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n56 ) ) ;
and ( 
    .Z ( config0_decoder13.U17.ZN ) ,
    .I0 ( config0_decoder13.U17.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_3 ) ,
    .IN ( config0_decoder13.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U87.AB ) ,
    .I0 ( config0_decoder13.n57 ) ,
    .I1 ( config0_decoder13.n54 ) ) ;
and ( 
    .Z ( config0_decoder13.U87.ZN ) ,
    .I0 ( config0_decoder13.U87.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_50 ) ,
    .IN ( config0_decoder13.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U57.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n58 ) ) ;
and ( 
    .Z ( config0_decoder13.U57.ZN ) ,
    .I0 ( config0_decoder13.U57.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_5 ) ,
    .IN ( config0_decoder13.U57.ZN ) ) ;
nor ( 
    .Z ( config0_decoder13.n46 ) ,
    .I0 ( config0_decoder13.n45 ) ,
    .I1 ( masks_hold_reg_11_9 ) ) ;
or ( 
    .Z ( config0_decoder13.U77.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n47 ) ) ;
and ( 
    .Z ( config0_decoder13.U77.ZN ) ,
    .I0 ( config0_decoder13.U77.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_11 ) ,
    .IN ( config0_decoder13.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U67.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n59 ) ) ;
and ( 
    .Z ( config0_decoder13.U67.ZN ) ,
    .I0 ( config0_decoder13.U67.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_10 ) ,
    .IN ( config0_decoder13.U67.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n55 ) ,
    .I0 ( config0_decoder13.n52 ) ,
    .I1 ( config0_decoder13.n51 ) ) ;
or ( 
    .Z ( config0_decoder13.U34.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U34.ZN ) ,
    .I0 ( config0_decoder13.U34.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_25 ) ,
    .IN ( config0_decoder13.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U26.AB ) ,
    .I0 ( config0_decoder13.n57 ) ,
    .I1 ( config0_decoder13.n53 ) ) ;
and ( 
    .Z ( config0_decoder13.U26.ZN ) ,
    .I0 ( config0_decoder13.U26.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_48 ) ,
    .IN ( config0_decoder13.U26.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n48 ) ,
    .I0 ( config0_decoder13.n46 ) ,
    .I1 ( config0_decoder13.n51 ) ) ;
or ( 
    .Z ( config0_decoder13.U86.AB ) ,
    .I0 ( config0_decoder13.n57 ) ,
    .I1 ( config0_decoder13.n56 ) ) ;
and ( 
    .Z ( config0_decoder13.U86.ZN ) ,
    .I0 ( config0_decoder13.U86.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_52 ) ,
    .IN ( config0_decoder13.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U58.AB ) ,
    .I0 ( config0_decoder13.n56 ) ,
    .I1 ( config0_decoder13.n55 ) ) ;
and ( 
    .Z ( config0_decoder13.U58.ZN ) ,
    .I0 ( config0_decoder13.U58.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_51 ) ,
    .IN ( config0_decoder13.U58.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n50 ) ,
    .I0 ( config0_decoder13.n40 ) ,
    .I1 ( masks_hold_reg_11_8 ) ) ;
or ( 
    .Z ( config0_decoder13.U74.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U74.ZN ) ,
    .I0 ( config0_decoder13.U74.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_42 ) ,
    .IN ( config0_decoder13.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U66.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n50 ) ) ;
and ( 
    .Z ( config0_decoder13.U66.ZN ) ,
    .I0 ( config0_decoder13.U66.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_14 ) ,
    .IN ( config0_decoder13.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U11.AB ) ,
    .I0 ( config0_decoder13.n50 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U11.ZN ) ,
    .I0 ( config0_decoder13.U11.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_30 ) ,
    .IN ( config0_decoder13.U11.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n56 ) ,
    .I0 ( config0_decoder13.n41 ) ,
    .I1 ( config0_decoder13.n39 ) ,
    .I2 ( masks_hold_reg_11_7 ) ) ;
or ( 
    .Z ( config0_decoder13.U35.AB ) ,
    .I0 ( config0_decoder13.n58 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U35.ZN ) ,
    .I0 ( config0_decoder13.U35.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_37 ) ,
    .IN ( config0_decoder13.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U2.AB ) ,
    .I0 ( config0_decoder13.n47 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U2.ZN ) ,
    .I0 ( config0_decoder13.U2.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_28 ) ,
    .IN ( config0_decoder13.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U81.AB ) ,
    .I0 ( config0_decoder13.n60 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U81.ZN ) ,
    .I0 ( config0_decoder13.U81.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_39 ) ,
    .IN ( config0_decoder13.U81.ZN ) ) ;
not ( 
    .O1 ( config0_decoder13.n39 ) ,
    .IN ( masks_hold_reg_11_8 ) ) ;
nand ( 
    .Z ( config0_decoder13.n57 ) ,
    .I0 ( masks_hold_reg_11_5 ) ,
    .I1 ( config0_decoder13.n52 ) ) ;
or ( 
    .Z ( config0_decoder13.U75.AB ) ,
    .I0 ( config0_decoder13.n58 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U75.ZN ) ,
    .I0 ( config0_decoder13.U75.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_21 ) ,
    .IN ( config0_decoder13.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U65.AB ) ,
    .I0 ( config0_decoder13.n56 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U65.ZN ) ,
    .I0 ( config0_decoder13.U65.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_36 ) ,
    .IN ( config0_decoder13.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U12.AB ) ,
    .I0 ( config0_decoder13.n58 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U12.ZN ) ,
    .I0 ( config0_decoder13.U12.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_22 ) ,
    .IN ( config0_decoder13.U12.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n47 ) ,
    .I0 ( masks_hold_reg_11_8 ) ,
    .I1 ( config0_decoder13.n41 ) ,
    .I2 ( masks_hold_reg_11_7 ) ) ;
or ( 
    .Z ( config0_decoder13.U32.AB ) ,
    .I0 ( config0_decoder13.n50 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U32.ZN ) ,
    .I0 ( config0_decoder13.U32.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_29 ) ,
    .IN ( config0_decoder13.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U29.AB ) ,
    .I0 ( config0_decoder13.n60 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U29.ZN ) ,
    .I0 ( config0_decoder13.U29.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_24 ) ,
    .IN ( config0_decoder13.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U80.AB ) ,
    .I0 ( config0_decoder13.n47 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U80.ZN ) ,
    .I0 ( config0_decoder13.U80.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_27 ) ,
    .IN ( config0_decoder13.U80.ZN ) ) ;
not ( 
    .O1 ( config0_decoder13.n36 ) ,
    .IN ( masks_hold_reg_11_9 ) ) ;
or ( 
    .Z ( config0_decoder13.U64.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n54 ) ) ;
and ( 
    .Z ( config0_decoder13.U64.ZN ) ,
    .I0 ( config0_decoder13.U64.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_1 ) ,
    .IN ( config0_decoder13.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U13.AB ) ,
    .I0 ( config0_decoder13.n60 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U13.ZN ) ,
    .I0 ( config0_decoder13.U13.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_23 ) ,
    .IN ( config0_decoder13.U13.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U33.AB ) ,
    .I0 ( config0_decoder13.n54 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U33.ZN ) ,
    .I0 ( config0_decoder13.U33.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_33 ) ,
    .IN ( config0_decoder13.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U28.AB ) ,
    .I0 ( config0_decoder13.n53 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U28.ZN ) ,
    .I0 ( config0_decoder13.U28.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_32 ) ,
    .IN ( config0_decoder13.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U83.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n50 ) ) ;
and ( 
    .Z ( config0_decoder13.U83.ZN ) ,
    .I0 ( config0_decoder13.U83.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_13 ) ,
    .IN ( config0_decoder13.U83.ZN ) ) ;
nor ( 
    .Z ( config0_decoder13.n38 ) ,
    .I0 ( masks_hold_reg_11_7 ) ,
    .I1 ( masks_hold_reg_11_8 ) ) ;
or ( 
    .Z ( config0_decoder13.U30.AB ) ,
    .I0 ( config0_decoder13.n54 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U30.ZN ) ,
    .I0 ( config0_decoder13.U30.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_34 ) ,
    .IN ( config0_decoder13.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U82.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n62 ) ) ;
and ( 
    .Z ( config0_decoder13.U82.ZN ) ,
    .I0 ( config0_decoder13.U82.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_9 ) ,
    .IN ( config0_decoder13.U82.ZN ) ) ;
nor ( 
    .Z ( config0_decoder13.n37 ) ,
    .I0 ( config0_decoder13.n36 ) ,
    .I1 ( masks_hold_reg_11_10 ) ) ;
nand ( 
    .Z ( config0_decoder13.n54 ) ,
    .I0 ( config0_decoder13.n38 ) ,
    .I1 ( masks_hold_reg_11_6 ) ) ;
or ( 
    .Z ( config0_decoder13.U78.AB ) ,
    .I0 ( config0_decoder13.n54 ) ,
    .I1 ( config0_decoder13.n43 ) ) ;
and ( 
    .Z ( config0_decoder13.U78.ZN ) ,
    .I0 ( config0_decoder13.U78.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_17 ) ,
    .IN ( config0_decoder13.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U31.AB ) ,
    .I0 ( config0_decoder13.n58 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U31.ZN ) ,
    .I0 ( config0_decoder13.U31.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_38 ) ,
    .IN ( config0_decoder13.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U21.AB ) ,
    .I0 ( config0_decoder13.n62 ) ,
    .I1 ( config0_decoder13.n60 ) ) ;
and ( 
    .Z ( config0_decoder13.U21.ZN ) ,
    .I0 ( config0_decoder13.U21.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_7 ) ,
    .IN ( config0_decoder13.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n43 ) ,
    .I0 ( config0_decoder13.n37 ) ,
    .I1 ( config0_decoder13.n51 ) ) ;
not ( 
    .O1 ( config0_decoder13.n51 ) ,
    .IN ( masks_hold_reg_11_5 ) ) ;
nand ( 
    .Z ( config0_decoder13.n59 ) ,
    .I0 ( masks_hold_reg_11_5 ) ,
    .I1 ( config0_decoder13.n35 ) ) ;
or ( 
    .Z ( config0_decoder13.U79.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U79.ZN ) ,
    .I0 ( config0_decoder13.U79.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_41 ) ,
    .IN ( config0_decoder13.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U72.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n47 ) ) ;
and ( 
    .Z ( config0_decoder13.U72.ZN ) ,
    .I0 ( config0_decoder13.U72.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_12 ) ,
    .IN ( config0_decoder13.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U69.AB ) ,
    .I0 ( config0_decoder13.n60 ) ,
    .I1 ( config0_decoder13.n49 ) ) ;
and ( 
    .Z ( config0_decoder13.U69.ZN ) ,
    .I0 ( config0_decoder13.U69.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_40 ) ,
    .IN ( config0_decoder13.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U20.AB ) ,
    .I0 ( config0_decoder13.n56 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U20.ZN ) ,
    .I0 ( config0_decoder13.U20.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_20 ) ,
    .IN ( config0_decoder13.U20.ZN ) ) ;
nor ( 
    .Z ( config0_decoder13.n52 ) ,
    .I0 ( config0_decoder13.n45 ) ,
    .I1 ( config0_decoder13.n36 ) ) ;
nand ( 
    .Z ( config0_decoder13.n62 ) ,
    .I0 ( config0_decoder13.n35 ) ,
    .I1 ( config0_decoder13.n51 ) ) ;
nor ( 
    .Z ( config0_decoder13.n42 ) ,
    .I0 ( config0_decoder13.n39 ) ,
    .I1 ( masks_hold_reg_11_7 ) ) ;
nand ( 
    .Z ( config0_decoder13.n44 ) ,
    .I0 ( config0_decoder13.n37 ) ,
    .I1 ( masks_hold_reg_11_5 ) ) ;
or ( 
    .Z ( config0_decoder13.U73.AB ) ,
    .I0 ( config0_decoder13.n54 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U73.ZN ) ,
    .I0 ( config0_decoder13.U73.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_18 ) ,
    .IN ( config0_decoder13.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U68.AB ) ,
    .I0 ( config0_decoder13.n53 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U68.ZN ) ,
    .I0 ( config0_decoder13.U68.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_16 ) ,
    .IN ( config0_decoder13.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U63.AB ) ,
    .I0 ( config0_decoder13.n50 ) ,
    .I1 ( config0_decoder13.n48 ) ) ;
and ( 
    .Z ( config0_decoder13.U63.ZN ) ,
    .I0 ( config0_decoder13.U63.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_45 ) ,
    .IN ( config0_decoder13.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder13.U14.AB ) ,
    .I0 ( config0_decoder13.n59 ) ,
    .I1 ( config0_decoder13.n56 ) ) ;
and ( 
    .Z ( config0_decoder13.U14.ZN ) ,
    .I0 ( config0_decoder13.U14.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_4 ) ,
    .IN ( config0_decoder13.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder13.n58 ) ,
    .I0 ( config0_decoder13.n40 ) ,
    .I1 ( config0_decoder13.n39 ) ) ;
nand ( 
    .Z ( config0_decoder13.n60 ) ,
    .I0 ( config0_decoder13.n42 ) ,
    .I1 ( config0_decoder13.n41 ) ) ;
not ( 
    .O1 ( config0_decoder13.n41 ) ,
    .IN ( masks_hold_reg_11_6 ) ) ;
nand ( 
    .Z ( config0_decoder13.n49 ) ,
    .I0 ( config0_decoder13.n46 ) ,
    .I1 ( masks_hold_reg_11_5 ) ) ;
or ( 
    .Z ( config0_decoder13.U70.AB ) ,
    .I0 ( config0_decoder13.n63 ) ,
    .I1 ( config0_decoder13.n44 ) ) ;
and ( 
    .Z ( config0_decoder13.U70.ZN ) ,
    .I0 ( config0_decoder13.U70.AB ) ,
    .I1 ( config0_decoder13.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_12_26 ) ,
    .IN ( config0_decoder13.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U28.AB ) ,
    .I0 ( config0_decoder10.n40 ) ,
    .I1 ( masks_hold_reg_8_5 ) ) ;
and ( 
    .Z ( config0_decoder10.U28.ZN ) ,
    .I0 ( config0_decoder10.U28.AB ) ,
    .I1 ( config0_decoder10.n52 ) ) ;
not ( 
    .O1 ( config0_decoder10.n1 ) ,
    .IN ( config0_decoder10.U28.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n55 ) ,
    .I0 ( config0_decoder10.n52 ) ,
    .I1 ( config0_decoder10.n51 ) ) ;
nor ( 
    .Z ( config0_decoder10.n52 ) ,
    .I0 ( config0_decoder10.n45 ) ,
    .I1 ( config0_decoder10.n36 ) ) ;
or ( 
    .Z ( config0_decoder10.U54.AB ) ,
    .I0 ( config0_decoder10.n49 ) ,
    .I1 ( config0_decoder10.n47 ) ) ;
and ( 
    .Z ( config0_decoder10.U54.ZN ) ,
    .I0 ( config0_decoder10.U54.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_44 ) ,
    .IN ( config0_decoder10.U54.ZN ) ) ;
nor ( 
    .Z ( config0_decoder10.n46 ) ,
    .I0 ( config0_decoder10.n45 ) ,
    .I1 ( masks_hold_reg_8_6 ) ) ;
or ( 
    .Z ( config0_decoder10.U70.AB ) ,
    .I0 ( config0_decoder10.n50 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U70.ZN ) ,
    .I0 ( config0_decoder10.U70.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_29 ) ,
    .IN ( config0_decoder10.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U62.AB ) ,
    .I0 ( config0_decoder10.n60 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U62.ZN ) ,
    .I0 ( config0_decoder10.U62.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_40 ) ,
    .IN ( config0_decoder10.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U18.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n53 ) ) ;
and ( 
    .Z ( config0_decoder10.U18.ZN ) ,
    .I0 ( config0_decoder10.U18.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_0 ) ,
    .IN ( config0_decoder10.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U15.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n56 ) ) ;
and ( 
    .Z ( config0_decoder10.U15.ZN ) ,
    .I0 ( config0_decoder10.U15.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_4 ) ,
    .IN ( config0_decoder10.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n58 ) ,
    .I0 ( config0_decoder10.n40 ) ,
    .I1 ( config0_decoder10.n39 ) ) ;
or ( 
    .Z ( config0_decoder10.U85.AB ) ,
    .I0 ( config0_decoder10.n56 ) ,
    .I1 ( config0_decoder10.n55 ) ) ;
and ( 
    .Z ( config0_decoder10.U85.ZN ) ,
    .I0 ( config0_decoder10.U85.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_51 ) ,
    .IN ( config0_decoder10.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U55.AB ) ,
    .I0 ( config0_decoder10.n50 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U55.ZN ) ,
    .I0 ( config0_decoder10.U55.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_45 ) ,
    .IN ( config0_decoder10.U55.ZN ) ) ;
nor ( 
    .Z ( config0_decoder10.n42 ) ,
    .I0 ( config0_decoder10.n39 ) ,
    .I1 ( masks_hold_reg_8_4 ) ) ;
or ( 
    .Z ( config0_decoder10.U71.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U71.ZN ) ,
    .I0 ( config0_decoder10.U71.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_25 ) ,
    .IN ( config0_decoder10.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U61.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n59 ) ) ;
and ( 
    .Z ( config0_decoder10.U61.ZN ) ,
    .I0 ( config0_decoder10.U61.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_10 ) ,
    .IN ( config0_decoder10.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U19.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n56 ) ) ;
and ( 
    .Z ( config0_decoder10.U19.ZN ) ,
    .I0 ( config0_decoder10.U19.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_3 ) ,
    .IN ( config0_decoder10.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U16.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n60 ) ) ;
and ( 
    .Z ( config0_decoder10.U16.ZN ) ,
    .I0 ( config0_decoder10.U16.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_7 ) ,
    .IN ( config0_decoder10.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n63 ) ,
    .I0 ( masks_hold_reg_8_3 ) ,
    .I1 ( config0_decoder10.n42 ) ) ;
nand ( 
    .Z ( config0_decoder10.n48 ) ,
    .I0 ( config0_decoder10.n46 ) ,
    .I1 ( config0_decoder10.n51 ) ) ;
or ( 
    .Z ( config0_decoder10.U84.AB ) ,
    .I0 ( config0_decoder10.n48 ) ,
    .I1 ( config0_decoder10.n47 ) ) ;
and ( 
    .Z ( config0_decoder10.U84.ZN ) ,
    .I0 ( config0_decoder10.U84.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_43 ) ,
    .IN ( config0_decoder10.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U56.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n54 ) ) ;
and ( 
    .Z ( config0_decoder10.U56.ZN ) ,
    .I0 ( config0_decoder10.U56.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_1 ) ,
    .IN ( config0_decoder10.U56.ZN ) ) ;
not ( 
    .O1 ( config0_decoder10.n45 ) ,
    .IN ( masks_hold_reg_8_7 ) ) ;
or ( 
    .Z ( config0_decoder10.U76.AB ) ,
    .I0 ( config0_decoder10.n53 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U76.ZN ) ,
    .I0 ( config0_decoder10.U76.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_15 ) ,
    .IN ( config0_decoder10.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U60.AB ) ,
    .I0 ( config0_decoder10.n56 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U60.ZN ) ,
    .I0 ( config0_decoder10.U60.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_20 ) ,
    .IN ( config0_decoder10.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U17.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n58 ) ) ;
and ( 
    .Z ( config0_decoder10.U17.ZN ) ,
    .I0 ( config0_decoder10.U17.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_6 ) ,
    .IN ( config0_decoder10.U17.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n57 ) ,
    .I0 ( masks_hold_reg_8_2 ) ,
    .I1 ( config0_decoder10.n52 ) ) ;
or ( 
    .Z ( config0_decoder10.U87.AB ) ,
    .I0 ( config0_decoder10.n57 ) ,
    .I1 ( config0_decoder10.n54 ) ) ;
and ( 
    .Z ( config0_decoder10.U87.ZN ) ,
    .I0 ( config0_decoder10.U87.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_50 ) ,
    .IN ( config0_decoder10.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U57.AB ) ,
    .I0 ( config0_decoder10.n60 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U57.ZN ) ,
    .I0 ( config0_decoder10.U57.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_24 ) ,
    .IN ( config0_decoder10.U57.ZN ) ) ;
not ( 
    .O1 ( config0_decoder10.n36 ) ,
    .IN ( masks_hold_reg_8_6 ) ) ;
or ( 
    .Z ( config0_decoder10.U77.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U77.ZN ) ,
    .I0 ( config0_decoder10.U77.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_41 ) ,
    .IN ( config0_decoder10.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U67.AB ) ,
    .I0 ( config0_decoder10.n60 ) ,
    .I1 ( config0_decoder10.n59 ) ) ;
and ( 
    .Z ( config0_decoder10.U67.ZN ) ,
    .I0 ( config0_decoder10.U67.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_8 ) ,
    .IN ( config0_decoder10.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U10.AB ) ,
    .I0 ( config0_decoder10.n50 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U10.ZN ) ,
    .I0 ( config0_decoder10.U10.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_30 ) ,
    .IN ( config0_decoder10.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n44 ) ,
    .I0 ( config0_decoder10.n37 ) ,
    .I1 ( masks_hold_reg_8_2 ) ) ;
nand ( 
    .Z ( config0_decoder10.n43 ) ,
    .I0 ( config0_decoder10.n37 ) ,
    .I1 ( config0_decoder10.n51 ) ) ;
or ( 
    .Z ( config0_decoder10.U86.AB ) ,
    .I0 ( config0_decoder10.n57 ) ,
    .I1 ( config0_decoder10.n56 ) ) ;
and ( 
    .Z ( config0_decoder10.U86.ZN ) ,
    .I0 ( config0_decoder10.U86.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_52 ) ,
    .IN ( config0_decoder10.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U58.AB ) ,
    .I0 ( config0_decoder10.n53 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U58.ZN ) ,
    .I0 ( config0_decoder10.U58.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_32 ) ,
    .IN ( config0_decoder10.U58.ZN ) ) ;
not ( 
    .O1 ( config0_decoder10.n41 ) ,
    .IN ( masks_hold_reg_8_3 ) ) ;
or ( 
    .Z ( config0_decoder10.U74.AB ) ,
    .I0 ( config0_decoder10.n54 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U74.ZN ) ,
    .I0 ( config0_decoder10.U74.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_17 ) ,
    .IN ( config0_decoder10.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U66.AB ) ,
    .I0 ( config0_decoder10.n58 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U66.ZN ) ,
    .I0 ( config0_decoder10.U66.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_22 ) ,
    .IN ( config0_decoder10.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U11.AB ) ,
    .I0 ( config0_decoder10.n53 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U11.ZN ) ,
    .I0 ( config0_decoder10.U11.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_31 ) ,
    .IN ( config0_decoder10.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder10.n35 ) ,
    .I0 ( masks_hold_reg_8_6 ) ,
    .I1 ( masks_hold_reg_8_7 ) ) ;
nand ( 
    .Z ( config0_decoder10.n50 ) ,
    .I0 ( config0_decoder10.n40 ) ,
    .I1 ( masks_hold_reg_8_5 ) ) ;
nand ( 
    .Z ( config0_decoder10.n62 ) ,
    .I0 ( config0_decoder10.n35 ) ,
    .I1 ( config0_decoder10.n51 ) ) ;
or ( 
    .Z ( config0_decoder10.U81.AB ) ,
    .I0 ( config0_decoder10.n60 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U81.ZN ) ,
    .I0 ( config0_decoder10.U81.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_23 ) ,
    .IN ( config0_decoder10.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U59.AB ) ,
    .I0 ( config0_decoder10.n56 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U59.ZN ) ,
    .I0 ( config0_decoder10.U59.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_36 ) ,
    .IN ( config0_decoder10.U59.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U49.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n47 ) ) ;
and ( 
    .Z ( config0_decoder10.U49.ZN ) ,
    .I0 ( config0_decoder10.U49.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_11 ) ,
    .IN ( config0_decoder10.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U75.AB ) ,
    .I0 ( config0_decoder10.n58 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U75.ZN ) ,
    .I0 ( config0_decoder10.U75.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_21 ) ,
    .IN ( config0_decoder10.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U65.AB ) ,
    .I0 ( config0_decoder10.n58 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U65.ZN ) ,
    .I0 ( config0_decoder10.U65.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_38 ) ,
    .IN ( config0_decoder10.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U12.AB ) ,
    .I0 ( config0_decoder10.n53 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U12.ZN ) ,
    .I0 ( config0_decoder10.U12.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_16 ) ,
    .IN ( config0_decoder10.U12.ZN ) ) ;
nor ( 
    .Z ( config0_decoder10.n37 ) ,
    .I0 ( config0_decoder10.n36 ) ,
    .I1 ( masks_hold_reg_8_7 ) ) ;
nand ( 
    .Z ( config0_decoder10.n49 ) ,
    .I0 ( config0_decoder10.n46 ) ,
    .I1 ( masks_hold_reg_8_2 ) ) ;
nand ( 
    .Z ( config0_decoder10.n56 ) ,
    .I0 ( config0_decoder10.n41 ) ,
    .I1 ( config0_decoder10.n39 ) ,
    .I2 ( masks_hold_reg_8_4 ) ) ;
or ( 
    .Z ( config0_decoder10.U80.AB ) ,
    .I0 ( config0_decoder10.n60 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U80.ZN ) ,
    .I0 ( config0_decoder10.U80.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_39 ) ,
    .IN ( config0_decoder10.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U48.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n50 ) ) ;
and ( 
    .Z ( config0_decoder10.U48.ZN ) ,
    .I0 ( config0_decoder10.U48.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_14 ) ,
    .IN ( config0_decoder10.U48.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U64.AB ) ,
    .I0 ( config0_decoder10.n54 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U64.ZN ) ,
    .I0 ( config0_decoder10.U64.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_34 ) ,
    .IN ( config0_decoder10.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U13.AB ) ,
    .I0 ( config0_decoder10.n54 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U13.ZN ) ,
    .I0 ( config0_decoder10.U13.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_18 ) ,
    .IN ( config0_decoder10.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n54 ) ,
    .I0 ( config0_decoder10.n38 ) ,
    .I1 ( masks_hold_reg_8_3 ) ) ;
or ( 
    .Z ( config0_decoder10.U83.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n50 ) ) ;
and ( 
    .Z ( config0_decoder10.U83.ZN ) ,
    .I0 ( config0_decoder10.U83.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_13 ) ,
    .IN ( config0_decoder10.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U50.AB ) ,
    .I0 ( config0_decoder10.n55 ) ,
    .I1 ( config0_decoder10.n53 ) ) ;
and ( 
    .Z ( config0_decoder10.U50.ZN ) ,
    .I0 ( config0_decoder10.U50.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_47 ) ,
    .IN ( config0_decoder10.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n47 ) ,
    .I0 ( masks_hold_reg_8_5 ) ,
    .I1 ( config0_decoder10.n41 ) ,
    .I2 ( masks_hold_reg_8_4 ) ) ;
or ( 
    .Z ( config0_decoder10.U22.AB ) ,
    .I0 ( config0_decoder10.n55 ) ,
    .I1 ( config0_decoder10.n54 ) ) ;
and ( 
    .Z ( config0_decoder10.U22.ZN ) ,
    .I0 ( config0_decoder10.U22.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_49 ) ,
    .IN ( config0_decoder10.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U82.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n62 ) ) ;
and ( 
    .Z ( config0_decoder10.U82.ZN ) ,
    .I0 ( config0_decoder10.U82.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_9 ) ,
    .IN ( config0_decoder10.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U51.AB ) ,
    .I0 ( config0_decoder10.n62 ) ,
    .I1 ( config0_decoder10.n58 ) ) ;
and ( 
    .Z ( config0_decoder10.U51.ZN ) ,
    .I0 ( config0_decoder10.U51.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_5 ) ,
    .IN ( config0_decoder10.U51.ZN ) ) ;
not ( 
    .O1 ( config0_decoder10.n39 ) ,
    .IN ( masks_hold_reg_8_5 ) ) ;
or ( 
    .Z ( config0_decoder10.U78.AB ) ,
    .I0 ( config0_decoder10.n47 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U78.ZN ) ,
    .I0 ( config0_decoder10.U78.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_27 ) ,
    .IN ( config0_decoder10.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n59 ) ,
    .I0 ( masks_hold_reg_8_2 ) ,
    .I1 ( config0_decoder10.n35 ) ) ;
or ( 
    .Z ( config0_decoder10.U21.AB ) ,
    .I0 ( config0_decoder10.n57 ) ,
    .I1 ( config0_decoder10.n53 ) ) ;
and ( 
    .Z ( config0_decoder10.U21.ZN ) ,
    .I0 ( config0_decoder10.U21.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_48 ) ,
    .IN ( config0_decoder10.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n60 ) ,
    .I0 ( config0_decoder10.n42 ) ,
    .I1 ( config0_decoder10.n41 ) ) ;
and ( 
    .Z ( config0_decoder10.n40 ) ,
    .I0 ( masks_hold_reg_8_4 ) ,
    .I1 ( masks_hold_reg_8_3 ) ) ;
nor ( 
    .Z ( config0_decoder10.n38 ) ,
    .I0 ( masks_hold_reg_8_4 ) ,
    .I1 ( masks_hold_reg_8_5 ) ) ;
or ( 
    .Z ( config0_decoder10.U79.AB ) ,
    .I0 ( config0_decoder10.n56 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U79.ZN ) ,
    .I0 ( config0_decoder10.U79.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_35 ) ,
    .IN ( config0_decoder10.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U72.AB ) ,
    .I0 ( config0_decoder10.n54 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U72.ZN ) ,
    .I0 ( config0_decoder10.U72.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_33 ) ,
    .IN ( config0_decoder10.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U69.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U69.ZN ) ,
    .I0 ( config0_decoder10.U69.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_42 ) ,
    .IN ( config0_decoder10.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U20.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n54 ) ) ;
and ( 
    .Z ( config0_decoder10.U20.ZN ) ,
    .I0 ( config0_decoder10.U20.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_2 ) ,
    .IN ( config0_decoder10.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U9.AB ) ,
    .I0 ( config0_decoder10.n47 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U9.ZN ) ,
    .I0 ( config0_decoder10.U9.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_28 ) ,
    .IN ( config0_decoder10.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder10.n53 ) ,
    .I0 ( config0_decoder10.n38 ) ,
    .I1 ( config0_decoder10.n41 ) ) ;
or ( 
    .Z ( config0_decoder10.U53.AB ) ,
    .I0 ( config0_decoder10.n50 ) ,
    .I1 ( config0_decoder10.n49 ) ) ;
and ( 
    .Z ( config0_decoder10.U53.ZN ) ,
    .I0 ( config0_decoder10.U53.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_46 ) ,
    .IN ( config0_decoder10.U53.ZN ) ) ;
not ( 
    .O1 ( config0_decoder10.n51 ) ,
    .IN ( masks_hold_reg_8_2 ) ) ;
or ( 
    .Z ( config0_decoder10.U73.AB ) ,
    .I0 ( config0_decoder10.n58 ) ,
    .I1 ( config0_decoder10.n48 ) ) ;
and ( 
    .Z ( config0_decoder10.U73.ZN ) ,
    .I0 ( config0_decoder10.U73.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_37 ) ,
    .IN ( config0_decoder10.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U68.AB ) ,
    .I0 ( config0_decoder10.n59 ) ,
    .I1 ( config0_decoder10.n47 ) ) ;
and ( 
    .Z ( config0_decoder10.U68.ZN ) ,
    .I0 ( config0_decoder10.U68.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_12 ) ,
    .IN ( config0_decoder10.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U63.AB ) ,
    .I0 ( config0_decoder10.n63 ) ,
    .I1 ( config0_decoder10.n44 ) ) ;
and ( 
    .Z ( config0_decoder10.U63.ZN ) ,
    .I0 ( config0_decoder10.U63.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_26 ) ,
    .IN ( config0_decoder10.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder10.U14.AB ) ,
    .I0 ( config0_decoder10.n56 ) ,
    .I1 ( config0_decoder10.n43 ) ) ;
and ( 
    .Z ( config0_decoder10.U14.ZN ) ,
    .I0 ( config0_decoder10.U14.AB ) ,
    .I1 ( config0_decoder10.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_9_19 ) ,
    .IN ( config0_decoder10.U14.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U38.AB ) ,
    .I0 ( config0_decoder11.n40 ) ,
    .I1 ( masks_hold_reg_9_6 ) ) ;
and ( 
    .Z ( config0_decoder11.U38.ZN ) ,
    .I0 ( config0_decoder11.U38.AB ) ,
    .I1 ( config0_decoder11.n52 ) ) ;
not ( 
    .O1 ( config0_decoder11.n1 ) ,
    .IN ( config0_decoder11.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U68.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n59 ) ) ;
and ( 
    .Z ( config0_decoder11.U68.ZN ) ,
    .I0 ( config0_decoder11.U68.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_10 ) ,
    .IN ( config0_decoder11.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U63.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n58 ) ) ;
and ( 
    .Z ( config0_decoder11.U63.ZN ) ,
    .I0 ( config0_decoder11.U63.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_5 ) ,
    .IN ( config0_decoder11.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U14.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n56 ) ) ;
and ( 
    .Z ( config0_decoder11.U14.ZN ) ,
    .I0 ( config0_decoder11.U14.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_4 ) ,
    .IN ( config0_decoder11.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n60 ) ,
    .I0 ( config0_decoder11.n42 ) ,
    .I1 ( config0_decoder11.n41 ) ) ;
nand ( 
    .Z ( config0_decoder11.n53 ) ,
    .I0 ( config0_decoder11.n38 ) ,
    .I1 ( config0_decoder11.n41 ) ) ;
nor ( 
    .Z ( config0_decoder11.n46 ) ,
    .I0 ( config0_decoder11.n45 ) ,
    .I1 ( masks_hold_reg_9_7 ) ) ;
nand ( 
    .Z ( config0_decoder11.n54 ) ,
    .I0 ( config0_decoder11.n38 ) ,
    .I1 ( masks_hold_reg_9_4 ) ) ;
or ( 
    .Z ( config0_decoder11.U70.AB ) ,
    .I0 ( config0_decoder11.n60 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U70.ZN ) ,
    .I0 ( config0_decoder11.U70.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_40 ) ,
    .IN ( config0_decoder11.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U62.AB ) ,
    .I0 ( config0_decoder11.n49 ) ,
    .I1 ( config0_decoder11.n47 ) ) ;
and ( 
    .Z ( config0_decoder11.U62.ZN ) ,
    .I0 ( config0_decoder11.U62.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_44 ) ,
    .IN ( config0_decoder11.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U18.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n56 ) ) ;
and ( 
    .Z ( config0_decoder11.U18.ZN ) ,
    .I0 ( config0_decoder11.U18.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_3 ) ,
    .IN ( config0_decoder11.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U15.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n60 ) ) ;
and ( 
    .Z ( config0_decoder11.U15.ZN ) ,
    .I0 ( config0_decoder11.U15.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_7 ) ,
    .IN ( config0_decoder11.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n62 ) ,
    .I0 ( config0_decoder11.n35 ) ,
    .I1 ( config0_decoder11.n51 ) ) ;
or ( 
    .Z ( config0_decoder11.U85.AB ) ,
    .I0 ( config0_decoder11.n56 ) ,
    .I1 ( config0_decoder11.n55 ) ) ;
and ( 
    .Z ( config0_decoder11.U85.ZN ) ,
    .I0 ( config0_decoder11.U85.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_51 ) ,
    .IN ( config0_decoder11.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U55.AB ) ,
    .I0 ( config0_decoder11.n58 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U55.ZN ) ,
    .I0 ( config0_decoder11.U55.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_21 ) ,
    .IN ( config0_decoder11.U55.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n63 ) ,
    .I0 ( masks_hold_reg_9_4 ) ,
    .I1 ( config0_decoder11.n42 ) ) ;
or ( 
    .Z ( config0_decoder11.U71.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U71.ZN ) ,
    .I0 ( config0_decoder11.U71.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_26 ) ,
    .IN ( config0_decoder11.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U61.AB ) ,
    .I0 ( config0_decoder11.n50 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U61.ZN ) ,
    .I0 ( config0_decoder11.U61.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_46 ) ,
    .IN ( config0_decoder11.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U19.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n54 ) ) ;
and ( 
    .Z ( config0_decoder11.U19.ZN ) ,
    .I0 ( config0_decoder11.U19.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_2 ) ,
    .IN ( config0_decoder11.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U16.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n58 ) ) ;
and ( 
    .Z ( config0_decoder11.U16.ZN ) ,
    .I0 ( config0_decoder11.U16.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_6 ) ,
    .IN ( config0_decoder11.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U36.AB ) ,
    .I0 ( config0_decoder11.n56 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U36.ZN ) ,
    .I0 ( config0_decoder11.U36.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_35 ) ,
    .IN ( config0_decoder11.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U1.AB ) ,
    .I0 ( config0_decoder11.n47 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U1.ZN ) ,
    .I0 ( config0_decoder11.U1.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_28 ) ,
    .IN ( config0_decoder11.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U84.AB ) ,
    .I0 ( config0_decoder11.n48 ) ,
    .I1 ( config0_decoder11.n47 ) ) ;
and ( 
    .Z ( config0_decoder11.U84.ZN ) ,
    .I0 ( config0_decoder11.U84.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_43 ) ,
    .IN ( config0_decoder11.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U56.AB ) ,
    .I0 ( config0_decoder11.n50 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U56.ZN ) ,
    .I0 ( config0_decoder11.U56.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_45 ) ,
    .IN ( config0_decoder11.U56.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n44 ) ,
    .I0 ( config0_decoder11.n37 ) ,
    .I1 ( masks_hold_reg_9_3 ) ) ;
or ( 
    .Z ( config0_decoder11.U76.AB ) ,
    .I0 ( config0_decoder11.n53 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U76.ZN ) ,
    .I0 ( config0_decoder11.U76.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_15 ) ,
    .IN ( config0_decoder11.U76.ZN ) ) ;
not ( 
    .O1 ( config0_decoder11.n45 ) ,
    .IN ( masks_hold_reg_9_8 ) ) ;
or ( 
    .Z ( config0_decoder11.U17.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n53 ) ) ;
and ( 
    .Z ( config0_decoder11.U17.ZN ) ,
    .I0 ( config0_decoder11.U17.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_0 ) ,
    .IN ( config0_decoder11.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U37.AB ) ,
    .I0 ( config0_decoder11.n47 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U37.ZN ) ,
    .I0 ( config0_decoder11.U37.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_27 ) ,
    .IN ( config0_decoder11.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U87.AB ) ,
    .I0 ( config0_decoder11.n57 ) ,
    .I1 ( config0_decoder11.n54 ) ) ;
and ( 
    .Z ( config0_decoder11.U87.ZN ) ,
    .I0 ( config0_decoder11.U87.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_50 ) ,
    .IN ( config0_decoder11.U87.ZN ) ) ;
not ( 
    .O1 ( config0_decoder11.n39 ) ,
    .IN ( masks_hold_reg_9_6 ) ) ;
nand ( 
    .Z ( config0_decoder11.n57 ) ,
    .I0 ( masks_hold_reg_9_3 ) ,
    .I1 ( config0_decoder11.n52 ) ) ;
or ( 
    .Z ( config0_decoder11.U77.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n47 ) ) ;
and ( 
    .Z ( config0_decoder11.U77.ZN ) ,
    .I0 ( config0_decoder11.U77.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_11 ) ,
    .IN ( config0_decoder11.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U67.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n50 ) ) ;
and ( 
    .Z ( config0_decoder11.U67.ZN ) ,
    .I0 ( config0_decoder11.U67.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_14 ) ,
    .IN ( config0_decoder11.U67.ZN ) ) ;
nor ( 
    .Z ( config0_decoder11.n52 ) ,
    .I0 ( config0_decoder11.n45 ) ,
    .I1 ( config0_decoder11.n36 ) ) ;
or ( 
    .Z ( config0_decoder11.U34.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U34.ZN ) ,
    .I0 ( config0_decoder11.U34.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_25 ) ,
    .IN ( config0_decoder11.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U3.AB ) ,
    .I0 ( config0_decoder11.n50 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U3.ZN ) ,
    .I0 ( config0_decoder11.U3.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_30 ) ,
    .IN ( config0_decoder11.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U86.AB ) ,
    .I0 ( config0_decoder11.n57 ) ,
    .I1 ( config0_decoder11.n56 ) ) ;
and ( 
    .Z ( config0_decoder11.U86.ZN ) ,
    .I0 ( config0_decoder11.U86.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_52 ) ,
    .IN ( config0_decoder11.U86.ZN ) ) ;
and ( 
    .Z ( config0_decoder11.n40 ) ,
    .I0 ( masks_hold_reg_9_5 ) ,
    .I1 ( masks_hold_reg_9_4 ) ) ;
nand ( 
    .Z ( config0_decoder11.n50 ) ,
    .I0 ( config0_decoder11.n40 ) ,
    .I1 ( masks_hold_reg_9_6 ) ) ;
or ( 
    .Z ( config0_decoder11.U74.AB ) ,
    .I0 ( config0_decoder11.n54 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U74.ZN ) ,
    .I0 ( config0_decoder11.U74.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_18 ) ,
    .IN ( config0_decoder11.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U66.AB ) ,
    .I0 ( config0_decoder11.n56 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U66.ZN ) ,
    .I0 ( config0_decoder11.U66.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_36 ) ,
    .IN ( config0_decoder11.U66.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n55 ) ,
    .I0 ( config0_decoder11.n52 ) ,
    .I1 ( config0_decoder11.n51 ) ) ;
or ( 
    .Z ( config0_decoder11.U35.AB ) ,
    .I0 ( config0_decoder11.n58 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U35.ZN ) ,
    .I0 ( config0_decoder11.U35.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_37 ) ,
    .IN ( config0_decoder11.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U2.AB ) ,
    .I0 ( config0_decoder11.n53 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U2.ZN ) ,
    .I0 ( config0_decoder11.U2.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_31 ) ,
    .IN ( config0_decoder11.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U81.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n62 ) ) ;
and ( 
    .Z ( config0_decoder11.U81.ZN ) ,
    .I0 ( config0_decoder11.U81.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_9 ) ,
    .IN ( config0_decoder11.U81.ZN ) ) ;
not ( 
    .O1 ( config0_decoder11.n36 ) ,
    .IN ( masks_hold_reg_9_7 ) ) ;
not ( 
    .O1 ( config0_decoder11.n51 ) ,
    .IN ( masks_hold_reg_9_3 ) ) ;
or ( 
    .Z ( config0_decoder11.U75.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U75.ZN ) ,
    .I0 ( config0_decoder11.U75.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_42 ) ,
    .IN ( config0_decoder11.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U65.AB ) ,
    .I0 ( config0_decoder11.n55 ) ,
    .I1 ( config0_decoder11.n53 ) ) ;
and ( 
    .Z ( config0_decoder11.U65.ZN ) ,
    .I0 ( config0_decoder11.U65.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_47 ) ,
    .IN ( config0_decoder11.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U12.AB ) ,
    .I0 ( config0_decoder11.n58 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U12.ZN ) ,
    .I0 ( config0_decoder11.U12.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_22 ) ,
    .IN ( config0_decoder11.U12.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n56 ) ,
    .I0 ( config0_decoder11.n41 ) ,
    .I1 ( config0_decoder11.n39 ) ,
    .I2 ( masks_hold_reg_9_5 ) ) ;
or ( 
    .Z ( config0_decoder11.U32.AB ) ,
    .I0 ( config0_decoder11.n50 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U32.ZN ) ,
    .I0 ( config0_decoder11.U32.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_29 ) ,
    .IN ( config0_decoder11.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U29.AB ) ,
    .I0 ( config0_decoder11.n53 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U29.ZN ) ,
    .I0 ( config0_decoder11.U29.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_32 ) ,
    .IN ( config0_decoder11.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U80.AB ) ,
    .I0 ( config0_decoder11.n60 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U80.ZN ) ,
    .I0 ( config0_decoder11.U80.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_39 ) ,
    .IN ( config0_decoder11.U80.ZN ) ) ;
nor ( 
    .Z ( config0_decoder11.n38 ) ,
    .I0 ( masks_hold_reg_9_5 ) ,
    .I1 ( masks_hold_reg_9_6 ) ) ;
or ( 
    .Z ( config0_decoder11.U64.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n54 ) ) ;
and ( 
    .Z ( config0_decoder11.U64.ZN ) ,
    .I0 ( config0_decoder11.U64.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_1 ) ,
    .IN ( config0_decoder11.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U13.AB ) ,
    .I0 ( config0_decoder11.n60 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U13.ZN ) ,
    .I0 ( config0_decoder11.U13.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_23 ) ,
    .IN ( config0_decoder11.U13.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U33.AB ) ,
    .I0 ( config0_decoder11.n54 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U33.ZN ) ,
    .I0 ( config0_decoder11.U33.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_33 ) ,
    .IN ( config0_decoder11.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U28.AB ) ,
    .I0 ( config0_decoder11.n60 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U28.ZN ) ,
    .I0 ( config0_decoder11.U28.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_24 ) ,
    .IN ( config0_decoder11.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U83.AB ) ,
    .I0 ( config0_decoder11.n56 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U83.ZN ) ,
    .I0 ( config0_decoder11.U83.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_19 ) ,
    .IN ( config0_decoder11.U83.ZN ) ) ;
nor ( 
    .Z ( config0_decoder11.n35 ) ,
    .I0 ( masks_hold_reg_9_7 ) ,
    .I1 ( masks_hold_reg_9_8 ) ) ;
or ( 
    .Z ( config0_decoder11.U30.AB ) ,
    .I0 ( config0_decoder11.n54 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U30.ZN ) ,
    .I0 ( config0_decoder11.U30.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_34 ) ,
    .IN ( config0_decoder11.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U22.AB ) ,
    .I0 ( config0_decoder11.n56 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U22.ZN ) ,
    .I0 ( config0_decoder11.U22.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_20 ) ,
    .IN ( config0_decoder11.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U82.AB ) ,
    .I0 ( config0_decoder11.n62 ) ,
    .I1 ( config0_decoder11.n50 ) ) ;
and ( 
    .Z ( config0_decoder11.U82.ZN ) ,
    .I0 ( config0_decoder11.U82.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_13 ) ,
    .IN ( config0_decoder11.U82.ZN ) ) ;
nor ( 
    .Z ( config0_decoder11.n42 ) ,
    .I0 ( config0_decoder11.n39 ) ,
    .I1 ( masks_hold_reg_9_5 ) ) ;
nand ( 
    .Z ( config0_decoder11.n59 ) ,
    .I0 ( masks_hold_reg_9_3 ) ,
    .I1 ( config0_decoder11.n35 ) ) ;
or ( 
    .Z ( config0_decoder11.U78.AB ) ,
    .I0 ( config0_decoder11.n54 ) ,
    .I1 ( config0_decoder11.n43 ) ) ;
and ( 
    .Z ( config0_decoder11.U78.ZN ) ,
    .I0 ( config0_decoder11.U78.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_17 ) ,
    .IN ( config0_decoder11.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U31.AB ) ,
    .I0 ( config0_decoder11.n58 ) ,
    .I1 ( config0_decoder11.n49 ) ) ;
and ( 
    .Z ( config0_decoder11.U31.ZN ) ,
    .I0 ( config0_decoder11.U31.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_38 ) ,
    .IN ( config0_decoder11.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U21.AB ) ,
    .I0 ( config0_decoder11.n55 ) ,
    .I1 ( config0_decoder11.n54 ) ) ;
and ( 
    .Z ( config0_decoder11.U21.ZN ) ,
    .I0 ( config0_decoder11.U21.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_49 ) ,
    .IN ( config0_decoder11.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n43 ) ,
    .I0 ( config0_decoder11.n37 ) ,
    .I1 ( config0_decoder11.n51 ) ) ;
not ( 
    .O1 ( config0_decoder11.n41 ) ,
    .IN ( masks_hold_reg_9_4 ) ) ;
nand ( 
    .Z ( config0_decoder11.n47 ) ,
    .I0 ( masks_hold_reg_9_6 ) ,
    .I1 ( config0_decoder11.n41 ) ,
    .I2 ( masks_hold_reg_9_5 ) ) ;
or ( 
    .Z ( config0_decoder11.U79.AB ) ,
    .I0 ( config0_decoder11.n63 ) ,
    .I1 ( config0_decoder11.n48 ) ) ;
and ( 
    .Z ( config0_decoder11.U79.ZN ) ,
    .I0 ( config0_decoder11.U79.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_41 ) ,
    .IN ( config0_decoder11.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U72.AB ) ,
    .I0 ( config0_decoder11.n60 ) ,
    .I1 ( config0_decoder11.n59 ) ) ;
and ( 
    .Z ( config0_decoder11.U72.ZN ) ,
    .I0 ( config0_decoder11.U72.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_8 ) ,
    .IN ( config0_decoder11.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U69.AB ) ,
    .I0 ( config0_decoder11.n53 ) ,
    .I1 ( config0_decoder11.n44 ) ) ;
and ( 
    .Z ( config0_decoder11.U69.ZN ) ,
    .I0 ( config0_decoder11.U69.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_16 ) ,
    .IN ( config0_decoder11.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder11.U20.AB ) ,
    .I0 ( config0_decoder11.n57 ) ,
    .I1 ( config0_decoder11.n53 ) ) ;
and ( 
    .Z ( config0_decoder11.U20.ZN ) ,
    .I0 ( config0_decoder11.U20.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_48 ) ,
    .IN ( config0_decoder11.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder11.n58 ) ,
    .I0 ( config0_decoder11.n40 ) ,
    .I1 ( config0_decoder11.n39 ) ) ;
nand ( 
    .Z ( config0_decoder11.n48 ) ,
    .I0 ( config0_decoder11.n46 ) ,
    .I1 ( config0_decoder11.n51 ) ) ;
nor ( 
    .Z ( config0_decoder11.n37 ) ,
    .I0 ( config0_decoder11.n36 ) ,
    .I1 ( masks_hold_reg_9_8 ) ) ;
nand ( 
    .Z ( config0_decoder11.n49 ) ,
    .I0 ( config0_decoder11.n46 ) ,
    .I1 ( masks_hold_reg_9_3 ) ) ;
or ( 
    .Z ( config0_decoder11.U73.AB ) ,
    .I0 ( config0_decoder11.n59 ) ,
    .I1 ( config0_decoder11.n47 ) ) ;
and ( 
    .Z ( config0_decoder11.U73.ZN ) ,
    .I0 ( config0_decoder11.U73.AB ) ,
    .I1 ( config0_decoder11.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_10_12 ) ,
    .IN ( config0_decoder11.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U28.AB ) ,
    .I0 ( config0_decoder14.n40 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
and ( 
    .Z ( config0_decoder14.U28.ZN ) ,
    .I0 ( config0_decoder14.U28.AB ) ,
    .I1 ( config0_decoder14.n52 ) ) ;
not ( 
    .O1 ( config0_decoder14.n1 ) ,
    .IN ( config0_decoder14.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U68.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U68.ZN ) ,
    .I0 ( config0_decoder14.U68.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_42 ) ,
    .IN ( config0_decoder14.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U63.AB ) ,
    .I0 ( config0_decoder14.n54 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U63.ZN ) ,
    .I0 ( config0_decoder14.U63.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_34 ) ,
    .IN ( config0_decoder14.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U14.AB ) ,
    .I0 ( config0_decoder14.n54 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U14.ZN ) ,
    .I0 ( config0_decoder14.U14.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_18 ) ,
    .IN ( config0_decoder14.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n55 ) ,
    .I0 ( config0_decoder14.n52 ) ,
    .I1 ( config0_decoder14.n51 ) ) ;
nor ( 
    .Z ( config0_decoder14.n52 ) ,
    .I0 ( config0_decoder14.n45 ) ,
    .I1 ( config0_decoder14.n36 ) ) ;
or ( 
    .Z ( config0_decoder14.U54.AB ) ,
    .I0 ( config0_decoder14.n49 ) ,
    .I1 ( config0_decoder14.n47 ) ) ;
and ( 
    .Z ( config0_decoder14.U54.ZN ) ,
    .I0 ( config0_decoder14.U54.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_44 ) ,
    .IN ( config0_decoder14.U54.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n57 ) ,
    .I0 ( masks_hold_reg_12_6 ) ,
    .I1 ( config0_decoder14.n52 ) ) ;
or ( 
    .Z ( config0_decoder14.U70.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U70.ZN ) ,
    .I0 ( config0_decoder14.U70.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_25 ) ,
    .IN ( config0_decoder14.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U62.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U62.ZN ) ,
    .I0 ( config0_decoder14.U62.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_26 ) ,
    .IN ( config0_decoder14.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U18.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n58 ) ) ;
and ( 
    .Z ( config0_decoder14.U18.ZN ) ,
    .I0 ( config0_decoder14.U18.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_6 ) ,
    .IN ( config0_decoder14.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U15.AB ) ,
    .I0 ( config0_decoder14.n56 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U15.ZN ) ,
    .I0 ( config0_decoder14.U15.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_19 ) ,
    .IN ( config0_decoder14.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n58 ) ,
    .I0 ( config0_decoder14.n40 ) ,
    .I1 ( config0_decoder14.n39 ) ) ;
or ( 
    .Z ( config0_decoder14.U85.AB ) ,
    .I0 ( config0_decoder14.n56 ) ,
    .I1 ( config0_decoder14.n55 ) ) ;
and ( 
    .Z ( config0_decoder14.U85.ZN ) ,
    .I0 ( config0_decoder14.U85.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_51 ) ,
    .IN ( config0_decoder14.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U55.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n58 ) ) ;
and ( 
    .Z ( config0_decoder14.U55.ZN ) ,
    .I0 ( config0_decoder14.U55.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_5 ) ,
    .IN ( config0_decoder14.U55.ZN ) ) ;
not ( 
    .O1 ( config0_decoder14.n51 ) ,
    .IN ( masks_hold_reg_12_6 ) ) ;
or ( 
    .Z ( config0_decoder14.U71.AB ) ,
    .I0 ( config0_decoder14.n54 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U71.ZN ) ,
    .I0 ( config0_decoder14.U71.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_33 ) ,
    .IN ( config0_decoder14.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U61.AB ) ,
    .I0 ( config0_decoder14.n60 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U61.ZN ) ,
    .I0 ( config0_decoder14.U61.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_40 ) ,
    .IN ( config0_decoder14.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U19.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n56 ) ) ;
and ( 
    .Z ( config0_decoder14.U19.ZN ) ,
    .I0 ( config0_decoder14.U19.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_3 ) ,
    .IN ( config0_decoder14.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U16.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n56 ) ) ;
and ( 
    .Z ( config0_decoder14.U16.ZN ) ,
    .I0 ( config0_decoder14.U16.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_4 ) ,
    .IN ( config0_decoder14.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n44 ) ,
    .I0 ( config0_decoder14.n37 ) ,
    .I1 ( masks_hold_reg_12_6 ) ) ;
nand ( 
    .Z ( config0_decoder14.n48 ) ,
    .I0 ( config0_decoder14.n46 ) ,
    .I1 ( config0_decoder14.n51 ) ) ;
or ( 
    .Z ( config0_decoder14.U84.AB ) ,
    .I0 ( config0_decoder14.n48 ) ,
    .I1 ( config0_decoder14.n47 ) ) ;
and ( 
    .Z ( config0_decoder14.U84.ZN ) ,
    .I0 ( config0_decoder14.U84.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_43 ) ,
    .IN ( config0_decoder14.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U56.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n54 ) ) ;
and ( 
    .Z ( config0_decoder14.U56.ZN ) ,
    .I0 ( config0_decoder14.U56.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_1 ) ,
    .IN ( config0_decoder14.U56.ZN ) ) ;
not ( 
    .O1 ( config0_decoder14.n41 ) ,
    .IN ( masks_hold_reg_12_7 ) ) ;
or ( 
    .Z ( config0_decoder14.U76.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n47 ) ) ;
and ( 
    .Z ( config0_decoder14.U76.ZN ) ,
    .I0 ( config0_decoder14.U76.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_11 ) ,
    .IN ( config0_decoder14.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U60.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n50 ) ) ;
and ( 
    .Z ( config0_decoder14.U60.ZN ) ,
    .I0 ( config0_decoder14.U60.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_14 ) ,
    .IN ( config0_decoder14.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U17.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n60 ) ) ;
and ( 
    .Z ( config0_decoder14.U17.ZN ) ,
    .I0 ( config0_decoder14.U17.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_7 ) ,
    .IN ( config0_decoder14.U17.ZN ) ) ;
nor ( 
    .Z ( config0_decoder14.n35 ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( masks_hold_reg_11_0 ) ) ;
or ( 
    .Z ( config0_decoder14.U87.AB ) ,
    .I0 ( config0_decoder14.n57 ) ,
    .I1 ( config0_decoder14.n54 ) ) ;
and ( 
    .Z ( config0_decoder14.U87.ZN ) ,
    .I0 ( config0_decoder14.U87.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_50 ) ,
    .IN ( config0_decoder14.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U57.AB ) ,
    .I0 ( config0_decoder14.n60 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U57.ZN ) ,
    .I0 ( config0_decoder14.U57.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_24 ) ,
    .IN ( config0_decoder14.U57.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U47.AB ) ,
    .I0 ( config0_decoder14.n53 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U47.ZN ) ,
    .I0 ( config0_decoder14.U47.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_32 ) ,
    .IN ( config0_decoder14.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U77.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U77.ZN ) ,
    .I0 ( config0_decoder14.U77.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_41 ) ,
    .IN ( config0_decoder14.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U67.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n47 ) ) ;
and ( 
    .Z ( config0_decoder14.U67.ZN ) ,
    .I0 ( config0_decoder14.U67.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_12 ) ,
    .IN ( config0_decoder14.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U10.AB ) ,
    .I0 ( config0_decoder14.n53 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U10.ZN ) ,
    .I0 ( config0_decoder14.U10.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_16 ) ,
    .IN ( config0_decoder14.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n63 ) ,
    .I0 ( masks_hold_reg_12_7 ) ,
    .I1 ( config0_decoder14.n42 ) ) ;
nand ( 
    .Z ( config0_decoder14.n43 ) ,
    .I0 ( config0_decoder14.n37 ) ,
    .I1 ( config0_decoder14.n51 ) ) ;
or ( 
    .Z ( config0_decoder14.U86.AB ) ,
    .I0 ( config0_decoder14.n57 ) ,
    .I1 ( config0_decoder14.n56 ) ) ;
and ( 
    .Z ( config0_decoder14.U86.ZN ) ,
    .I0 ( config0_decoder14.U86.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_52 ) ,
    .IN ( config0_decoder14.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U58.AB ) ,
    .I0 ( config0_decoder14.n56 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U58.ZN ) ,
    .I0 ( config0_decoder14.U58.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_36 ) ,
    .IN ( config0_decoder14.U58.ZN ) ) ;
nor ( 
    .Z ( config0_decoder14.n37 ) ,
    .I0 ( config0_decoder14.n36 ) ,
    .I1 ( masks_hold_reg_11_0 ) ) ;
or ( 
    .Z ( config0_decoder14.U74.AB ) ,
    .I0 ( config0_decoder14.n58 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U74.ZN ) ,
    .I0 ( config0_decoder14.U74.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_21 ) ,
    .IN ( config0_decoder14.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U66.AB ) ,
    .I0 ( config0_decoder14.n60 ) ,
    .I1 ( config0_decoder14.n59 ) ) ;
and ( 
    .Z ( config0_decoder14.U66.ZN ) ,
    .I0 ( config0_decoder14.U66.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_8 ) ,
    .IN ( config0_decoder14.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U11.AB ) ,
    .I0 ( config0_decoder14.n47 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U11.ZN ) ,
    .I0 ( config0_decoder14.U11.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_28 ) ,
    .IN ( config0_decoder14.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder14.n46 ) ,
    .I0 ( config0_decoder14.n45 ) ,
    .I1 ( masks_hold_reg_12_10 ) ) ;
nand ( 
    .Z ( config0_decoder14.n49 ) ,
    .I0 ( config0_decoder14.n46 ) ,
    .I1 ( masks_hold_reg_12_6 ) ) ;
nand ( 
    .Z ( config0_decoder14.n62 ) ,
    .I0 ( config0_decoder14.n35 ) ,
    .I1 ( config0_decoder14.n51 ) ) ;
or ( 
    .Z ( config0_decoder14.U81.AB ) ,
    .I0 ( config0_decoder14.n60 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U81.ZN ) ,
    .I0 ( config0_decoder14.U81.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_23 ) ,
    .IN ( config0_decoder14.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U59.AB ) ,
    .I0 ( config0_decoder14.n56 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U59.ZN ) ,
    .I0 ( config0_decoder14.U59.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_20 ) ,
    .IN ( config0_decoder14.U59.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U49.AB ) ,
    .I0 ( config0_decoder14.n55 ) ,
    .I1 ( config0_decoder14.n53 ) ) ;
and ( 
    .Z ( config0_decoder14.U49.ZN ) ,
    .I0 ( config0_decoder14.U49.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_47 ) ,
    .IN ( config0_decoder14.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U75.AB ) ,
    .I0 ( config0_decoder14.n53 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U75.ZN ) ,
    .I0 ( config0_decoder14.U75.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_15 ) ,
    .IN ( config0_decoder14.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U65.AB ) ,
    .I0 ( config0_decoder14.n58 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U65.ZN ) ,
    .I0 ( config0_decoder14.U65.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_22 ) ,
    .IN ( config0_decoder14.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U12.AB ) ,
    .I0 ( config0_decoder14.n50 ) ,
    .I1 ( config0_decoder14.n44 ) ) ;
and ( 
    .Z ( config0_decoder14.U12.ZN ) ,
    .I0 ( config0_decoder14.U12.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_30 ) ,
    .IN ( config0_decoder14.U12.ZN ) ) ;
nor ( 
    .Z ( config0_decoder14.n38 ) ,
    .I0 ( masks_hold_reg_12_8 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
nand ( 
    .Z ( config0_decoder14.n50 ) ,
    .I0 ( config0_decoder14.n40 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
nand ( 
    .Z ( config0_decoder14.n56 ) ,
    .I0 ( config0_decoder14.n41 ) ,
    .I1 ( config0_decoder14.n39 ) ,
    .I2 ( masks_hold_reg_12_8 ) ) ;
or ( 
    .Z ( config0_decoder14.U80.AB ) ,
    .I0 ( config0_decoder14.n60 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U80.ZN ) ,
    .I0 ( config0_decoder14.U80.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_39 ) ,
    .IN ( config0_decoder14.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U48.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n59 ) ) ;
and ( 
    .Z ( config0_decoder14.U48.ZN ) ,
    .I0 ( config0_decoder14.U48.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_10 ) ,
    .IN ( config0_decoder14.U48.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U64.AB ) ,
    .I0 ( config0_decoder14.n58 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U64.ZN ) ,
    .I0 ( config0_decoder14.U64.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_38 ) ,
    .IN ( config0_decoder14.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U13.AB ) ,
    .I0 ( config0_decoder14.n53 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U13.ZN ) ,
    .I0 ( config0_decoder14.U13.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_31 ) ,
    .IN ( config0_decoder14.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n54 ) ,
    .I0 ( config0_decoder14.n38 ) ,
    .I1 ( masks_hold_reg_12_7 ) ) ;
or ( 
    .Z ( config0_decoder14.U83.AB ) ,
    .I0 ( config0_decoder14.n62 ) ,
    .I1 ( config0_decoder14.n50 ) ) ;
and ( 
    .Z ( config0_decoder14.U83.ZN ) ,
    .I0 ( config0_decoder14.U83.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_13 ) ,
    .IN ( config0_decoder14.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U50.AB ) ,
    .I0 ( config0_decoder14.n50 ) ,
    .I1 ( config0_decoder14.n49 ) ) ;
and ( 
    .Z ( config0_decoder14.U50.ZN ) ,
    .I0 ( config0_decoder14.U50.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_46 ) ,
    .IN ( config0_decoder14.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n47 ) ,
    .I0 ( masks_hold_reg_12_9 ) ,
    .I1 ( config0_decoder14.n41 ) ,
    .I2 ( masks_hold_reg_12_8 ) ) ;
or ( 
    .Z ( config0_decoder14.U22.AB ) ,
    .I0 ( config0_decoder14.n55 ) ,
    .I1 ( config0_decoder14.n54 ) ) ;
and ( 
    .Z ( config0_decoder14.U22.ZN ) ,
    .I0 ( config0_decoder14.U22.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_49 ) ,
    .IN ( config0_decoder14.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U82.AB ) ,
    .I0 ( config0_decoder14.n63 ) ,
    .I1 ( config0_decoder14.n62 ) ) ;
and ( 
    .Z ( config0_decoder14.U82.ZN ) ,
    .I0 ( config0_decoder14.U82.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_9 ) ,
    .IN ( config0_decoder14.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U51.AB ) ,
    .I0 ( config0_decoder14.n50 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U51.ZN ) ,
    .I0 ( config0_decoder14.U51.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_45 ) ,
    .IN ( config0_decoder14.U51.ZN ) ) ;
not ( 
    .O1 ( config0_decoder14.n36 ) ,
    .IN ( masks_hold_reg_12_10 ) ) ;
or ( 
    .Z ( config0_decoder14.U78.AB ) ,
    .I0 ( config0_decoder14.n47 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U78.ZN ) ,
    .I0 ( config0_decoder14.U78.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_27 ) ,
    .IN ( config0_decoder14.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n59 ) ,
    .I0 ( masks_hold_reg_12_6 ) ,
    .I1 ( config0_decoder14.n35 ) ) ;
or ( 
    .Z ( config0_decoder14.U21.AB ) ,
    .I0 ( config0_decoder14.n57 ) ,
    .I1 ( config0_decoder14.n53 ) ) ;
and ( 
    .Z ( config0_decoder14.U21.ZN ) ,
    .I0 ( config0_decoder14.U21.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_48 ) ,
    .IN ( config0_decoder14.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n60 ) ,
    .I0 ( config0_decoder14.n42 ) ,
    .I1 ( config0_decoder14.n41 ) ) ;
and ( 
    .Z ( config0_decoder14.n40 ) ,
    .I0 ( masks_hold_reg_12_8 ) ,
    .I1 ( masks_hold_reg_12_7 ) ) ;
not ( 
    .O1 ( config0_decoder14.n39 ) ,
    .IN ( masks_hold_reg_12_9 ) ) ;
or ( 
    .Z ( config0_decoder14.U79.AB ) ,
    .I0 ( config0_decoder14.n56 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U79.ZN ) ,
    .I0 ( config0_decoder14.U79.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_35 ) ,
    .IN ( config0_decoder14.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U72.AB ) ,
    .I0 ( config0_decoder14.n58 ) ,
    .I1 ( config0_decoder14.n48 ) ) ;
and ( 
    .Z ( config0_decoder14.U72.ZN ) ,
    .I0 ( config0_decoder14.U72.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_37 ) ,
    .IN ( config0_decoder14.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U69.AB ) ,
    .I0 ( config0_decoder14.n50 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U69.ZN ) ,
    .I0 ( config0_decoder14.U69.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_29 ) ,
    .IN ( config0_decoder14.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U20.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n54 ) ) ;
and ( 
    .Z ( config0_decoder14.U20.ZN ) ,
    .I0 ( config0_decoder14.U20.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_2 ) ,
    .IN ( config0_decoder14.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder14.U9.AB ) ,
    .I0 ( config0_decoder14.n59 ) ,
    .I1 ( config0_decoder14.n53 ) ) ;
and ( 
    .Z ( config0_decoder14.U9.ZN ) ,
    .I0 ( config0_decoder14.U9.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_0 ) ,
    .IN ( config0_decoder14.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder14.n53 ) ,
    .I0 ( config0_decoder14.n38 ) ,
    .I1 ( config0_decoder14.n41 ) ) ;
not ( 
    .O1 ( config0_decoder14.n45 ) ,
    .IN ( masks_hold_reg_11_0 ) ) ;
nor ( 
    .Z ( config0_decoder14.n42 ) ,
    .I0 ( config0_decoder14.n39 ) ,
    .I1 ( masks_hold_reg_12_8 ) ) ;
or ( 
    .Z ( config0_decoder14.U73.AB ) ,
    .I0 ( config0_decoder14.n54 ) ,
    .I1 ( config0_decoder14.n43 ) ) ;
and ( 
    .Z ( config0_decoder14.U73.ZN ) ,
    .I0 ( config0_decoder14.U73.AB ) ,
    .I1 ( config0_decoder14.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_13_17 ) ,
    .IN ( config0_decoder14.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U42.AB ) ,
    .I0 ( config0_decoder15.n40 ) ,
    .I1 ( masks_hold_reg_13_7 ) ) ;
and ( 
    .Z ( config0_decoder15.U42.ZN ) ,
    .I0 ( config0_decoder15.U42.AB ) ,
    .I1 ( config0_decoder15.n52 ) ) ;
not ( 
    .O1 ( config0_decoder15.n1 ) ,
    .IN ( config0_decoder15.U42.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U68.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n58 ) ) ;
and ( 
    .Z ( config0_decoder15.U68.ZN ) ,
    .I0 ( config0_decoder15.U68.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_5 ) ,
    .IN ( config0_decoder15.U68.ZN ) ) ;
and ( 
    .Z ( config0_decoder15.n40 ) ,
    .I0 ( masks_hold_reg_13_6 ) ,
    .I1 ( masks_hold_reg_13_5 ) ) ;
or ( 
    .Z ( config0_decoder15.U14.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n56 ) ) ;
and ( 
    .Z ( config0_decoder15.U14.ZN ) ,
    .I0 ( config0_decoder15.U14.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_4 ) ,
    .IN ( config0_decoder15.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n60 ) ,
    .I0 ( config0_decoder15.n42 ) ,
    .I1 ( config0_decoder15.n41 ) ) ;
nand ( 
    .Z ( config0_decoder15.n53 ) ,
    .I0 ( config0_decoder15.n38 ) ,
    .I1 ( config0_decoder15.n41 ) ) ;
nor ( 
    .Z ( config0_decoder15.n35 ) ,
    .I0 ( masks_hold_reg_12_0 ) ,
    .I1 ( masks_hold_reg_12_1 ) ) ;
or ( 
    .Z ( config0_decoder15.U70.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n50 ) ) ;
and ( 
    .Z ( config0_decoder15.U70.ZN ) ,
    .I0 ( config0_decoder15.U70.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_14 ) ,
    .IN ( config0_decoder15.U70.ZN ) ) ;
not ( 
    .O1 ( config0_decoder15.n39 ) ,
    .IN ( masks_hold_reg_13_7 ) ) ;
or ( 
    .Z ( config0_decoder15.U18.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n56 ) ) ;
and ( 
    .Z ( config0_decoder15.U18.ZN ) ,
    .I0 ( config0_decoder15.U18.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_3 ) ,
    .IN ( config0_decoder15.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U15.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n60 ) ) ;
and ( 
    .Z ( config0_decoder15.U15.ZN ) ,
    .I0 ( config0_decoder15.U15.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_7 ) ,
    .IN ( config0_decoder15.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n62 ) ,
    .I0 ( config0_decoder15.n35 ) ,
    .I1 ( config0_decoder15.n51 ) ) ;
or ( 
    .Z ( config0_decoder15.U85.AB ) ,
    .I0 ( config0_decoder15.n48 ) ,
    .I1 ( config0_decoder15.n47 ) ) ;
and ( 
    .Z ( config0_decoder15.U85.ZN ) ,
    .I0 ( config0_decoder15.U85.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_43 ) ,
    .IN ( config0_decoder15.U85.ZN ) ) ;
nor ( 
    .Z ( config0_decoder15.n42 ) ,
    .I0 ( config0_decoder15.n39 ) ,
    .I1 ( masks_hold_reg_13_6 ) ) ;
nand ( 
    .Z ( config0_decoder15.n59 ) ,
    .I0 ( masks_hold_reg_13_4 ) ,
    .I1 ( config0_decoder15.n35 ) ) ;
or ( 
    .Z ( config0_decoder15.U71.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n59 ) ) ;
and ( 
    .Z ( config0_decoder15.U71.ZN ) ,
    .I0 ( config0_decoder15.U71.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_10 ) ,
    .IN ( config0_decoder15.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U61.AB ) ,
    .I0 ( config0_decoder15.n56 ) ,
    .I1 ( config0_decoder15.n55 ) ) ;
and ( 
    .Z ( config0_decoder15.U61.ZN ) ,
    .I0 ( config0_decoder15.U61.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_51 ) ,
    .IN ( config0_decoder15.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U19.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n54 ) ) ;
and ( 
    .Z ( config0_decoder15.U19.ZN ) ,
    .I0 ( config0_decoder15.U19.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_2 ) ,
    .IN ( config0_decoder15.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U16.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n58 ) ) ;
and ( 
    .Z ( config0_decoder15.U16.ZN ) ,
    .I0 ( config0_decoder15.U16.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_6 ) ,
    .IN ( config0_decoder15.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U36.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U36.ZN ) ,
    .I0 ( config0_decoder15.U36.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_25 ) ,
    .IN ( config0_decoder15.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U1.AB ) ,
    .I0 ( config0_decoder15.n53 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U1.ZN ) ,
    .I0 ( config0_decoder15.U1.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_31 ) ,
    .IN ( config0_decoder15.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U84.AB ) ,
    .I0 ( config0_decoder15.n56 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U84.ZN ) ,
    .I0 ( config0_decoder15.U84.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_19 ) ,
    .IN ( config0_decoder15.U84.ZN ) ) ;
not ( 
    .O1 ( config0_decoder15.n41 ) ,
    .IN ( masks_hold_reg_13_5 ) ) ;
nand ( 
    .Z ( config0_decoder15.n47 ) ,
    .I0 ( masks_hold_reg_13_7 ) ,
    .I1 ( config0_decoder15.n41 ) ,
    .I2 ( masks_hold_reg_13_6 ) ) ;
or ( 
    .Z ( config0_decoder15.U76.AB ) ,
    .I0 ( config0_decoder15.n54 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U76.ZN ) ,
    .I0 ( config0_decoder15.U76.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_18 ) ,
    .IN ( config0_decoder15.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U60.AB ) ,
    .I0 ( config0_decoder15.n50 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U60.ZN ) ,
    .I0 ( config0_decoder15.U60.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_46 ) ,
    .IN ( config0_decoder15.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U17.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n53 ) ) ;
and ( 
    .Z ( config0_decoder15.U17.ZN ) ,
    .I0 ( config0_decoder15.U17.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_0 ) ,
    .IN ( config0_decoder15.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U37.AB ) ,
    .I0 ( config0_decoder15.n58 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U37.ZN ) ,
    .I0 ( config0_decoder15.U37.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_37 ) ,
    .IN ( config0_decoder15.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U87.AB ) ,
    .I0 ( config0_decoder15.n57 ) ,
    .I1 ( config0_decoder15.n54 ) ) ;
and ( 
    .Z ( config0_decoder15.U87.ZN ) ,
    .I0 ( config0_decoder15.U87.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_50 ) ,
    .IN ( config0_decoder15.U87.ZN ) ) ;
nor ( 
    .Z ( config0_decoder15.n37 ) ,
    .I0 ( config0_decoder15.n36 ) ,
    .I1 ( masks_hold_reg_12_1 ) ) ;
nand ( 
    .Z ( config0_decoder15.n49 ) ,
    .I0 ( config0_decoder15.n46 ) ,
    .I1 ( masks_hold_reg_13_4 ) ) ;
or ( 
    .Z ( config0_decoder15.U77.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U77.ZN ) ,
    .I0 ( config0_decoder15.U77.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_42 ) ,
    .IN ( config0_decoder15.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U67.AB ) ,
    .I0 ( config0_decoder15.n50 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U67.ZN ) ,
    .I0 ( config0_decoder15.U67.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_45 ) ,
    .IN ( config0_decoder15.U67.ZN ) ) ;
nor ( 
    .Z ( config0_decoder15.n52 ) ,
    .I0 ( config0_decoder15.n45 ) ,
    .I1 ( config0_decoder15.n36 ) ) ;
or ( 
    .Z ( config0_decoder15.U34.AB ) ,
    .I0 ( config0_decoder15.n50 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U34.ZN ) ,
    .I0 ( config0_decoder15.U34.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_29 ) ,
    .IN ( config0_decoder15.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U3.AB ) ,
    .I0 ( config0_decoder15.n47 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U3.ZN ) ,
    .I0 ( config0_decoder15.U3.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_28 ) ,
    .IN ( config0_decoder15.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U86.AB ) ,
    .I0 ( config0_decoder15.n57 ) ,
    .I1 ( config0_decoder15.n56 ) ) ;
and ( 
    .Z ( config0_decoder15.U86.ZN ) ,
    .I0 ( config0_decoder15.U86.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_52 ) ,
    .IN ( config0_decoder15.U86.ZN ) ) ;
nor ( 
    .Z ( config0_decoder15.n46 ) ,
    .I0 ( config0_decoder15.n45 ) ,
    .I1 ( masks_hold_reg_12_0 ) ) ;
nand ( 
    .Z ( config0_decoder15.n54 ) ,
    .I0 ( config0_decoder15.n38 ) ,
    .I1 ( masks_hold_reg_13_5 ) ) ;
or ( 
    .Z ( config0_decoder15.U74.AB ) ,
    .I0 ( config0_decoder15.n60 ) ,
    .I1 ( config0_decoder15.n59 ) ) ;
and ( 
    .Z ( config0_decoder15.U74.ZN ) ,
    .I0 ( config0_decoder15.U74.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_8 ) ,
    .IN ( config0_decoder15.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U66.AB ) ,
    .I0 ( config0_decoder15.n49 ) ,
    .I1 ( config0_decoder15.n47 ) ) ;
and ( 
    .Z ( config0_decoder15.U66.ZN ) ,
    .I0 ( config0_decoder15.U66.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_44 ) ,
    .IN ( config0_decoder15.U66.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n55 ) ,
    .I0 ( config0_decoder15.n52 ) ,
    .I1 ( config0_decoder15.n51 ) ) ;
or ( 
    .Z ( config0_decoder15.U38.AB ) ,
    .I0 ( config0_decoder15.n58 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U38.ZN ) ,
    .I0 ( config0_decoder15.U38.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_21 ) ,
    .IN ( config0_decoder15.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U35.AB ) ,
    .I0 ( config0_decoder15.n54 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U35.ZN ) ,
    .I0 ( config0_decoder15.U35.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_33 ) ,
    .IN ( config0_decoder15.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U2.AB ) ,
    .I0 ( config0_decoder15.n50 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U2.ZN ) ,
    .I0 ( config0_decoder15.U2.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_30 ) ,
    .IN ( config0_decoder15.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U81.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U81.ZN ) ,
    .I0 ( config0_decoder15.U81.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_41 ) ,
    .IN ( config0_decoder15.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U59.AB ) ,
    .I0 ( config0_decoder15.n55 ) ,
    .I1 ( config0_decoder15.n53 ) ) ;
and ( 
    .Z ( config0_decoder15.U59.ZN ) ,
    .I0 ( config0_decoder15.U59.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_47 ) ,
    .IN ( config0_decoder15.U59.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n63 ) ,
    .I0 ( masks_hold_reg_13_5 ) ,
    .I1 ( config0_decoder15.n42 ) ) ;
or ( 
    .Z ( config0_decoder15.U75.AB ) ,
    .I0 ( config0_decoder15.n59 ) ,
    .I1 ( config0_decoder15.n47 ) ) ;
and ( 
    .Z ( config0_decoder15.U75.ZN ) ,
    .I0 ( config0_decoder15.U75.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_12 ) ,
    .IN ( config0_decoder15.U75.ZN ) ) ;
not ( 
    .O1 ( config0_decoder15.n45 ) ,
    .IN ( masks_hold_reg_12_1 ) ) ;
or ( 
    .Z ( config0_decoder15.U12.AB ) ,
    .I0 ( config0_decoder15.n58 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U12.ZN ) ,
    .I0 ( config0_decoder15.U12.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_22 ) ,
    .IN ( config0_decoder15.U12.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U39.AB ) ,
    .I0 ( config0_decoder15.n56 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U39.ZN ) ,
    .I0 ( config0_decoder15.U39.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_35 ) ,
    .IN ( config0_decoder15.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U32.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U32.ZN ) ,
    .I0 ( config0_decoder15.U32.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_26 ) ,
    .IN ( config0_decoder15.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U29.AB ) ,
    .I0 ( config0_decoder15.n60 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U29.ZN ) ,
    .I0 ( config0_decoder15.U29.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_24 ) ,
    .IN ( config0_decoder15.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U80.AB ) ,
    .I0 ( config0_decoder15.n54 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U80.ZN ) ,
    .I0 ( config0_decoder15.U80.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_17 ) ,
    .IN ( config0_decoder15.U80.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n44 ) ,
    .I0 ( config0_decoder15.n37 ) ,
    .I1 ( masks_hold_reg_13_4 ) ) ;
not ( 
    .O1 ( config0_decoder15.n36 ) ,
    .IN ( masks_hold_reg_12_0 ) ) ;
or ( 
    .Z ( config0_decoder15.U13.AB ) ,
    .I0 ( config0_decoder15.n60 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U13.ZN ) ,
    .I0 ( config0_decoder15.U13.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_23 ) ,
    .IN ( config0_decoder15.U13.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U33.AB ) ,
    .I0 ( config0_decoder15.n58 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U33.ZN ) ,
    .I0 ( config0_decoder15.U33.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_38 ) ,
    .IN ( config0_decoder15.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U28.AB ) ,
    .I0 ( config0_decoder15.n53 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U28.ZN ) ,
    .I0 ( config0_decoder15.U28.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_32 ) ,
    .IN ( config0_decoder15.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U83.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n50 ) ) ;
and ( 
    .Z ( config0_decoder15.U83.ZN ) ,
    .I0 ( config0_decoder15.U83.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_13 ) ,
    .IN ( config0_decoder15.U83.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n50 ) ,
    .I0 ( config0_decoder15.n40 ) ,
    .I1 ( masks_hold_reg_13_7 ) ) ;
or ( 
    .Z ( config0_decoder15.U30.AB ) ,
    .I0 ( config0_decoder15.n56 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U30.ZN ) ,
    .I0 ( config0_decoder15.U30.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_36 ) ,
    .IN ( config0_decoder15.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U22.AB ) ,
    .I0 ( config0_decoder15.n56 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U22.ZN ) ,
    .I0 ( config0_decoder15.U22.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_20 ) ,
    .IN ( config0_decoder15.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U82.AB ) ,
    .I0 ( config0_decoder15.n63 ) ,
    .I1 ( config0_decoder15.n62 ) ) ;
and ( 
    .Z ( config0_decoder15.U82.ZN ) ,
    .I0 ( config0_decoder15.U82.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_9 ) ,
    .IN ( config0_decoder15.U82.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n57 ) ,
    .I0 ( masks_hold_reg_13_4 ) ,
    .I1 ( config0_decoder15.n52 ) ) ;
or ( 
    .Z ( config0_decoder15.U41.AB ) ,
    .I0 ( config0_decoder15.n60 ) ,
    .I1 ( config0_decoder15.n48 ) ) ;
and ( 
    .Z ( config0_decoder15.U41.ZN ) ,
    .I0 ( config0_decoder15.U41.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_39 ) ,
    .IN ( config0_decoder15.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U78.AB ) ,
    .I0 ( config0_decoder15.n53 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U78.ZN ) ,
    .I0 ( config0_decoder15.U78.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_15 ) ,
    .IN ( config0_decoder15.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U31.AB ) ,
    .I0 ( config0_decoder15.n54 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U31.ZN ) ,
    .I0 ( config0_decoder15.U31.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_34 ) ,
    .IN ( config0_decoder15.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U21.AB ) ,
    .I0 ( config0_decoder15.n55 ) ,
    .I1 ( config0_decoder15.n54 ) ) ;
and ( 
    .Z ( config0_decoder15.U21.ZN ) ,
    .I0 ( config0_decoder15.U21.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_49 ) ,
    .IN ( config0_decoder15.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n43 ) ,
    .I0 ( config0_decoder15.n37 ) ,
    .I1 ( config0_decoder15.n51 ) ) ;
nor ( 
    .Z ( config0_decoder15.n38 ) ,
    .I0 ( masks_hold_reg_13_6 ) ,
    .I1 ( masks_hold_reg_13_7 ) ) ;
or ( 
    .Z ( config0_decoder15.U40.AB ) ,
    .I0 ( config0_decoder15.n47 ) ,
    .I1 ( config0_decoder15.n43 ) ) ;
and ( 
    .Z ( config0_decoder15.U40.ZN ) ,
    .I0 ( config0_decoder15.U40.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_27 ) ,
    .IN ( config0_decoder15.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U79.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n47 ) ) ;
and ( 
    .Z ( config0_decoder15.U79.ZN ) ,
    .I0 ( config0_decoder15.U79.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_11 ) ,
    .IN ( config0_decoder15.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U72.AB ) ,
    .I0 ( config0_decoder15.n53 ) ,
    .I1 ( config0_decoder15.n44 ) ) ;
and ( 
    .Z ( config0_decoder15.U72.ZN ) ,
    .I0 ( config0_decoder15.U72.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_16 ) ,
    .IN ( config0_decoder15.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U69.AB ) ,
    .I0 ( config0_decoder15.n62 ) ,
    .I1 ( config0_decoder15.n54 ) ) ;
and ( 
    .Z ( config0_decoder15.U69.ZN ) ,
    .I0 ( config0_decoder15.U69.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_1 ) ,
    .IN ( config0_decoder15.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder15.U20.AB ) ,
    .I0 ( config0_decoder15.n57 ) ,
    .I1 ( config0_decoder15.n53 ) ) ;
and ( 
    .Z ( config0_decoder15.U20.ZN ) ,
    .I0 ( config0_decoder15.U20.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_48 ) ,
    .IN ( config0_decoder15.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder15.n58 ) ,
    .I0 ( config0_decoder15.n40 ) ,
    .I1 ( config0_decoder15.n39 ) ) ;
nand ( 
    .Z ( config0_decoder15.n48 ) ,
    .I0 ( config0_decoder15.n46 ) ,
    .I1 ( config0_decoder15.n51 ) ) ;
not ( 
    .O1 ( config0_decoder15.n51 ) ,
    .IN ( masks_hold_reg_13_4 ) ) ;
nand ( 
    .Z ( config0_decoder15.n56 ) ,
    .I0 ( config0_decoder15.n41 ) ,
    .I1 ( config0_decoder15.n39 ) ,
    .I2 ( masks_hold_reg_13_6 ) ) ;
or ( 
    .Z ( config0_decoder15.U73.AB ) ,
    .I0 ( config0_decoder15.n60 ) ,
    .I1 ( config0_decoder15.n49 ) ) ;
and ( 
    .Z ( config0_decoder15.U73.ZN ) ,
    .I0 ( config0_decoder15.U73.AB ) ,
    .I1 ( config0_decoder15.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_14_40 ) ,
    .IN ( config0_decoder15.U73.ZN ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_10 ) ,
    .IN ( masks_hold_reg_1_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_140 ) ,
    .IN ( masks_hold_reg_12_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_130 ) ,
    .IN ( masks_hold_reg_10_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_100 ) ,
    .IN ( masks_hold_reg_8_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_110 ) ,
    .IN ( masks_hold_reg_9_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_120 ) ,
    .IN ( masks_hold_reg_10_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_70 ) ,
    .IN ( masks_hold_reg_6_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_80 ) ,
    .IN ( masks_hold_reg_6_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_90 ) ,
    .IN ( masks_hold_reg_7_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_60 ) ,
    .IN ( masks_hold_reg_5_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_136 ) ,
    .IN ( masks_hold_reg_12_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_137 ) ,
    .IN ( masks_hold_reg_12_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_30 ) ,
    .IN ( masks_hold_reg_2_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_11 ) ,
    .IN ( masks_hold_reg_1_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_138 ) ,
    .IN ( masks_hold_reg_12_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_13 ) ,
    .IN ( masks_hold_reg_2_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_12 ) ,
    .IN ( masks_hold_reg_2_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_131 ) ,
    .IN ( masks_hold_reg_11_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_141 ) ,
    .IN ( masks_hold_reg_12_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_139 ) ,
    .IN ( masks_hold_reg_12_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_134 ) ,
    .IN ( masks_hold_reg_12_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_133 ) ,
    .IN ( masks_hold_reg_12_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_132 ) ,
    .IN ( masks_hold_reg_11_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_112 ) ,
    .IN ( masks_hold_reg_10_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_121 ) ,
    .IN ( masks_hold_reg_10_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_135 ) ,
    .IN ( masks_hold_reg_12_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_115 ) ,
    .IN ( masks_hold_reg_10_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_114 ) ,
    .IN ( masks_hold_reg_10_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_113 ) ,
    .IN ( masks_hold_reg_10_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_118 ) ,
    .IN ( masks_hold_reg_10_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_117 ) ,
    .IN ( masks_hold_reg_10_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_116 ) ,
    .IN ( masks_hold_reg_10_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_96 ) ,
    .IN ( masks_hold_reg_8_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_111 ) ,
    .IN ( masks_hold_reg_9_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_119 ) ,
    .IN ( masks_hold_reg_10_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_99 ) ,
    .IN ( masks_hold_reg_8_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_98 ) ,
    .IN ( masks_hold_reg_8_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_97 ) ,
    .IN ( masks_hold_reg_8_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_92 ) ,
    .IN ( masks_hold_reg_8_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_91 ) ,
    .IN ( masks_hold_reg_8_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_101 ) ,
    .IN ( masks_hold_reg_8_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_95 ) ,
    .IN ( masks_hold_reg_8_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_94 ) ,
    .IN ( masks_hold_reg_8_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_93 ) ,
    .IN ( masks_hold_reg_8_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_73 ) ,
    .IN ( masks_hold_reg_6_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_72 ) ,
    .IN ( masks_hold_reg_6_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_81 ) ,
    .IN ( masks_hold_reg_7_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_76 ) ,
    .IN ( masks_hold_reg_6_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_75 ) ,
    .IN ( masks_hold_reg_6_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_74 ) ,
    .IN ( masks_hold_reg_6_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_79 ) ,
    .IN ( masks_hold_reg_6_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_78 ) ,
    .IN ( masks_hold_reg_6_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_77 ) ,
    .IN ( masks_hold_reg_6_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_50 ) ,
    .IN ( n92 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_61 ) ,
    .IN ( masks_hold_reg_5_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_71 ) ,
    .IN ( masks_hold_reg_6_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_40 ) ,
    .IN ( masks_hold_reg_3_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_35 ) ,
    .IN ( masks_hold_reg_2_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_34 ) ,
    .IN ( masks_hold_reg_2_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_33 ) ,
    .IN ( masks_hold_reg_2_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_38 ) ,
    .IN ( masks_hold_reg_2_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_37 ) ,
    .IN ( masks_hold_reg_2_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_36 ) ,
    .IN ( masks_hold_reg_2_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_8 ) ,
    .IN ( masks_hold_reg_0_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_31 ) ,
    .IN ( masks_hold_reg_2_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_39 ) ,
    .IN ( masks_hold_reg_3_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_1 ) ,
    .IN ( masks_hold_reg_0_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_0 ) ,
    .IN ( masks_hold_reg_0_9 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_9 ) ,
    .IN ( masks_hold_reg_0_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_7 ) ,
    .IN ( masks_hold_reg_0_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_6 ) ,
    .IN ( masks_hold_reg_0_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_5 ) ,
    .IN ( masks_hold_reg_0_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_32 ) ,
    .IN ( n79 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_56 ) ,
    .IN ( masks_hold_reg_4_3 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_59 ) ,
    .IN ( masks_hold_reg_4_0 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_58 ) ,
    .IN ( masks_hold_reg_4_1 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_57 ) ,
    .IN ( masks_hold_reg_4_2 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_53 ) ,
    .IN ( masks_hold_reg_4_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_52 ) ,
    .IN ( masks_hold_reg_4_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_51 ) ,
    .IN ( masks_hold_reg_4_8 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_41 ) ,
    .IN ( masks_hold_reg_4_10 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_55 ) ,
    .IN ( masks_hold_reg_4_4 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_54 ) ,
    .IN ( masks_hold_reg_4_5 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_3 ) ,
    .IN ( masks_hold_reg_0_6 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_2 ) ,
    .IN ( masks_hold_reg_0_7 ) ) ;
buf ( 
    .O1 ( config1_xor_encoded_masks_4 ) ,
    .IN ( masks_hold_reg_0_5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_68 ) ,
    .I0 ( masks_hold_reg_4_1 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_69 ) ,
    .I0 ( masks_hold_reg_4_0 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_64 ) ,
    .I0 ( masks_hold_reg_4_5 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_67 ) ,
    .I0 ( masks_hold_reg_4_2 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_62 ) ,
    .I0 ( masks_hold_reg_4_7 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_63 ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_20 ) ,
    .I0 ( masks_hold_reg_0_1 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_19 ) ,
    .I0 ( masks_hold_reg_0_2 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n8 ) ,
    .I0 ( masks_hold_reg_8_10 ) ,
    .I1 ( masks_hold_reg_7_9 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_103 ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_102 ) ,
    .I0 ( masks_hold_reg_8_9 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_148 ) ,
    .I0 ( masks_hold_reg_12_5 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_46 ) ,
    .I0 ( masks_hold_reg_2_2 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_149 ) ,
    .I0 ( masks_hold_reg_12_4 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_66 ) ,
    .I0 ( masks_hold_reg_4_3 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_47 ) ,
    .I0 ( masks_hold_reg_2_1 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_146 ) ,
    .I0 ( masks_hold_reg_12_7 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_48 ) ,
    .I0 ( masks_hold_reg_2_0 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_147 ) ,
    .I0 ( masks_hold_reg_12_6 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n2 ) ,
    .I0 ( masks_hold_reg_4_8 ) ,
    .I1 ( n92 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_49 ) ,
    .I0 ( masks_hold_reg_3_10 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_28 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( plugin_xor_decoder.n4 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_29 ) ,
    .I0 ( masks_hold_reg_0_3 ) ,
    .I1 ( plugin_xor_decoder.n4 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_85 ) ,
    .I0 ( masks_hold_reg_6_5 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_86 ) ,
    .I0 ( masks_hold_reg_6_4 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_83 ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_84 ) ,
    .I0 ( masks_hold_reg_6_6 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_89 ) ,
    .I0 ( masks_hold_reg_6_1 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_87 ) ,
    .I0 ( masks_hold_reg_6_3 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_88 ) ,
    .I0 ( masks_hold_reg_6_2 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n1 ) ,
    .I0 ( masks_hold_reg_6_9 ) ,
    .I1 ( masks_hold_reg_6_10 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_82 ) ,
    .I0 ( masks_hold_reg_6_8 ) ,
    .I1 ( plugin_xor_decoder.n1 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_145 ) ,
    .I0 ( masks_hold_reg_12_8 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_144 ) ,
    .I0 ( masks_hold_reg_12_9 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n7 ) ,
    .I0 ( masks_hold_reg_9_9 ) ,
    .I1 ( masks_hold_reg_9_10 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_22 ) ,
    .I0 ( masks_hold_reg_1_10 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_143 ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_122 ) ,
    .I0 ( masks_hold_reg_10_10 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_21 ) ,
    .I0 ( masks_hold_reg_0_0 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_142 ) ,
    .I0 ( masks_hold_reg_11_9 ) ,
    .I1 ( plugin_xor_decoder.n6 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_123 ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_24 ) ,
    .I0 ( masks_hold_reg_2_10 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n6 ) ,
    .I0 ( masks_hold_reg_11_10 ) ,
    .I1 ( masks_hold_reg_10_0 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_124 ) ,
    .I0 ( masks_hold_reg_10_8 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_23 ) ,
    .I0 ( masks_hold_reg_1_9 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_129 ) ,
    .I0 ( masks_hold_reg_10_3 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_106 ) ,
    .I0 ( masks_hold_reg_8_5 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n4 ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_128 ) ,
    .I0 ( masks_hold_reg_10_4 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_107 ) ,
    .I0 ( masks_hold_reg_8_4 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_25 ) ,
    .I0 ( masks_hold_reg_2_9 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_127 ) ,
    .I0 ( masks_hold_reg_10_5 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_108 ) ,
    .I0 ( masks_hold_reg_8_3 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_27 ) ,
    .I0 ( masks_hold_reg_0_5 ) ,
    .I1 ( plugin_xor_decoder.n4 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_126 ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_109 ) ,
    .I0 ( masks_hold_reg_8_2 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_26 ) ,
    .I0 ( masks_hold_reg_0_6 ) ,
    .I1 ( plugin_xor_decoder.n4 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_125 ) ,
    .I0 ( masks_hold_reg_10_7 ) ,
    .I1 ( plugin_xor_decoder.n7 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_104 ) ,
    .I0 ( masks_hold_reg_8_7 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_105 ) ,
    .I0 ( masks_hold_reg_8_6 ) ,
    .I1 ( plugin_xor_decoder.n8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_17 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_65 ) ,
    .I0 ( masks_hold_reg_4_4 ) ,
    .I1 ( plugin_xor_decoder.n2 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_18 ) ,
    .I0 ( masks_hold_reg_0_3 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n3 ) ,
    .I0 ( masks_hold_reg_2_7 ) ,
    .I1 ( masks_hold_reg_2_8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_15 ) ,
    .I0 ( masks_hold_reg_0_6 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_42 ) ,
    .I0 ( n79 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_16 ) ,
    .I0 ( masks_hold_reg_0_5 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_43 ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( plugin_xor_decoder.n5 ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_44 ) ,
    .I0 ( masks_hold_reg_2_4 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_14 ) ,
    .I0 ( masks_hold_reg_0_7 ) ,
    .I1 ( plugin_xor_decoder.n5 ) ) ;
xor ( 
    .Z ( config1_xor_encoded_masks_45 ) ,
    .I0 ( masks_hold_reg_2_3 ) ,
    .I1 ( plugin_xor_decoder.n3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U606.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_350 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U606.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_317 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.decoder.n61 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U666.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_30 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U666.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_40 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n68 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U527.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_402 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U527.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_374 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n175 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U983.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_103 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U983.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U693.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_293 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U693.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n56 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n61 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.n360 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_312 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n125 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U516.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_410 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U516.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U524.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_405 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U524.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_549 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n29 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n178 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_515 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n139 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n180 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U402.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_492 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U402.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U456.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_451 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U456.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_445 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n164 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U932.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_133 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U932.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n29 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U944.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_126 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U944.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n130 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_512 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n83 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_308 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n180 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_490 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n150 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_450 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n34 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U465.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_446 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U465.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n101 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_560 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n128 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_554 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n128 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U945.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_125 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U945.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_313 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n40 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n123 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_64 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n26 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n14 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_677 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n78 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n92 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_613 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.n108 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U728.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_270 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.decoder.U728.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U984.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_102 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U984.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U698.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.n913 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_28 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U698.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U191.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_654 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.decoder.U191.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_681 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n77 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_676 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n79 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_583 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n92 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U719.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_277 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U719.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U729.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_26 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U729.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U511.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_414 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U511.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U985.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_101 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U985.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U699.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_289 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U699.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_352 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n180 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U190.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_655 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U190.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_682 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n76 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n77 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.n813 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_278 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n74 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U510.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_415 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U510.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n33 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U986.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_100 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.U986.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U602.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_353 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U602.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n20 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_652 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n93 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_584 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n77 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_60 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n110 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U513.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_412 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U513.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U523.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_406 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U523.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U577.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_370 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U577.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_0 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n132 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U601.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_354 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U601.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_314 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n130 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_653 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n92 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n104 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U108.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_724 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U108.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_673 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n82 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U280.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_585 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U280.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_616 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n9 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n52 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_232 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n159 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U512.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_413 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U512.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U520.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_408 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U520.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U576.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_371 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U576.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n136 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U600.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_355 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U600.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U948.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_123 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U948.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U654.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_316 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U654.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_310 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n104 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_723 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n54 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U169.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_672 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U169.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n9 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U778.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_233 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U778.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n93 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.n461 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_407 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n33 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U575.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_372 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U575.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_104 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n85 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_34 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.decoder.n181 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U949.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_122 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U949.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_315 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n20 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U667.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_309 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U667.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_411 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n93 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_403 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n131 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U574.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_373 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U574.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n85 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n59 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_510 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n108 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_425 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n88 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_488 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.n152 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n114 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n166 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_200 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n192 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_778 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n24 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U10.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_91 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U10.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_79 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n16 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_509 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n115 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n88 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_209 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n132 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n46 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_227 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.decoder.n168 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_779 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n23 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_90 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.n5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_7 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n15 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_50 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n140 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U496.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_424 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U496.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U115.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_718 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U115.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U816.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_208 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U816.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_640 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n48 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_201 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n46 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U872.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_173 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U872.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n168 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_776 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n25 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U731.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_268 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U731.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_8 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U746.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.n381 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_257 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U746.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U22.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_80 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U22.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_423 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n94 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U114.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_719 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U114.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_709 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n60 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U817.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_207 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U817.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_641 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.n97 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n169 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_607 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_172 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n188 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U46.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_777 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U46.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U730.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.n331 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_269 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U730.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_89 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_256 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n190 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_81 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n14 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_548 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n32 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_716 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n56 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_375 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n174 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n170 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_351 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n56 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_318 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n106 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n40 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U519.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_409 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U519.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_404 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n168 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n82 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_294 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.n59 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U939.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_12 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U939.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n106 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_311 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n185 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n94 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n68 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_376 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.n82 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U696.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_291 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U696.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n120 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n125 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U499.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_422 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U499.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U697.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_290 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U697.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_130 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n120 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n58 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_401 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n51 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n132 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_292 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n182 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U317.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_557 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U317.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n100 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_349 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n58 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U940.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_129 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U940.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_493 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n149 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n51 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n182 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.n331 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_558 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n98 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_131 ) ,
    .I0 ( constant_shift_controller_i.n320 ) ,
    .I1 ( constant_shift_controller_i.decoder.n100 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_550 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n54 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U941.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_128 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.decoder.U941.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U400.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_494 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U400.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U454.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_453 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U454.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_559 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n126 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n118 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U325.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_54 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U325.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_127 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n178 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U371.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_514 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U371.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_491 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n60 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U455.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_452 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U455.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_444 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n137 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U314.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_55 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U314.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_132 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n118 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_671 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n15 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U469.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_443 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.U469.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_574 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n121 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_20 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.n166 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U202.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_645 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U202.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n25 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_603 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n114 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U877.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_16 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U877.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U262.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_59 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.U262.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n110 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U734.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_265 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U734.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_259 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n99 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U113.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_71 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U113.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n5 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_666 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n86 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n137 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U297.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_573 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U297.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_646 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n96 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_204 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n25 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U257.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_602 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U257.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n188 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_598 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.decoder.n115 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U783.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_230 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U783.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U737.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_262 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U737.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U18.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_84 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U18.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n4 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_720 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.decoder.n55 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_713 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n58 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_667 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n85 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_575 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n80 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U200.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_647 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U200.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U254.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_605 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.decoder.U254.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U875.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_171 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U875.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n89 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n159 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U736.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_263 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U736.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_83 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.decoder.n12 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_25 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n175 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U588.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_363 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.U588.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_712 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n59 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U175.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_668 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U175.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n80 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U255.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.n913 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_604 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U255.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U267.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_596 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U267.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_231 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n110 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_260 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_362 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n37 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U174.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_669 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U174.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U372.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_513 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U372.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U490.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_428 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.U490.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n60 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U450.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_456 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U450.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n73 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U818.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_206 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U818.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_169 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n141 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U41.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_781 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U41.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_88 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n8 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_36 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n101 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U311.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_561 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U311.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_134 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n128 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U321.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.n813 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_553 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U321.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_124 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n157 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_511 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n91 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U491.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_427 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U491.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U407.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_489 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U407.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_455 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n162 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_447 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n73 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U819.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.n461 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_205 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U819.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n141 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U40.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_782 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U40.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_87 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n9 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_793 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n17 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_562 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n125 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_552 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n129 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n157 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n83 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_426 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n151 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_48 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n151 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_454 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n160 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U462.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_448 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.decoder.U462.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U43.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_77 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U43.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_86 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n10 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U26.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_794 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U26.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U323.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_551 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U323.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n108 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n151 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U409.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_487 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U409.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n160 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_449 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n163 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U829.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U829.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U42.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_780 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U42.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_85 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n11 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U25.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_795 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U25.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_117 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n63 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_337 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n131 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n164 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U118.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_715 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U118.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_665 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n50 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_97 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_400 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n148 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n156 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U616.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_342 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.U616.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n172 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U622.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_338 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U622.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_303 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n186 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_639 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n99 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U7.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_94 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U7.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U748.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_255 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U748.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_397 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n140 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_391 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n100 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U617.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_341 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U617.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U625.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.n381 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_336 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U625.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_302 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n187 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_707 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.n62 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_63 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n98 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_95 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U749.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_254 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U749.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U580.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_369 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U580.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U536.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_398 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U536.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_395 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n109 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U908.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_14 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U908.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U614.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_344 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.decoder.U614.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n131 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U968.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_111 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U968.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_307 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n144 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_706 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.n63 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U1.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_9 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U1.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U581.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_368 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U581.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U535.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_399 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U535.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n109 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U909.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_149 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U909.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U615.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_343 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U615.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n30 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_110 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n62 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n144 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_367 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n176 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n21 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_394 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n87 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_335 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n30 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U672.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_306 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U672.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_98 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_366 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n43 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_708 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n61 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n34 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_66 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n84 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n187 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U205.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_642 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U205.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_202 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n169 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U253.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_606 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U253.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U870.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_175 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.U870.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U261.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_5 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U261.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_774 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n27 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_266 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n124 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n99 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_82 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n13 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_555 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n17 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n32 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U116.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_717 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U116.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U124.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_710 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U124.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_44 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n114 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_670 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n83 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U298.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_572 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U298.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U811.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_211 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U811.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_643 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n51 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n186 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_609 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n111 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U871.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_174 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U871.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U260.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_600 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U260.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_775 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.n26 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U732.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_267 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U732.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U745.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_258 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U745.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_556 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n127 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U111.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_721 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U111.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U125.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_70 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U125.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n15 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_571 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n122 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U812.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_210 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U812.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U203.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_644 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U203.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_203 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n186 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_608 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n112 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U876.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_170 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U876.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_599 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n89 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_264 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n168 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n175 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.n401 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U110.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_722 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U110.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_711 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n54 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_120 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n189 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_486 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n8 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n76 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n72 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n140 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n91 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_543 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n125 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U950.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_121 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U950.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n152 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n8 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.n913 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n53 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n22 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_364 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n177 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U907.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_150 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U907.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_544 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n131 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_11 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n165 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U342.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_537 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U342.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U963.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_115 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U963.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U412.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_485 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U412.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_477 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.n53 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_439 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n26 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_164 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n22 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U548.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_390 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U548.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U900.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.n441 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_154 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U900.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_541 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n133 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n189 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_536 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n136 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n63 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_301 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n57 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_484 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n153 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U421.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_478 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U421.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n26 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.n401 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_167 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n192 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_188 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n191 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U9.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_92 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U9.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U549.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_38 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U549.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_502 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n143 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_153 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n155 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_542 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n132 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_119 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n117 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_539 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n135 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_116 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.n152 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n57 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U414.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_483 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U414.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_479 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n118 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_440 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n165 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U880.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_168 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U880.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U848.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_189 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U848.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U8.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_93 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U8.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_501 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.decoder.n144 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n155 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_546 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.decoder.n44 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n165 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U341.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_538 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U341.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n177 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U415.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_482 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U415.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U427.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_474 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U427.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U475.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_43 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U475.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_166 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n76 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U50.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_773 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U50.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U386.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_504 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U386.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_577 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n81 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_597 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n67 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U786.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_229 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U786.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U738.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_261 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U738.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_791 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.n19 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U612.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_346 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U612.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U293.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_576 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U293.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U269.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_594 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U269.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U787.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_228 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U787.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_792 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.n18 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_39 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n21 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U613.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_345 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U613.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U621.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_339 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U621.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_579 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n120 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_601 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n71 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U268.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_595 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U268.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_22 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n112 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_3 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n169 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U544.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_393 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U544.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U610.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_348 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U610.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_33 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n182 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_304 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n164 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_714 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n57 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_664 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n87 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U291.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_578 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U291.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n71 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n112 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_96 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n148 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_392 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n156 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U611.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_347 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U611.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n192 ) ,
    .I0 ( constant_shift_controller_i.n320 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_772 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U63.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_763 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U63.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_786 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.decoder.n11 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U387.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_503 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U387.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_545 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n120 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n117 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U347.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_532 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U347.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U964.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_114 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U964.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U417.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_480 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U417.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_475 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n96 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n146 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n7 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_764 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n30 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_785 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n21 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n66 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n44 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U344.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_535 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U344.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_113 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n177 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_47 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.decoder.n6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U424.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_476 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U424.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_442 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n135 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U838.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_195 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U838.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_73 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n46 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_771 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U61.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_765 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U61.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U34.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_788 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U34.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U385.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.n1013 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_505 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U385.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_534 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n137 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n6 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n135 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U839.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_194 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U839.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U88.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_740 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U88.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n3 ) ,
    .I0 ( constant_shift_controller_i.n320 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U60.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_766 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U60.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_787 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n20 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_507 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n142 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n81 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.n331 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U799.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_219 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U799.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_770 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n28 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U67.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_75 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U67.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_789 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_506 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n66 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U429.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.n381 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_472 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U429.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U889.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_162 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U889.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U216.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_632 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U216.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U837.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_196 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U837.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n190 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U798.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_21 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U798.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U56.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_76 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.decoder.U56.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U702.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_287 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U702.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_760 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n32 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U757.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_248 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U757.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n2 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n115 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_531 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_6 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n66 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_473 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n155 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U888.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_163 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U888.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_631 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n12 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U834.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_198 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U834.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U225.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_627 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U225.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_193 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n190 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_743 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n43 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_769 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n29 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_286 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n67 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U65.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_761 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.U65.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U756.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_249 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U756.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U30.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_790 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U30.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n42 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.n461 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_508 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n141 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_53 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n134 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U349.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_530 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U349.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_656 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n11 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U136.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_700 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U136.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_698 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n69 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_634 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n102 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_197 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n81 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U224.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_628 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U224.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n167 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U270.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_593 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U270.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n87 ) ,
    .I0 ( constant_shift_controller_i.n320 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U629.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_333 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U629.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U673.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_305 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U673.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U2.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_99 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U2.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n43 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n149 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_340 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n54 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_334 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n169 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U885.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_165 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.decoder.U885.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_365 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n72 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_396 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n170 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_151 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n91 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n11 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n41 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .I1 ( constant_shift_controller_i.n441 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_697 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n70 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U215.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_633 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.decoder.U215.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_199 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n121 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_625 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n86 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_192 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n167 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U271.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_592 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U271.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_741 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n45 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U59.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_767 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U59.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n162 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n111 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.n401 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U766.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_241 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U766.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_701 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n41 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U142.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_696 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U142.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_636 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n100 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n121 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_626 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.decoder.n104 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_190 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n126 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_591 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.n116 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_742 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n44 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n183 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_250 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n111 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U767.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_240 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U767.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U133.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_702 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U133.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_695 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n66 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U478.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_438 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U478.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_635 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n101 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_19 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n171 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_62 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.n35 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U844.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_191 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U844.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U273.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_590 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U273.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n122 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U81.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_747 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U81.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_284 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n158 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_758 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n34 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U752.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_251 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U752.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U760.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_245 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U760.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U184.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_65 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U184.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_703 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n65 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_694 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.decoder.n71 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U479.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_437 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U479.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U210.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_638 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U210.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n171 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n10 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U847.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_18 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U847.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U274.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_58 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U274.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_224 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n122 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_748 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n39 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n67 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_759 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n33 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U751.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_252 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U751.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_244 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n161 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_659 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n90 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_704 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n64 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_693 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n72 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U211.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.n1013 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_637 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.U211.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_629 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n103 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n126 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.n391 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U275.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_589 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U275.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U791.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_225 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U791.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_745 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n41 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_285 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n183 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U750.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_253 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U750.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n161 ) ,
    .I0 ( constant_shift_controller_i.n320 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U599.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_356 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U599.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_658 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n91 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U130.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_705 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U130.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_692 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n73 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n35 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .I1 ( constant_shift_controller_i.n391 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U276.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_588 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U276.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U790.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_226 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.U790.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_746 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n40 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_243 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n42 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_357 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n179 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U187.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_657 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U187.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_691 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n74 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_587 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n117 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U797.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_220 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U797.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U38.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_784 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U38.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_295 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n170 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U180.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_663 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U180.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U148.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_690 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U148.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_586 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n27 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U796.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.n1013 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_221 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U796.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_152 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n149 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_547 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n130 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_118 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n172 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U346.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_533 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U346.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U967.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_112 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U967.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_481 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n154 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n96 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_441 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n146 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U869.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_176 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U869.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_755 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.n36 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n64 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U396.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_497 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U396.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n158 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_783 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n22 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_421 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n107 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U688.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_296 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U688.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U630.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_332 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U630.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U181.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_662 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U181.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U149.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_68 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U149.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n27 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U795.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_222 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U795.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U709.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_283 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U709.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n107 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_386 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n172 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_331 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n17 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_31 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n163 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_661 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.decoder.n88 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U794.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_223 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.U794.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_420 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n167 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n65 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n23 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n17 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.n461 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_320 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n183 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_660 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n89 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U229.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_624 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U229.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_23 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n49 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_41 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n139 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U557.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_384 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.U557.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U567.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_378 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U567.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U633.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.n1013 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_330 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U633.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U645.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_321 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U645.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n12 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n86 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.n331 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U759.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_246 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U759.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n49 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n139 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_385 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n173 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U564.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_37 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U564.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U634.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_32 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U634.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n47 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_699 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n68 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_630 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n10 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U758.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_247 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U758.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_361 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n134 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_419 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n56 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_388 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n116 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_379 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n23 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U683.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_29 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U683.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_141 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n185 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_329 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n119 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_105 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n136 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_322 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n47 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_69 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n67 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n37 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U506.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_418 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U506.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_389 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n171 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_380 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.decoder.n150 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_2 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n188 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U918.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.n381 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_142 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U918.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n119 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n75 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.n451 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U642.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_323 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U642.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U593.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_360 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U593.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_417 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n147 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_387 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n65 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n150 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n129 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U637.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_328 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U637.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U641.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_324 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U641.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n134 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n147 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n116 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U560.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_382 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U560.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_300 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.n129 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n74 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.n913 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U638.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_327 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U638.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U640.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_325 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U640.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n79 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_359 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n18 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U509.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_416 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U509.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U561.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_381 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U561.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U687.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_297 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U687.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U915.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_144 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U915.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_744 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n42 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U58.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_768 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U58.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_288 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n162 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_762 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n31 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_24 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n191 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U31.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_78 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U31.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U765.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_242 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U765.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U338.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_540 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U338.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_752 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n37 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n36 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n55 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_648 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n69 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U106.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.n351 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_726 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.U106.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U150.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_689 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U150.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_457 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.decoder.n161 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U162.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_679 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U162.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_217 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n133 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U236.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_618 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U236.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U853.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_185 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U853.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_614 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n13 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_180 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n102 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_733 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n19 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U710.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_282 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U710.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U722.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_275 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U722.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U777.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_234 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U777.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_563 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n45 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U929.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_135 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U929.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U639.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_326 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U639.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_429 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n79 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_158 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n103 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_35 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n178 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n145 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.n441 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U914.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_145 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U914.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U926.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_137 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.U926.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n103 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U597.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_358 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U597.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_298 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.n145 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n179 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.n461 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_565 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n124 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_136 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n74 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n173 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_46 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n156 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U896.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_157 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U896.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n18 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U684.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.decoder.U684.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_143 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n179 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U307.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_564 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U307.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U924.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_139 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U924.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_528 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n30 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_109 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n173 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_469 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n138 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U445.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_460 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.U445.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_156 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n124 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n39 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n16 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_567 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n123 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U925.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_138 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U925.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U352.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_529 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.decoder.U352.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U971.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_10 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U971.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_522 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n38 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_471 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n139 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n95 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U890.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n431 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_161 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U890.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n105 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_383 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n39 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_495 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n148 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_148 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n16 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_566 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n36 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_13 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n24 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n62 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n38 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U431.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_470 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U431.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U447.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_459 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U447.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U891.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_160 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U891.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_181 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.decoder.n174 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n48 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U913.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_146 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U913.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U302.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_569 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U302.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n113 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.n391 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_52 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n24 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_106 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n75 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_319 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n184 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U362.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_521 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.decoder.U362.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n98 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_45 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n160 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U892.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_15 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U892.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_377 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n64 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_496 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n48 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U912.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_147 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.U912.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U303.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_568 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U303.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n185 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U357.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_524 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U357.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n70 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n163 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_520 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n51 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U481.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_435 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U481.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_467 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n157 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U441.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_463 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U441.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U893.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_159 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U893.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_212 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.decoder.n187 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_729 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n31 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_685 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n75 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_675 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n80 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_581 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n119 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U232.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_621 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U232.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_182 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n105 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U246.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_611 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U246.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_178 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n142 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U92.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_737 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U92.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_27 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n176 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n154 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_237 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n55 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_649 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n95 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n31 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U157.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_683 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U157.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_674 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n81 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_582 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n118 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U233.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_620 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U233.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_612 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n109 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U864.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_179 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U864.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U93.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_736 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U93.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_271 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.decoder.n169 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U300.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_570 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U300.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U921.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_140 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U921.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U356.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_525 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U356.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_107 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n70 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_51 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n138 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_436 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.decoder.n166 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n138 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_464 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n159 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U808.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_213 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U808.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n181 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.n813 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U73.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_754 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U73.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_498 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n147 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U301.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n461 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_56 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U301.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U355.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_526 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U355.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U974.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .I1 ( constant_shift_controller_i.n331 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_108 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U974.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_519 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.n119 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U483.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_433 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U483.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_468 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n98 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_461 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.n95 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U98.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_732 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U98.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U70.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.n410 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_757 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U70.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_499 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n146 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U354.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_527 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U354.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U366.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_518 ) ,
    .I0 ( constant_shift_controller_i.n410 ) ,
    .I1 ( constant_shift_controller_i.decoder.U366.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_434 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n91 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U442.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_462 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U442.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_731 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n51 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_756 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n35 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n28 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_517 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.decoder.n78 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_431 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n141 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_215 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n84 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_751 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n38 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_49 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n28 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n78 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U484.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_432 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U484.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U438.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_466 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U438.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n124 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n143 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n191 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n184 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U77.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_750 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U77.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_4 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n87 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n50 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U369.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n913 ) ,
    .I1 ( constant_shift_controller_i.n320 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_516 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U369.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U487.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_42 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U487.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U104.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_728 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U104.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_465 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n158 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U899.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_155 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U899.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U807.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.n913 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_214 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U807.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_61 ) ,
    .I0 ( constant_shift_controller_i.n351 ) ,
    .I1 ( constant_shift_controller_i.decoder.n107 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U851.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_187 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U851.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U863.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_17 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U863.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_735 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n49 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_280 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n184 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U74.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.n441 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_753 ) ,
    .I0 ( constant_shift_controller_i.n391 ) ,
    .I1 ( constant_shift_controller_i.decoder.U74.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_276 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.decoder.n36 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U775.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_236 ) ,
    .I0 ( constant_shift_controller_i.n371 ) ,
    .I1 ( constant_shift_controller_i.decoder.U775.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_500 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n145 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_523 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.n50 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n69 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U486.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_430 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U486.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_727 ) ,
    .I0 ( constant_shift_controller_i.n331 ) ,
    .I1 ( constant_shift_controller_i.decoder.n53 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U151.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_688 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U151.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n84 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U235.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_619 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U235.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U852.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.n371 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_186 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U852.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n13 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n102 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_734 ) ,
    .I0 ( constant_shift_controller_i.n381 ) ,
    .I1 ( constant_shift_controller_i.decoder.n50 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U711.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_281 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.U711.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U107.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_725 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U107.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U153.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_686 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U153.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U448.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_458 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U448.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U163.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_678 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U163.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U289.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_57 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U289.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U800.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n451 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_218 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.U800.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U237.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_617 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U237.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_184 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n127 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n97 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n174 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n19 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n153 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_274 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n189 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U776.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n401 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_235 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U776.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n45 ) ,
    .I0 ( constant_shift_controller_i.n421 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_730 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n52 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U152.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n340 ) ,
    .I1 ( constant_shift_controller_i.n421 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_687 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.U152.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U160.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n1113 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_4 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_680 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U160.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n90 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_216 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n143 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_623 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n105 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n127 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_615 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n97 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_177 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n181 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_739 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.n47 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_279 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n153 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U78.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_74 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.U78.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_273 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.n46 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_238 ) ,
    .I0 ( constant_shift_controller_i.n813 ) ,
    .I1 ( constant_shift_controller_i.decoder.n123 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_650 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .I1 ( constant_shift_controller_i.decoder.n94 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U101.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_72 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .I1 ( constant_shift_controller_i.decoder.U101.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_684 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.n14 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U161.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .I1 ( constant_shift_controller_i.n340 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_67 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .I1 ( constant_shift_controller_i.decoder.U161.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_580 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .I1 ( constant_shift_controller_i.decoder.n90 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n133 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_622 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n106 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U856.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.n441 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_183 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U856.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_610 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .I1 ( constant_shift_controller_i.decoder.n52 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n142 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .I1 ( constant_shift_controller_i.n1113 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_738 ) ,
    .I0 ( constant_shift_controller_i.n1013 ) ,
    .I1 ( constant_shift_controller_i.decoder.n48 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.n176 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_0 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U79.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_749 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .I1 ( constant_shift_controller_i.decoder.U79.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_272 ) ,
    .I0 ( constant_shift_controller_i.n360 ) ,
    .I1 ( constant_shift_controller_i.decoder.n154 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U770.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_239 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.decoder.U770.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.decoder.U194.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ) ;
xor ( 
    .Z ( constant_shift_controller_i.bias_inputs_651 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .I1 ( constant_shift_controller_i.decoder.U194.SYNTEST_VL_xor_28002_299 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n1113 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n1013 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n913 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n813 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_0 ) ) ;
and ( 
    .Z ( edt_scan_in_759 ) ,
    .I0 ( edt_decompressor_out_759 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_759 ) ) ;
and ( 
    .Z ( edt_scan_in_530 ) ,
    .I0 ( edt_decompressor_out_530 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_530 ) ) ;
and ( 
    .Z ( edt_scan_in_242 ) ,
    .I0 ( edt_decompressor_out_242 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_242 ) ) ;
and ( 
    .Z ( edt_scan_in_197 ) ,
    .I0 ( edt_decompressor_out_197 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_197 ) ) ;
and ( 
    .Z ( edt_scan_in_335 ) ,
    .I0 ( edt_decompressor_out_335 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_335 ) ) ;
and ( 
    .Z ( edt_scan_in_38 ) ,
    .I0 ( edt_decompressor_out_38 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_38 ) ) ;
and ( 
    .Z ( edt_scan_in_263 ) ,
    .I0 ( edt_decompressor_out_263 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_263 ) ) ;
and ( 
    .Z ( edt_scan_in_257 ) ,
    .I0 ( edt_decompressor_out_257 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_257 ) ) ;
and ( 
    .Z ( edt_scan_in_205 ) ,
    .I0 ( edt_decompressor_out_205 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_205 ) ) ;
and ( 
    .Z ( edt_scan_in_198 ) ,
    .I0 ( edt_decompressor_out_198 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_198 ) ) ;
and ( 
    .Z ( edt_scan_in_606 ) ,
    .I0 ( edt_decompressor_out_606 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_606 ) ) ;
and ( 
    .Z ( edt_scan_in_83 ) ,
    .I0 ( edt_decompressor_out_83 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_83 ) ) ;
and ( 
    .Z ( edt_scan_in_298 ) ,
    .I0 ( edt_decompressor_out_298 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_298 ) ) ;
and ( 
    .Z ( edt_scan_in_265 ) ,
    .I0 ( edt_decompressor_out_265 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_265 ) ) ;
and ( 
    .Z ( edt_scan_in_272 ) ,
    .I0 ( edt_decompressor_out_272 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_272 ) ) ;
and ( 
    .Z ( edt_scan_in_201 ) ,
    .I0 ( edt_decompressor_out_201 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_201 ) ) ;
and ( 
    .Z ( edt_scan_in_119 ) ,
    .I0 ( edt_decompressor_out_119 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_119 ) ) ;
and ( 
    .Z ( edt_scan_in_81 ) ,
    .I0 ( edt_decompressor_out_81 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_81 ) ) ;
and ( 
    .Z ( edt_scan_in_399 ) ,
    .I0 ( edt_decompressor_out_399 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_399 ) ) ;
and ( 
    .Z ( edt_scan_in_111 ) ,
    .I0 ( edt_decompressor_out_111 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_111 ) ) ;
and ( 
    .Z ( edt_scan_in_154 ) ,
    .I0 ( edt_decompressor_out_154 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_154 ) ) ;
and ( 
    .Z ( edt_scan_in_126 ) ,
    .I0 ( edt_decompressor_out_126 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_126 ) ) ;
and ( 
    .Z ( edt_scan_in_244 ) ,
    .I0 ( edt_decompressor_out_244 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_244 ) ) ;
and ( 
    .Z ( edt_scan_in_151 ) ,
    .I0 ( edt_decompressor_out_151 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_151 ) ) ;
and ( 
    .Z ( edt_scan_in_438 ) ,
    .I0 ( edt_decompressor_out_438 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_438 ) ) ;
and ( 
    .Z ( edt_scan_in_170 ) ,
    .I0 ( edt_decompressor_out_170 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_170 ) ) ;
and ( 
    .Z ( edt_scan_in_749 ) ,
    .I0 ( edt_decompressor_out_749 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_749 ) ) ;
and ( 
    .Z ( edt_scan_in_204 ) ,
    .I0 ( edt_decompressor_out_204 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_204 ) ) ;
and ( 
    .Z ( edt_scan_in_294 ) ,
    .I0 ( edt_decompressor_out_294 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_294 ) ) ;
and ( 
    .Z ( edt_scan_in_196 ) ,
    .I0 ( edt_decompressor_out_196 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_196 ) ) ;
and ( 
    .Z ( edt_scan_in_49 ) ,
    .I0 ( edt_decompressor_out_49 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_49 ) ) ;
and ( 
    .Z ( edt_scan_in_381 ) ,
    .I0 ( edt_decompressor_out_381 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_381 ) ) ;
and ( 
    .Z ( edt_scan_in_523 ) ,
    .I0 ( edt_decompressor_out_523 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_523 ) ) ;
and ( 
    .Z ( edt_scan_in_619 ) ,
    .I0 ( edt_decompressor_out_619 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_619 ) ) ;
and ( 
    .Z ( edt_scan_in_339 ) ,
    .I0 ( edt_decompressor_out_339 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_339 ) ) ;
and ( 
    .Z ( edt_scan_in_481 ) ,
    .I0 ( edt_decompressor_out_481 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_481 ) ) ;
and ( 
    .Z ( edt_scan_in_136 ) ,
    .I0 ( edt_decompressor_out_136 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_136 ) ) ;
and ( 
    .Z ( edt_scan_in_60 ) ,
    .I0 ( edt_decompressor_out_60 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_60 ) ) ;
and ( 
    .Z ( edt_scan_in_618 ) ,
    .I0 ( edt_decompressor_out_618 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_618 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n812 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n912 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n1012 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n1112 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n127 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n250 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n290 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n300 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_3 ) ) ;
and ( 
    .Z ( edt_scan_in_300 ) ,
    .I0 ( edt_decompressor_out_300 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_300 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n650 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N80 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n3 ) ) ;
and ( 
    .Z ( edt_scan_in_301 ) ,
    .I0 ( edt_decompressor_out_301 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_301 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N71 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n650 ) ) ;
and ( 
    .Z ( edt_scan_in_302 ) ,
    .I0 ( edt_decompressor_out_302 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_302 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N91 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n170 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N88 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n370 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N72 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n6 ) ) ;
and ( 
    .Z ( edt_scan_in_268 ) ,
    .I0 ( edt_decompressor_out_268 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_268 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N46 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n260 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n300 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_2 ) ) ;
and ( 
    .Z ( edt_scan_in_267 ) ,
    .I0 ( edt_decompressor_out_267 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_267 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N106 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1400 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_3 ) ) ;
and ( 
    .Z ( edt_scan_in_266 ) ,
    .I0 ( edt_decompressor_out_266 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_266 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N10 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1420 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n471 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1420 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_1 ) ) ;
and ( 
    .Z ( edt_scan_in_273 ) ,
    .I0 ( edt_decompressor_out_273 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_273 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N95 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n450 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N64 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n810 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n450 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N96 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n350 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N238 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_7 ) ) ;
and ( 
    .Z ( edt_scan_in_579 ) ,
    .I0 ( edt_decompressor_out_579 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_579 ) ) ;
and ( 
    .Z ( edt_scan_in_271 ) ,
    .I0 ( edt_decompressor_out_271 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_271 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N94 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n460 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N36 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_4 ) ) ;
and ( 
    .Z ( edt_scan_in_580 ) ,
    .I0 ( edt_decompressor_out_580 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_580 ) ) ;
and ( 
    .Z ( edt_scan_in_269 ) ,
    .I0 ( edt_decompressor_out_269 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_269 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n460 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N37 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_5.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n311 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_13_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_13_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_13_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_13_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_13_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N93 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n470 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N38 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_6.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n470 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N39 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_575 ) ,
    .I0 ( edt_decompressor_out_575 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_575 ) ) ;
and ( 
    .Z ( edt_scan_in_275 ) ,
    .I0 ( edt_decompressor_out_275 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_275 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N92 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n480 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N32 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_576 ) ,
    .I0 ( edt_decompressor_out_576 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_576 ) ) ;
and ( 
    .Z ( edt_scan_in_274 ) ,
    .I0 ( edt_decompressor_out_274 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_274 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n480 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N33 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_577 ) ,
    .I0 ( edt_decompressor_out_577 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_577 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N34 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_578 ) ,
    .I0 ( edt_decompressor_out_578 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_578 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N35 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_3_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_3_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_3_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_3_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_3_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_571 ) ,
    .I0 ( edt_decompressor_out_571 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_571 ) ) ;
and ( 
    .Z ( edt_scan_in_572 ) ,
    .I0 ( edt_decompressor_out_572 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_572 ) ) ;
and ( 
    .Z ( edt_scan_in_573 ) ,
    .I0 ( edt_decompressor_out_573 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_573 ) ) ;
and ( 
    .Z ( edt_scan_in_574 ) ,
    .I0 ( edt_decompressor_out_574 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_574 ) ) ;
and ( 
    .Z ( edt_scan_in_592 ) ,
    .I0 ( edt_decompressor_out_592 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_592 ) ) ;
and ( 
    .Z ( edt_scan_in_511 ) ,
    .I0 ( edt_decompressor_out_511 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_511 ) ) ;
and ( 
    .Z ( edt_scan_in_510 ) ,
    .I0 ( edt_decompressor_out_510 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_510 ) ) ;
and ( 
    .Z ( edt_scan_in_513 ) ,
    .I0 ( edt_decompressor_out_513 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_513 ) ) ;
and ( 
    .Z ( edt_scan_in_512 ) ,
    .I0 ( edt_decompressor_out_512 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_512 ) ) ;
and ( 
    .Z ( edt_scan_in_515 ) ,
    .I0 ( edt_decompressor_out_515 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_515 ) ) ;
and ( 
    .Z ( edt_scan_in_714 ) ,
    .I0 ( edt_decompressor_out_714 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_714 ) ) ;
and ( 
    .Z ( edt_scan_in_514 ) ,
    .I0 ( edt_decompressor_out_514 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_514 ) ) ;
and ( 
    .Z ( edt_scan_in_380 ) ,
    .I0 ( edt_decompressor_out_380 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_380 ) ) ;
and ( 
    .Z ( edt_scan_in_715 ) ,
    .I0 ( edt_decompressor_out_715 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_715 ) ) ;
and ( 
    .Z ( edt_scan_in_517 ) ,
    .I0 ( edt_decompressor_out_517 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_517 ) ) ;
and ( 
    .Z ( edt_scan_in_379 ) ,
    .I0 ( edt_decompressor_out_379 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_379 ) ) ;
and ( 
    .Z ( edt_scan_in_716 ) ,
    .I0 ( edt_decompressor_out_716 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_716 ) ) ;
and ( 
    .Z ( edt_scan_in_516 ) ,
    .I0 ( edt_decompressor_out_516 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_516 ) ) ;
and ( 
    .Z ( edt_scan_in_377 ) ,
    .I0 ( edt_decompressor_out_377 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_377 ) ) ;
and ( 
    .Z ( edt_scan_in_717 ) ,
    .I0 ( edt_decompressor_out_717 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_717 ) ) ;
and ( 
    .Z ( edt_scan_in_385 ) ,
    .I0 ( edt_decompressor_out_385 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_385 ) ) ;
and ( 
    .Z ( edt_scan_in_718 ) ,
    .I0 ( edt_decompressor_out_718 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_718 ) ) ;
and ( 
    .Z ( edt_scan_in_384 ) ,
    .I0 ( edt_decompressor_out_384 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_384 ) ) ;
and ( 
    .Z ( edt_scan_in_719 ) ,
    .I0 ( edt_decompressor_out_719 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_719 ) ) ;
and ( 
    .Z ( edt_scan_in_383 ) ,
    .I0 ( edt_decompressor_out_383 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_383 ) ) ;
and ( 
    .Z ( edt_scan_in_720 ) ,
    .I0 ( edt_decompressor_out_720 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_720 ) ) ;
and ( 
    .Z ( edt_scan_in_382 ) ,
    .I0 ( edt_decompressor_out_382 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_382 ) ) ;
and ( 
    .Z ( edt_scan_in_721 ) ,
    .I0 ( edt_decompressor_out_721 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_721 ) ) ;
and ( 
    .Z ( edt_scan_in_722 ) ,
    .I0 ( edt_decompressor_out_722 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_722 ) ) ;
and ( 
    .Z ( edt_scan_in_296 ) ,
    .I0 ( edt_decompressor_out_296 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_296 ) ) ;
and ( 
    .Z ( edt_scan_in_723 ) ,
    .I0 ( edt_decompressor_out_723 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_723 ) ) ;
and ( 
    .Z ( edt_scan_in_297 ) ,
    .I0 ( edt_decompressor_out_297 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_297 ) ) ;
and ( 
    .Z ( edt_scan_in_387 ) ,
    .I0 ( edt_decompressor_out_387 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_387 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n500 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_1 ) ) ;
and ( 
    .Z ( edt_scan_in_386 ) ,
    .I0 ( edt_decompressor_out_386 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_386 ) ) ;
and ( 
    .Z ( edt_scan_in_299 ) ,
    .I0 ( edt_decompressor_out_299 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_299 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N9 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n500 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N106 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_585 ) ,
    .I0 ( edt_decompressor_out_585 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_585 ) ) ;
and ( 
    .Z ( edt_scan_in_285 ) ,
    .I0 ( edt_decompressor_out_285 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N107 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_588 ) ,
    .I0 ( edt_decompressor_out_588 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_588 ) ) ;
and ( 
    .Z ( edt_scan_in_245 ) ,
    .I0 ( edt_decompressor_out_245 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_245 ) ) ;
and ( 
    .Z ( edt_scan_in_587 ) ,
    .I0 ( edt_decompressor_out_587 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_587 ) ) ;
and ( 
    .Z ( edt_scan_in_246 ) ,
    .I0 ( edt_decompressor_out_246 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_246 ) ) ;
and ( 
    .Z ( edt_scan_in_582 ) ,
    .I0 ( edt_decompressor_out_582 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_582 ) ) ;
and ( 
    .Z ( edt_scan_in_247 ) ,
    .I0 ( edt_decompressor_out_247 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_247 ) ) ;
and ( 
    .Z ( edt_scan_in_581 ) ,
    .I0 ( edt_decompressor_out_581 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_581 ) ) ;
and ( 
    .Z ( edt_scan_in_248 ) ,
    .I0 ( edt_decompressor_out_248 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_248 ) ) ;
and ( 
    .Z ( edt_scan_in_584 ) ,
    .I0 ( edt_decompressor_out_584 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_584 ) ) ;
and ( 
    .Z ( edt_scan_in_249 ) ,
    .I0 ( edt_decompressor_out_249 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_249 ) ) ;
and ( 
    .Z ( edt_scan_in_583 ) ,
    .I0 ( edt_decompressor_out_583 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_583 ) ) ;
and ( 
    .Z ( edt_scan_in_508 ) ,
    .I0 ( edt_decompressor_out_508 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_508 ) ) ;
and ( 
    .Z ( edt_scan_in_250 ) ,
    .I0 ( edt_decompressor_out_250 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_250 ) ) ;
and ( 
    .Z ( edt_scan_in_509 ) ,
    .I0 ( edt_decompressor_out_509 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_509 ) ) ;
and ( 
    .Z ( edt_scan_in_251 ) ,
    .I0 ( edt_decompressor_out_251 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_251 ) ) ;
and ( 
    .Z ( edt_scan_in_506 ) ,
    .I0 ( edt_decompressor_out_506 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_506 ) ) ;
and ( 
    .Z ( edt_scan_in_252 ) ,
    .I0 ( edt_decompressor_out_252 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_252 ) ) ;
and ( 
    .Z ( edt_scan_in_507 ) ,
    .I0 ( edt_decompressor_out_507 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_507 ) ) ;
and ( 
    .Z ( edt_scan_in_504 ) ,
    .I0 ( edt_decompressor_out_504 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_504 ) ) ;
and ( 
    .Z ( edt_scan_in_505 ) ,
    .I0 ( edt_decompressor_out_505 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_505 ) ) ;
and ( 
    .Z ( edt_scan_in_502 ) ,
    .I0 ( edt_decompressor_out_502 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_502 ) ) ;
and ( 
    .Z ( edt_scan_in_503 ) ,
    .I0 ( edt_decompressor_out_503 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_503 ) ) ;
and ( 
    .Z ( edt_scan_in_500 ) ,
    .I0 ( edt_decompressor_out_500 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_500 ) ) ;
and ( 
    .Z ( edt_scan_in_501 ) ,
    .I0 ( edt_decompressor_out_501 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_501 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U50.AB ) ,
    .I0 ( constant_shift_controller_i.n210 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U50.CD ) ,
    .I0 ( edt_channels_in_4 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U50.ZN ) ,
    .I0 ( constant_shift_controller_i.U50.AB ) ,
    .I1 ( constant_shift_controller_i.U50.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N166 ) ,
    .IN ( constant_shift_controller_i.U50.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U51.AB ) ,
    .I0 ( constant_shift_controller_i.n240 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U51.CD ) ,
    .I0 ( edt_channels_in_3 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U51.ZN ) ,
    .I0 ( constant_shift_controller_i.U51.AB ) ,
    .I1 ( constant_shift_controller_i.U51.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N158 ) ,
    .IN ( constant_shift_controller_i.U51.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_774 ) ,
    .I0 ( edt_decompressor_out_774 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_774 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U52.AB ) ,
    .I0 ( edt_channels_in_1 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U52.CD ) ,
    .I0 ( constant_shift_controller_i.n380 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U52.ZN ) ,
    .I0 ( constant_shift_controller_i.U52.AB ) ,
    .I1 ( constant_shift_controller_i.U52.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N149 ) ,
    .IN ( constant_shift_controller_i.U52.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_773 ) ,
    .I0 ( edt_decompressor_out_773 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_773 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U53.AB ) ,
    .I0 ( constant_shift_controller_i.n270 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U53.CD ) ,
    .I0 ( edt_channels_in_2 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U53.ZN ) ,
    .I0 ( constant_shift_controller_i.U53.AB ) ,
    .I1 ( constant_shift_controller_i.U53.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N150 ) ,
    .IN ( constant_shift_controller_i.U53.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U54.AB ) ,
    .I0 ( constant_shift_controller_i.n390 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U54.CD ) ,
    .I0 ( edt_channels_in_1 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U54.ZN ) ,
    .I0 ( constant_shift_controller_i.U54.AB ) ,
    .I1 ( constant_shift_controller_i.U54.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N142 ) ,
    .IN ( constant_shift_controller_i.U54.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U55.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_8 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U55.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U55.ZN ) ,
    .I0 ( constant_shift_controller_i.U55.AB ) ,
    .I1 ( constant_shift_controller_i.U55.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_8 ) ,
    .IN ( constant_shift_controller_i.U55.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_770 ) ,
    .I0 ( edt_decompressor_out_770 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_770 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U56.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_10 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U56.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n370 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U56.ZN ) ,
    .I0 ( constant_shift_controller_i.U56.AB ) ,
    .I1 ( constant_shift_controller_i.U56.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_10 ) ,
    .IN ( constant_shift_controller_i.U56.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_769 ) ,
    .I0 ( edt_decompressor_out_769 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_769 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U57.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_12 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U57.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n330 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U57.ZN ) ,
    .I0 ( constant_shift_controller_i.U57.AB ) ,
    .I1 ( constant_shift_controller_i.U57.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_12 ) ,
    .IN ( constant_shift_controller_i.U57.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_772 ) ,
    .I0 ( edt_decompressor_out_772 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_772 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U58.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_13 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U58.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n310 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U58.ZN ) ,
    .I0 ( constant_shift_controller_i.U58.AB ) ,
    .I1 ( constant_shift_controller_i.U58.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_13 ) ,
    .IN ( constant_shift_controller_i.U58.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_771 ) ,
    .I0 ( edt_decompressor_out_771 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_771 ) ) ;
and ( 
    .Z ( edt_scan_in_766 ) ,
    .I0 ( edt_decompressor_out_766 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_766 ) ) ;
and ( 
    .Z ( edt_scan_in_765 ) ,
    .I0 ( edt_decompressor_out_765 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_765 ) ) ;
and ( 
    .Z ( edt_scan_in_264 ) ,
    .I0 ( edt_decompressor_out_264 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_264 ) ) ;
and ( 
    .Z ( edt_scan_in_768 ) ,
    .I0 ( edt_decompressor_out_768 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_768 ) ) ;
and ( 
    .Z ( edt_scan_in_767 ) ,
    .I0 ( edt_decompressor_out_767 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_767 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N43 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N42 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N41 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_1.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n660 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_6 ) ) ;
and ( 
    .Z ( edt_scan_in_303 ) ,
    .I0 ( edt_decompressor_out_303 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_303 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N70 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n660 ) ) ;
and ( 
    .Z ( edt_scan_in_611 ) ,
    .I0 ( edt_decompressor_out_611 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_611 ) ) ;
and ( 
    .Z ( edt_scan_in_304 ) ,
    .I0 ( edt_decompressor_out_304 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_304 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n670 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_5 ) ) ;
and ( 
    .Z ( edt_scan_in_610 ) ,
    .I0 ( edt_decompressor_out_610 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_610 ) ) ;
and ( 
    .Z ( edt_scan_in_305 ) ,
    .I0 ( edt_decompressor_out_305 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_305 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N69 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n670 ) ) ;
and ( 
    .Z ( edt_scan_in_609 ) ,
    .I0 ( edt_decompressor_out_609 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_609 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n680 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_4 ) ) ;
and ( 
    .Z ( edt_scan_in_608 ) ,
    .I0 ( edt_decompressor_out_608 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_608 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N68 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n680 ) ) ;
and ( 
    .Z ( edt_scan_in_528 ) ,
    .I0 ( edt_decompressor_out_528 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_528 ) ) ;
and ( 
    .Z ( edt_scan_in_607 ) ,
    .I0 ( edt_decompressor_out_607 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_607 ) ) ;
and ( 
    .Z ( edt_scan_in_529 ) ,
    .I0 ( edt_decompressor_out_529 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_529 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N79 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_605 ) ,
    .I0 ( edt_decompressor_out_605 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_605 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N78 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_604 ) ,
    .I0 ( edt_decompressor_out_604 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_604 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N77 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_603 ) ,
    .I0 ( edt_decompressor_out_603 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_603 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N76 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_602 ) ,
    .I0 ( edt_decompressor_out_602 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_602 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N75 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N74 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N73 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_520 ) ,
    .I0 ( edt_decompressor_out_520 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_520 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N72 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_8_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_8_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_8_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_8_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_8_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_521 ) ,
    .I0 ( edt_decompressor_out_521 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_521 ) ) ;
and ( 
    .Z ( edt_scan_in_522 ) ,
    .I0 ( edt_decompressor_out_522 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_522 ) ) ;
and ( 
    .Z ( edt_scan_in_524 ) ,
    .I0 ( edt_decompressor_out_524 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_524 ) ) ;
and ( 
    .Z ( edt_scan_in_525 ) ,
    .I0 ( edt_decompressor_out_525 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_525 ) ) ;
and ( 
    .Z ( edt_scan_in_526 ) ,
    .I0 ( edt_decompressor_out_526 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_526 ) ) ;
and ( 
    .Z ( edt_scan_in_527 ) ,
    .I0 ( edt_decompressor_out_527 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_527 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N76 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n200 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N61 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n231 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N31 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n380 ) ) ;
and ( 
    .Z ( edt_scan_in_758 ) ,
    .I0 ( edt_decompressor_out_758 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_758 ) ) ;
and ( 
    .Z ( edt_scan_in_152 ) ,
    .I0 ( edt_decompressor_out_152 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_152 ) ) ;
and ( 
    .Z ( edt_scan_in_488 ) ,
    .I0 ( edt_decompressor_out_488 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_488 ) ) ;
and ( 
    .Z ( edt_scan_in_489 ) ,
    .I0 ( edt_decompressor_out_489 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_489 ) ) ;
and ( 
    .Z ( edt_scan_in_483 ) ,
    .I0 ( edt_decompressor_out_483 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_483 ) ) ;
and ( 
    .Z ( edt_scan_in_484 ) ,
    .I0 ( edt_decompressor_out_484 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_484 ) ) ;
and ( 
    .Z ( edt_scan_in_485 ) ,
    .I0 ( edt_decompressor_out_485 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_485 ) ) ;
and ( 
    .Z ( edt_scan_in_144 ) ,
    .I0 ( edt_decompressor_out_144 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_144 ) ) ;
and ( 
    .Z ( edt_scan_in_487 ) ,
    .I0 ( edt_decompressor_out_487 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_487 ) ) ;
and ( 
    .Z ( edt_scan_in_143 ) ,
    .I0 ( edt_decompressor_out_143 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_143 ) ) ;
and ( 
    .Z ( edt_scan_in_479 ) ,
    .I0 ( edt_decompressor_out_479 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_479 ) ) ;
and ( 
    .Z ( edt_scan_in_146 ) ,
    .I0 ( edt_decompressor_out_146 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_146 ) ) ;
and ( 
    .Z ( edt_scan_in_480 ) ,
    .I0 ( edt_decompressor_out_480 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_480 ) ) ;
and ( 
    .Z ( edt_scan_in_145 ) ,
    .I0 ( edt_decompressor_out_145 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_145 ) ) ;
and ( 
    .Z ( edt_scan_in_148 ) ,
    .I0 ( edt_decompressor_out_148 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_148 ) ) ;
and ( 
    .Z ( edt_scan_in_482 ) ,
    .I0 ( edt_decompressor_out_482 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_482 ) ) ;
and ( 
    .Z ( edt_scan_in_147 ) ,
    .I0 ( edt_decompressor_out_147 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_147 ) ) ;
and ( 
    .Z ( edt_scan_in_150 ) ,
    .I0 ( edt_decompressor_out_150 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_150 ) ) ;
and ( 
    .Z ( edt_scan_in_149 ) ,
    .I0 ( edt_decompressor_out_149 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_149 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n290 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n481 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N149 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_6.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N122 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N150 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N123 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N120 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_2_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_2_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_2_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_2_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_2_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N121 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_1.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N126 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_6.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N124 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N125 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_14_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_14_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_14_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_14_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_14_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_161 ) ,
    .I0 ( edt_decompressor_out_161 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_161 ) ) ;
and ( 
    .Z ( edt_scan_in_163 ) ,
    .I0 ( edt_decompressor_out_163 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_163 ) ) ;
and ( 
    .Z ( edt_scan_in_153 ) ,
    .I0 ( edt_decompressor_out_153 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_153 ) ) ;
and ( 
    .Z ( edt_scan_in_155 ) ,
    .I0 ( edt_decompressor_out_155 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_155 ) ) ;
and ( 
    .Z ( edt_scan_in_156 ) ,
    .I0 ( edt_decompressor_out_156 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_156 ) ) ;
and ( 
    .Z ( edt_scan_in_157 ) ,
    .I0 ( edt_decompressor_out_157 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_157 ) ) ;
and ( 
    .Z ( edt_scan_in_158 ) ,
    .I0 ( edt_decompressor_out_158 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_158 ) ) ;
and ( 
    .Z ( edt_scan_in_159 ) ,
    .I0 ( edt_decompressor_out_159 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_159 ) ) ;
and ( 
    .Z ( edt_scan_in_160 ) ,
    .I0 ( edt_decompressor_out_160 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_160 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N120 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1010 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N8 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n390 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N32 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n210 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N40 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n180 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N16 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n270 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N24 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n240 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N112 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n310 ) ) ;
and ( 
    .Z ( edt_scan_in_499 ) ,
    .I0 ( edt_decompressor_out_499 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_499 ) ) ;
and ( 
    .Z ( edt_scan_in_498 ) ,
    .I0 ( edt_decompressor_out_498 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_498 ) ) ;
and ( 
    .Z ( edt_scan_in_497 ) ,
    .I0 ( edt_decompressor_out_497 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_497 ) ) ;
and ( 
    .Z ( edt_scan_in_496 ) ,
    .I0 ( edt_decompressor_out_496 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_496 ) ) ;
and ( 
    .Z ( edt_scan_in_495 ) ,
    .I0 ( edt_decompressor_out_495 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_495 ) ) ;
and ( 
    .Z ( edt_scan_in_494 ) ,
    .I0 ( edt_decompressor_out_494 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_494 ) ) ;
and ( 
    .Z ( edt_scan_in_493 ) ,
    .I0 ( edt_decompressor_out_493 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_493 ) ) ;
and ( 
    .Z ( edt_scan_in_492 ) ,
    .I0 ( edt_decompressor_out_492 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_492 ) ) ;
and ( 
    .Z ( edt_scan_in_491 ) ,
    .I0 ( edt_decompressor_out_491 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_491 ) ) ;
and ( 
    .Z ( edt_scan_in_490 ) ,
    .I0 ( edt_decompressor_out_490 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_490 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U41.AB ) ,
    .I0 ( constant_shift_controller_i.n3 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U41.CD ) ,
    .I0 ( edt_channels_in_10 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U41.ZN ) ,
    .I0 ( constant_shift_controller_i.U41.AB ) ,
    .I1 ( constant_shift_controller_i.U41.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N214 ) ,
    .IN ( constant_shift_controller_i.U41.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U40.AB ) ,
    .I0 ( edt_channels_in_5 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U40.CD ) ,
    .I0 ( constant_shift_controller_i.n170 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U40.ZN ) ,
    .I0 ( constant_shift_controller_i.U40.AB ) ,
    .I1 ( constant_shift_controller_i.U40.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N209 ) ,
    .IN ( constant_shift_controller_i.U40.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U43.AB ) ,
    .I0 ( edt_channels_in_4 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U43.CD ) ,
    .I0 ( constant_shift_controller_i.n200 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U43.ZN ) ,
    .I0 ( constant_shift_controller_i.U43.AB ) ,
    .I1 ( constant_shift_controller_i.U43.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N194 ) ,
    .IN ( constant_shift_controller_i.U43.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U42.AB ) ,
    .I0 ( constant_shift_controller_i.n6 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U42.CD ) ,
    .I0 ( edt_channels_in_9 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U42.ZN ) ,
    .I0 ( constant_shift_controller_i.U42.AB ) ,
    .I1 ( constant_shift_controller_i.U42.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N206 ) ,
    .IN ( constant_shift_controller_i.U42.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U45.AB ) ,
    .I0 ( constant_shift_controller_i.n1270 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U45.CD ) ,
    .I0 ( edt_channels_in_7 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U45.ZN ) ,
    .I0 ( constant_shift_controller_i.U45.AB ) ,
    .I1 ( constant_shift_controller_i.U45.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N190 ) ,
    .IN ( constant_shift_controller_i.U45.ZN ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U44.AB ) ,
    .I0 ( constant_shift_controller_i.n810 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U44.CD ) ,
    .I0 ( edt_channels_in_8 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U44.ZN ) ,
    .I0 ( constant_shift_controller_i.U44.AB ) ,
    .I1 ( constant_shift_controller_i.U44.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N198 ) ,
    .IN ( constant_shift_controller_i.U44.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_278 ) ,
    .I0 ( edt_decompressor_out_278 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_278 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U47.AB ) ,
    .I0 ( constant_shift_controller_i.n1510 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U47.CD ) ,
    .I0 ( edt_channels_in_6 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U47.ZN ) ,
    .I0 ( constant_shift_controller_i.U47.AB ) ,
    .I1 ( constant_shift_controller_i.U47.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N182 ) ,
    .IN ( constant_shift_controller_i.U47.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_279 ) ,
    .I0 ( edt_decompressor_out_279 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_279 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U46.AB ) ,
    .I0 ( edt_channels_in_3 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U46.CD ) ,
    .I0 ( constant_shift_controller_i.n231 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U46.ZN ) ,
    .I0 ( constant_shift_controller_i.U46.AB ) ,
    .I1 ( constant_shift_controller_i.U46.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N179 ) ,
    .IN ( constant_shift_controller_i.U46.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_276 ) ,
    .I0 ( edt_decompressor_out_276 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_276 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U49.AB ) ,
    .I0 ( edt_channels_in_2 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U49.CD ) ,
    .I0 ( constant_shift_controller_i.n260 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U49.ZN ) ,
    .I0 ( constant_shift_controller_i.U49.AB ) ,
    .I1 ( constant_shift_controller_i.U49.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N164 ) ,
    .IN ( constant_shift_controller_i.U49.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_277 ) ,
    .I0 ( edt_decompressor_out_277 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_277 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U48.AB ) ,
    .I0 ( constant_shift_controller_i.n180 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U48.CD ) ,
    .I0 ( edt_channels_in_5 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U48.ZN ) ,
    .I0 ( constant_shift_controller_i.U48.AB ) ,
    .I1 ( constant_shift_controller_i.U48.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N174 ) ,
    .IN ( constant_shift_controller_i.U48.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_282 ) ,
    .I0 ( edt_decompressor_out_282 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_282 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N108 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_253 ) ,
    .I0 ( edt_decompressor_out_253 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_253 ) ) ;
and ( 
    .Z ( edt_scan_in_283 ) ,
    .I0 ( edt_decompressor_out_283 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_283 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N109 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_254 ) ,
    .I0 ( edt_decompressor_out_254 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_254 ) ) ;
and ( 
    .Z ( edt_scan_in_590 ) ,
    .I0 ( edt_decompressor_out_590 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_590 ) ) ;
and ( 
    .Z ( edt_scan_in_280 ) ,
    .I0 ( edt_decompressor_out_280 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_280 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N110 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_589 ) ,
    .I0 ( edt_decompressor_out_589 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_589 ) ) ;
and ( 
    .Z ( edt_scan_in_281 ) ,
    .I0 ( edt_decompressor_out_281 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N111 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N104 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N105 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_12_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_12_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_12_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_12_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_12_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_586 ) ,
    .I0 ( edt_decompressor_out_586 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_586 ) ) ;
and ( 
    .Z ( edt_scan_in_284 ) ,
    .I0 ( edt_decompressor_out_284 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_4 ) ) ;
and ( 
    .Z ( edt_scan_in_468 ) ,
    .I0 ( edt_decompressor_out_468 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_468 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N206 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_7 ) ) ;
and ( 
    .Z ( edt_scan_in_467 ) ,
    .I0 ( edt_decompressor_out_467 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_467 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_6 ) ) ;
and ( 
    .Z ( edt_scan_in_462 ) ,
    .I0 ( edt_decompressor_out_462 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_462 ) ) ;
and ( 
    .Z ( edt_scan_in_461 ) ,
    .I0 ( edt_decompressor_out_461 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_461 ) ) ;
and ( 
    .Z ( edt_scan_in_460 ) ,
    .I0 ( edt_decompressor_out_460 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_460 ) ) ;
and ( 
    .Z ( edt_scan_in_459 ) ,
    .I0 ( edt_decompressor_out_459 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_459 ) ) ;
and ( 
    .Z ( edt_scan_in_466 ) ,
    .I0 ( edt_decompressor_out_466 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_466 ) ) ;
and ( 
    .Z ( edt_scan_in_465 ) ,
    .I0 ( edt_decompressor_out_465 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_465 ) ) ;
and ( 
    .Z ( edt_scan_in_464 ) ,
    .I0 ( edt_decompressor_out_464 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_464 ) ) ;
and ( 
    .Z ( edt_scan_in_463 ) ,
    .I0 ( edt_decompressor_out_463 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_463 ) ) ;
and ( 
    .Z ( edt_scan_in_657 ) ,
    .I0 ( edt_decompressor_out_657 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_657 ) ) ;
and ( 
    .Z ( edt_scan_in_356 ) ,
    .I0 ( edt_decompressor_out_356 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_356 ) ) ;
and ( 
    .Z ( edt_scan_in_658 ) ,
    .I0 ( edt_decompressor_out_658 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_658 ) ) ;
and ( 
    .Z ( edt_scan_in_355 ) ,
    .I0 ( edt_decompressor_out_355 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_355 ) ) ;
and ( 
    .Z ( edt_scan_in_659 ) ,
    .I0 ( edt_decompressor_out_659 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_659 ) ) ;
and ( 
    .Z ( edt_scan_in_660 ) ,
    .I0 ( edt_decompressor_out_660 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_660 ) ) ;
and ( 
    .Z ( edt_scan_in_653 ) ,
    .I0 ( edt_decompressor_out_653 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_653 ) ) ;
and ( 
    .Z ( edt_scan_in_654 ) ,
    .I0 ( edt_decompressor_out_654 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_654 ) ) ;
and ( 
    .Z ( edt_scan_in_655 ) ,
    .I0 ( edt_decompressor_out_655 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_655 ) ) ;
and ( 
    .Z ( edt_scan_in_350 ) ,
    .I0 ( edt_decompressor_out_350 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_350 ) ) ;
and ( 
    .Z ( edt_scan_in_656 ) ,
    .I0 ( edt_decompressor_out_656 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_656 ) ) ;
and ( 
    .Z ( edt_scan_in_349 ) ,
    .I0 ( edt_decompressor_out_349 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_349 ) ) ;
and ( 
    .Z ( edt_scan_in_348 ) ,
    .I0 ( edt_decompressor_out_348 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_348 ) ) ;
and ( 
    .Z ( edt_scan_in_347 ) ,
    .I0 ( edt_decompressor_out_347 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_347 ) ) ;
and ( 
    .Z ( edt_scan_in_354 ) ,
    .I0 ( edt_decompressor_out_354 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_354 ) ) ;
and ( 
    .Z ( edt_scan_in_353 ) ,
    .I0 ( edt_decompressor_out_353 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_353 ) ) ;
and ( 
    .Z ( edt_scan_in_661 ) ,
    .I0 ( edt_decompressor_out_661 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_661 ) ) ;
and ( 
    .Z ( edt_scan_in_352 ) ,
    .I0 ( edt_decompressor_out_352 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_352 ) ) ;
and ( 
    .Z ( edt_scan_in_662 ) ,
    .I0 ( edt_decompressor_out_662 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_662 ) ) ;
and ( 
    .Z ( edt_scan_in_351 ) ,
    .I0 ( edt_decompressor_out_351 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_351 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N57 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_1.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N56 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N59 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N58 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N61 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_5.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N60 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N63 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N62 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_6_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_6_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_6_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_6_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_6_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_668 ) ,
    .I0 ( edt_decompressor_out_668 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_668 ) ) ;
and ( 
    .Z ( edt_scan_in_365 ) ,
    .I0 ( edt_decompressor_out_365 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_365 ) ) ;
and ( 
    .Z ( edt_scan_in_667 ) ,
    .I0 ( edt_decompressor_out_667 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_667 ) ) ;
and ( 
    .Z ( edt_scan_in_366 ) ,
    .I0 ( edt_decompressor_out_366 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_366 ) ) ;
and ( 
    .Z ( edt_scan_in_670 ) ,
    .I0 ( edt_decompressor_out_670 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_670 ) ) ;
and ( 
    .Z ( edt_scan_in_669 ) ,
    .I0 ( edt_decompressor_out_669 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_669 ) ) ;
and ( 
    .Z ( edt_scan_in_664 ) ,
    .I0 ( edt_decompressor_out_664 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_664 ) ) ;
and ( 
    .Z ( edt_scan_in_663 ) ,
    .I0 ( edt_decompressor_out_663 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_663 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N40 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_256 ) ,
    .I0 ( edt_decompressor_out_256 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_256 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N47 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_255 ) ,
    .I0 ( edt_decompressor_out_255 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_255 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N46 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_258 ) ,
    .I0 ( edt_decompressor_out_258 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_258 ) ) ;
and ( 
    .Z ( edt_scan_in_478 ) ,
    .I0 ( edt_decompressor_out_478 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_478 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N45 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_477 ) ,
    .I0 ( edt_decompressor_out_477 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_477 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N44 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_4_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_4_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_4_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_4_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_4_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_260 ) ,
    .I0 ( edt_decompressor_out_260 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_260 ) ) ;
and ( 
    .Z ( edt_scan_in_259 ) ,
    .I0 ( edt_decompressor_out_259 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_259 ) ) ;
and ( 
    .Z ( edt_scan_in_262 ) ,
    .I0 ( edt_decompressor_out_262 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_262 ) ) ;
and ( 
    .Z ( edt_scan_in_474 ) ,
    .I0 ( edt_decompressor_out_474 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_474 ) ) ;
and ( 
    .Z ( edt_scan_in_261 ) ,
    .I0 ( edt_decompressor_out_261 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_261 ) ) ;
and ( 
    .Z ( edt_scan_in_473 ) ,
    .I0 ( edt_decompressor_out_473 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_473 ) ) ;
and ( 
    .Z ( edt_scan_in_476 ) ,
    .I0 ( edt_decompressor_out_476 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_476 ) ) ;
and ( 
    .Z ( edt_scan_in_475 ) ,
    .I0 ( edt_decompressor_out_475 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_475 ) ) ;
and ( 
    .Z ( edt_scan_in_470 ) ,
    .I0 ( edt_decompressor_out_470 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_470 ) ) ;
and ( 
    .Z ( edt_scan_in_469 ) ,
    .I0 ( edt_decompressor_out_469 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_469 ) ) ;
and ( 
    .Z ( edt_scan_in_472 ) ,
    .I0 ( edt_decompressor_out_472 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_472 ) ) ;
and ( 
    .Z ( edt_scan_in_471 ) ,
    .I0 ( edt_decompressor_out_471 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_471 ) ) ;
and ( 
    .Z ( edt_scan_in_763 ) ,
    .I0 ( edt_decompressor_out_763 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_763 ) ) ;
and ( 
    .Z ( edt_scan_in_764 ) ,
    .I0 ( edt_decompressor_out_764 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_764 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n250 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_0 ) ) ;
and ( 
    .Z ( edt_scan_in_760 ) ,
    .I0 ( edt_decompressor_out_760 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_760 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_3 ) ) ;
and ( 
    .Z ( edt_scan_in_761 ) ,
    .I0 ( edt_decompressor_out_761 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N209 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_2.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_2 ) ) ;
and ( 
    .Z ( edt_scan_in_762 ) ,
    .I0 ( edt_decompressor_out_762 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_762 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_5 ) ) ;
and ( 
    .Z ( edt_scan_in_754 ) ,
    .I0 ( edt_decompressor_out_754 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_754 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_4 ) ) ;
and ( 
    .Z ( edt_scan_in_755 ) ,
    .I0 ( edt_decompressor_out_755 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_755 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N214 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_7 ) ) ;
and ( 
    .Z ( edt_scan_in_757 ) ,
    .I0 ( edt_decompressor_out_757 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_757 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_10_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_10_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_10_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_10_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_10_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N33 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n970 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n970 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N15 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N14 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_6.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N13 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_5.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N12 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N11 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N10 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N9 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_1.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N8 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_0_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_0_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_0_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_0_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_0_reg_0.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n950 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N35 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n950 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n960 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N34 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n960 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N245 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_6.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n930 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N37 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n930 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n940 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n127 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N36 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n940 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_14_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_14_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_14_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_14_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_14_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_14_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n920 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N38 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n920 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N63 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n720 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n720 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N182 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N49 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n840 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N179 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_4.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n840 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N50 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n830 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N94 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_6.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n830 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N95 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_7.QT ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N51 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n820 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N92 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_4.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n820 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_6_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_6_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_6_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_6_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_6_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N93 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_5.QT ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N52 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n811 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N90 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_2.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n811 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N91 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N88 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N89 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_10_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_10_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_10_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_10_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_10_reg_1.QT ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N104 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n330 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N48 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1510 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N56 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1270 ) ) ;
and ( 
    .Z ( edt_scan_in_457 ) ,
    .I0 ( edt_decompressor_out_457 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_457 ) ) ;
and ( 
    .Z ( edt_scan_in_458 ) ,
    .I0 ( edt_decompressor_out_458 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_458 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n912 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n231 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_2 ) ) ;
and ( 
    .Z ( edt_scan_in_451 ) ,
    .I0 ( edt_decompressor_out_451 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_451 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N174 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n260 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N224 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_1.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_1 ) ) ;
and ( 
    .Z ( edt_scan_in_452 ) ,
    .I0 ( edt_decompressor_out_452 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_452 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_0 ) ) ;
and ( 
    .Z ( edt_scan_in_449 ) ,
    .I0 ( edt_decompressor_out_449 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_449 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N230 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_7 ) ) ;
and ( 
    .Z ( edt_scan_in_450 ) ,
    .I0 ( edt_decompressor_out_450 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_450 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n491 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n380 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_6 ) ) ;
and ( 
    .Z ( edt_scan_in_455 ) ,
    .I0 ( edt_decompressor_out_455 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_455 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1400 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_5 ) ) ;
and ( 
    .Z ( edt_scan_in_456 ) ,
    .I0 ( edt_decompressor_out_456 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_456 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_5_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_5_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_5_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_5_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_5_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n170 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_12_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_12_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_12_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_12_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_12_4 ) ) ;
and ( 
    .Z ( edt_scan_in_453 ) ,
    .I0 ( edt_decompressor_out_453 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_453 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n200 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_4 ) ) ;
and ( 
    .Z ( edt_scan_in_454 ) ,
    .I0 ( edt_decompressor_out_454 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_454 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U90.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n380 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U90.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n390 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U90.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n400 ) ) ;
nand ( 
    .Z ( edt_channels_out_from_constant_shift_control_0 ) ,
    .I0 ( constant_shift_controller_i.U90.AB ) ,
    .I1 ( constant_shift_controller_i.U90.CD ) ,
    .I2 ( constant_shift_controller_i.U90.EF ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n400 ) ,
    .IN ( constant_shift_controller_i.n130 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U92.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_14 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U92.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n1010 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U92.ZN ) ,
    .I0 ( constant_shift_controller_i.U92.AB ) ,
    .I1 ( constant_shift_controller_i.U92.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_14 ) ,
    .IN ( constant_shift_controller_i.U92.ZN ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n3 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_9_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_9_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_9_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_9_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_9_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n130 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_7.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_7.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_7.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_7.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_7.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N83 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n560 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N117 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_5.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n560 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N116 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N119 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N118 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_21 ) ,
    .I0 ( edt_decompressor_out_21 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_21 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N113 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_22 ) ,
    .I0 ( edt_decompressor_out_22 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_22 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N112 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_23 ) ,
    .I0 ( edt_decompressor_out_23 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_23 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N115 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_24 ) ,
    .I0 ( edt_decompressor_out_24 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_24 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N114 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_13_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_13_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_13_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_13_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_13_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_25 ) ,
    .I0 ( edt_decompressor_out_25 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_25 ) ) ;
and ( 
    .Z ( edt_scan_in_26 ) ,
    .I0 ( edt_decompressor_out_26 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_26 ) ) ;
and ( 
    .Z ( edt_scan_in_27 ) ,
    .I0 ( edt_decompressor_out_27 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_27 ) ) ;
and ( 
    .Z ( edt_scan_in_28 ) ,
    .I0 ( edt_decompressor_out_28 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_28 ) ) ;
and ( 
    .Z ( edt_scan_in_29 ) ,
    .I0 ( edt_decompressor_out_29 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_29 ) ) ;
and ( 
    .Z ( edt_scan_in_30 ) ,
    .I0 ( edt_decompressor_out_30 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_30 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n740 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N60 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n740 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n750 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N59 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n750 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n760 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N58 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n760 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n770 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N57 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n770 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n730 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N62 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n730 ) ) ;
and ( 
    .Z ( edt_scan_in_32 ) ,
    .I0 ( edt_decompressor_out_32 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_32 ) ) ;
and ( 
    .Z ( edt_scan_in_31 ) ,
    .I0 ( edt_decompressor_out_31 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_31 ) ) ;
and ( 
    .Z ( edt_scan_in_34 ) ,
    .I0 ( edt_decompressor_out_34 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_34 ) ) ;
and ( 
    .Z ( edt_scan_in_33 ) ,
    .I0 ( edt_decompressor_out_33 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_33 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N50 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_3 ) ) ;
and ( 
    .Z ( edt_scan_in_36 ) ,
    .I0 ( edt_decompressor_out_36 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_36 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N51 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_2 ) ) ;
and ( 
    .Z ( edt_scan_in_35 ) ,
    .I0 ( edt_decompressor_out_35 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_35 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N48 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N49 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_1.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_0 ) ) ;
and ( 
    .Z ( edt_scan_in_37 ) ,
    .I0 ( edt_decompressor_out_37 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_37 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_6.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N158 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_7 ) ) ;
and ( 
    .Z ( edt_scan_in_40 ) ,
    .I0 ( edt_decompressor_out_40 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_40 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N55 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_6 ) ) ;
and ( 
    .Z ( edt_scan_in_39 ) ,
    .I0 ( edt_decompressor_out_39 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_39 ) ) ;
and ( 
    .Z ( edt_scan_in_666 ) ,
    .I0 ( edt_decompressor_out_666 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_666 ) ) ;
and ( 
    .Z ( edt_scan_in_359 ) ,
    .I0 ( edt_decompressor_out_359 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_359 ) ) ;
and ( 
    .Z ( edt_scan_in_665 ) ,
    .I0 ( edt_decompressor_out_665 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_665 ) ) ;
and ( 
    .Z ( edt_scan_in_360 ) ,
    .I0 ( edt_decompressor_out_360 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_360 ) ) ;
and ( 
    .Z ( edt_scan_in_357 ) ,
    .I0 ( edt_decompressor_out_357 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_357 ) ) ;
and ( 
    .Z ( edt_scan_in_358 ) ,
    .I0 ( edt_decompressor_out_358 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_358 ) ) ;
and ( 
    .Z ( edt_scan_in_363 ) ,
    .I0 ( edt_decompressor_out_363 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_363 ) ) ;
and ( 
    .Z ( edt_scan_in_364 ) ,
    .I0 ( edt_decompressor_out_364 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_364 ) ) ;
and ( 
    .Z ( edt_scan_in_672 ) ,
    .I0 ( edt_decompressor_out_672 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_672 ) ) ;
and ( 
    .Z ( edt_scan_in_361 ) ,
    .I0 ( edt_decompressor_out_361 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_361 ) ) ;
and ( 
    .Z ( edt_scan_in_671 ) ,
    .I0 ( edt_decompressor_out_671 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_671 ) ) ;
and ( 
    .Z ( edt_scan_in_362 ) ,
    .I0 ( edt_decompressor_out_362 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_362 ) ) ;
and ( 
    .Z ( edt_scan_in_556 ) ,
    .I0 ( edt_decompressor_out_556 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_556 ) ) ;
and ( 
    .Z ( edt_scan_in_555 ) ,
    .I0 ( edt_decompressor_out_555 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_555 ) ) ;
and ( 
    .Z ( edt_scan_in_558 ) ,
    .I0 ( edt_decompressor_out_558 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_558 ) ) ;
and ( 
    .Z ( edt_scan_in_557 ) ,
    .I0 ( edt_decompressor_out_557 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_557 ) ) ;
and ( 
    .Z ( edt_scan_in_552 ) ,
    .I0 ( edt_decompressor_out_552 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_552 ) ) ;
and ( 
    .Z ( edt_scan_in_551 ) ,
    .I0 ( edt_decompressor_out_551 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_551 ) ) ;
and ( 
    .Z ( edt_scan_in_554 ) ,
    .I0 ( edt_decompressor_out_554 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_554 ) ) ;
and ( 
    .Z ( edt_scan_in_553 ) ,
    .I0 ( edt_decompressor_out_553 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_553 ) ) ;
and ( 
    .Z ( edt_scan_in_560 ) ,
    .I0 ( edt_decompressor_out_560 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_560 ) ) ;
and ( 
    .Z ( edt_scan_in_559 ) ,
    .I0 ( edt_decompressor_out_559 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_559 ) ) ;
and ( 
    .Z ( edt_scan_in_565 ) ,
    .I0 ( edt_decompressor_out_565 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_565 ) ) ;
and ( 
    .Z ( edt_scan_in_566 ) ,
    .I0 ( edt_decompressor_out_566 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_566 ) ) ;
and ( 
    .Z ( edt_scan_in_567 ) ,
    .I0 ( edt_decompressor_out_567 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_567 ) ) ;
and ( 
    .Z ( edt_scan_in_568 ) ,
    .I0 ( edt_decompressor_out_568 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_568 ) ) ;
and ( 
    .Z ( edt_scan_in_561 ) ,
    .I0 ( edt_decompressor_out_561 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_561 ) ) ;
and ( 
    .Z ( edt_scan_in_562 ) ,
    .I0 ( edt_decompressor_out_562 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_562 ) ) ;
and ( 
    .Z ( edt_scan_in_563 ) ,
    .I0 ( edt_decompressor_out_563 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_563 ) ) ;
and ( 
    .Z ( edt_scan_in_564 ) ,
    .I0 ( edt_decompressor_out_564 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_564 ) ) ;
and ( 
    .Z ( edt_scan_in_569 ) ,
    .I0 ( edt_decompressor_out_569 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_569 ) ) ;
and ( 
    .Z ( edt_scan_in_570 ) ,
    .I0 ( edt_decompressor_out_570 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_570 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N44 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n870 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n870 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N43 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n880 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n880 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N47 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n850 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n850 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N45 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n860 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n860 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N31 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_1 ) ,
    .I0 ( edt_decompressor_out_1 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_2 ) ,
    .I0 ( edt_decompressor_out_2 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N25 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_7 ) ,
    .I0 ( edt_decompressor_out_7 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N24 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_8 ) ,
    .I0 ( edt_decompressor_out_8 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_8 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N27 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_5 ) ,
    .I0 ( edt_decompressor_out_5 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_6 ) ,
    .I0 ( edt_decompressor_out_6 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n520 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_7 ) ) ;
and ( 
    .Z ( edt_scan_in_9 ) ,
    .I0 ( edt_decompressor_out_9 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_9 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N87 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n520 ) ) ;
and ( 
    .Z ( edt_scan_in_10 ) ,
    .I0 ( edt_decompressor_out_10 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_10 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n640 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N73 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n640 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n630 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N74 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n630 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n620 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N75 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n620 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n610 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n270 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_0 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N77 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n610 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n240 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1010 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n390 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_0 ) ) ;
and ( 
    .Z ( edt_scan_in_14 ) ,
    .I0 ( edt_decompressor_out_14 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_14 ) ) ;
and ( 
    .Z ( edt_scan_in_13 ) ,
    .I0 ( edt_decompressor_out_13 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_13 ) ) ;
and ( 
    .Z ( edt_scan_in_12 ) ,
    .I0 ( edt_decompressor_out_12 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_12 ) ) ;
and ( 
    .Z ( edt_scan_in_11 ) ,
    .I0 ( edt_decompressor_out_11 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_11 ) ) ;
and ( 
    .Z ( edt_scan_in_18 ) ,
    .I0 ( edt_decompressor_out_18 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_18 ) ) ;
and ( 
    .Z ( edt_scan_in_17 ) ,
    .I0 ( edt_decompressor_out_17 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_17 ) ) ;
and ( 
    .Z ( edt_scan_in_16 ) ,
    .I0 ( edt_decompressor_out_16 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_16 ) ) ;
and ( 
    .Z ( edt_scan_in_15 ) ,
    .I0 ( edt_decompressor_out_15 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_15 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N78 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n600 ) ) ;
and ( 
    .Z ( edt_scan_in_20 ) ,
    .I0 ( edt_decompressor_out_20 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_20 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n600 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_6 ) ) ;
and ( 
    .Z ( edt_scan_in_19 ) ,
    .I0 ( edt_decompressor_out_19 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_19 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N79 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n590 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n590 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N65 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n710 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n710 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N66 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n700 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n700 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N67 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n690 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n690 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_3 ) ) ;
and ( 
    .Z ( edt_scan_in_54 ) ,
    .I0 ( edt_decompressor_out_54 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_54 ) ) ;
and ( 
    .Z ( edt_scan_in_108 ) ,
    .I0 ( edt_decompressor_out_108 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_108 ) ) ;
and ( 
    .Z ( edt_scan_in_162 ) ,
    .I0 ( edt_decompressor_out_162 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_162 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N108 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1230 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1230 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N109 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1220 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1220 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1130 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N118 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1130 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1140 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_5 ) ) ;
and ( 
    .Z ( edt_scan_in_216 ) ,
    .I0 ( edt_decompressor_out_216 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_216 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N117 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1140 ) ) ;
and ( 
    .Z ( edt_scan_in_270 ) ,
    .I0 ( edt_decompressor_out_270 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_270 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n510 ) ,
    .IN ( constant_shift_controller_i.n250 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N89 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n510 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1120 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N119 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1120 ) ) ;
and ( 
    .Z ( edt_scan_in_231 ) ,
    .I0 ( edt_decompressor_out_231 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_231 ) ) ;
and ( 
    .Z ( edt_scan_in_232 ) ,
    .I0 ( edt_decompressor_out_232 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_232 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n490 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N86 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_6.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N87 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_7.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N84 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N85 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_5.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N82 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_2.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N83 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N80 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N81 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_9_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_9_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_9_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_9_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_9_reg_1.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n800 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N53 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n800 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n790 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N54 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n790 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n780 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N55 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n780 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n900 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N41 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n900 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n890 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N42 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n890 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_0_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_0_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_0_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_0_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_0_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n570 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N81 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n580 ) ) ;
and ( 
    .Z ( edt_scan_in_0 ) ,
    .I0 ( edt_decompressor_out_0 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n580 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_1 ) ) ;
and ( 
    .Z ( edt_scan_in_756 ) ,
    .I0 ( edt_decompressor_out_756 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_756 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N85 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n540 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n540 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N84 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n550 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n550 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_4 ) ) ;
and ( 
    .Z ( edt_scan_in_241 ) ,
    .I0 ( edt_decompressor_out_241 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_241 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N86 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n530 ) ) ;
and ( 
    .Z ( edt_scan_in_240 ) ,
    .I0 ( edt_decompressor_out_240 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_240 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n530 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_6 ) ) ;
and ( 
    .Z ( edt_scan_in_239 ) ,
    .I0 ( edt_decompressor_out_239 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_239 ) ) ;
and ( 
    .Z ( edt_scan_in_238 ) ,
    .I0 ( edt_decompressor_out_238 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_238 ) ) ;
and ( 
    .Z ( edt_scan_in_237 ) ,
    .I0 ( edt_decompressor_out_237 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_237 ) ) ;
and ( 
    .Z ( edt_scan_in_236 ) ,
    .I0 ( edt_decompressor_out_236 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_236 ) ) ;
and ( 
    .Z ( edt_scan_in_235 ) ,
    .I0 ( edt_decompressor_out_235 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_235 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N103 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1260 ) ) ;
and ( 
    .Z ( edt_scan_in_243 ) ,
    .I0 ( edt_decompressor_out_243 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_243 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1260 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N99 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n420 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n420 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N98 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n430 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n430 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N97 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n440 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n440 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1070 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N125 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1070 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1060 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N126 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1060 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1090 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N105 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1250 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N123 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1090 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1250 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1080 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N124 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1080 ) ) ;
and ( 
    .Z ( edt_scan_in_208 ) ,
    .I0 ( edt_decompressor_out_208 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_208 ) ) ;
and ( 
    .Z ( edt_scan_in_209 ) ,
    .I0 ( edt_decompressor_out_209 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_209 ) ) ;
and ( 
    .Z ( edt_scan_in_210 ) ,
    .I0 ( edt_decompressor_out_210 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_210 ) ) ;
and ( 
    .Z ( edt_scan_in_211 ) ,
    .I0 ( edt_decompressor_out_211 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_211 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1210 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N110 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1210 ) ) ;
and ( 
    .Z ( edt_scan_in_206 ) ,
    .I0 ( edt_decompressor_out_206 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_206 ) ) ;
and ( 
    .Z ( edt_scan_in_207 ) ,
    .I0 ( edt_decompressor_out_207 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_207 ) ) ;
and ( 
    .Z ( edt_scan_in_130 ) ,
    .I0 ( edt_decompressor_out_130 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_130 ) ) ;
and ( 
    .Z ( edt_scan_in_129 ) ,
    .I0 ( edt_decompressor_out_129 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_129 ) ) ;
and ( 
    .Z ( edt_scan_in_128 ) ,
    .I0 ( edt_decompressor_out_128 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_128 ) ) ;
and ( 
    .Z ( edt_scan_in_212 ) ,
    .I0 ( edt_decompressor_out_212 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_212 ) ) ;
and ( 
    .Z ( edt_scan_in_127 ) ,
    .I0 ( edt_decompressor_out_127 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_127 ) ) ;
and ( 
    .Z ( edt_scan_in_213 ) ,
    .I0 ( edt_decompressor_out_213 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_213 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n12700 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_6 ) ) ;
and ( 
    .Z ( edt_scan_in_125 ) ,
    .I0 ( edt_decompressor_out_125 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_125 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N102 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n12700 ) ) ;
and ( 
    .Z ( edt_scan_in_124 ) ,
    .I0 ( edt_decompressor_out_124 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_124 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n129 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_5 ) ) ;
and ( 
    .Z ( edt_scan_in_123 ) ,
    .I0 ( edt_decompressor_out_123 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_123 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N101 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n129 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n13000 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N100 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n13000 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n141 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N11 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n141 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N64 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_0.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N65 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_132 ) ,
    .I0 ( edt_decompressor_out_132 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_132 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N114 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1170 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N66 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_131 ) ,
    .I0 ( edt_decompressor_out_131 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_131 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1170 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N67 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_3.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N52 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_4.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N53 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_5_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_5_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_5_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_5_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_5_reg_5.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_3_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_3_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_3_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_3_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_3_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n810 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n310 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1270 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_6_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1510 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n330 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n350 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n370 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_10_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n6 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n180 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n210 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N29 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_3 ) ,
    .I0 ( edt_decompressor_out_3 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N28 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_2_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_2_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_2_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_2_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_2_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_4 ) ,
    .I0 ( edt_decompressor_out_4 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1150 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_4 ) ) ;
and ( 
    .Z ( edt_scan_in_214 ) ,
    .I0 ( edt_decompressor_out_214 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_214 ) ) ;
and ( 
    .Z ( edt_scan_in_218 ) ,
    .I0 ( edt_decompressor_out_218 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_218 ) ) ;
and ( 
    .Z ( edt_scan_in_217 ) ,
    .I0 ( edt_decompressor_out_217 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_217 ) ) ;
and ( 
    .Z ( edt_scan_in_139 ) ,
    .I0 ( edt_decompressor_out_139 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_139 ) ) ;
and ( 
    .Z ( edt_scan_in_140 ) ,
    .I0 ( edt_decompressor_out_140 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_140 ) ) ;
and ( 
    .Z ( edt_scan_in_137 ) ,
    .I0 ( edt_decompressor_out_137 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_137 ) ) ;
and ( 
    .Z ( edt_scan_in_224 ) ,
    .I0 ( edt_decompressor_out_224 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_224 ) ) ;
and ( 
    .Z ( edt_scan_in_138 ) ,
    .I0 ( edt_decompressor_out_138 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_138 ) ) ;
and ( 
    .Z ( edt_scan_in_223 ) ,
    .I0 ( edt_decompressor_out_223 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_223 ) ) ;
and ( 
    .Z ( edt_scan_in_135 ) ,
    .I0 ( edt_decompressor_out_135 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_135 ) ) ;
and ( 
    .Z ( edt_scan_in_133 ) ,
    .I0 ( edt_decompressor_out_133 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_133 ) ) ;
and ( 
    .Z ( edt_scan_in_134 ) ,
    .I0 ( edt_decompressor_out_134 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_134 ) ) ;
and ( 
    .Z ( edt_scan_in_141 ) ,
    .I0 ( edt_decompressor_out_141 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_141 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1190 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_7 ) ) ;
and ( 
    .Z ( edt_scan_in_142 ) ,
    .I0 ( edt_decompressor_out_142 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_142 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N23 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1190 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n128 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_6 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N22 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n128 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n131 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N21 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n131 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n132 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_4 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N20 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n132 ) ) ;
and ( 
    .Z ( edt_scan_in_186 ) ,
    .I0 ( edt_decompressor_out_186 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_186 ) ) ;
and ( 
    .Z ( edt_scan_in_187 ) ,
    .I0 ( edt_decompressor_out_187 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_187 ) ) ;
and ( 
    .Z ( edt_scan_in_184 ) ,
    .I0 ( edt_decompressor_out_184 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_184 ) ) ;
and ( 
    .Z ( edt_scan_in_185 ) ,
    .I0 ( edt_decompressor_out_185 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_185 ) ) ;
and ( 
    .Z ( edt_scan_in_190 ) ,
    .I0 ( edt_decompressor_out_190 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_190 ) ) ;
and ( 
    .Z ( edt_scan_in_191 ) ,
    .I0 ( edt_decompressor_out_191 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_191 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n14000 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_4 ) ) ;
and ( 
    .Z ( edt_scan_in_188 ) ,
    .I0 ( edt_decompressor_out_188 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_188 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N12 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n14000 ) ) ;
and ( 
    .Z ( edt_scan_in_189 ) ,
    .I0 ( edt_decompressor_out_189 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_189 ) ) ;
and ( 
    .Z ( edt_scan_in_107 ) ,
    .I0 ( edt_decompressor_out_107 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_107 ) ) ;
and ( 
    .Z ( edt_scan_in_192 ) ,
    .I0 ( edt_decompressor_out_192 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_192 ) ) ;
and ( 
    .Z ( edt_scan_in_106 ) ,
    .I0 ( edt_decompressor_out_106 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_106 ) ) ;
and ( 
    .Z ( edt_scan_in_193 ) ,
    .I0 ( edt_decompressor_out_193 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_193 ) ) ;
and ( 
    .Z ( edt_scan_in_110 ) ,
    .I0 ( edt_decompressor_out_110 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_110 ) ) ;
and ( 
    .Z ( edt_scan_in_109 ) ,
    .I0 ( edt_decompressor_out_109 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_109 ) ) ;
and ( 
    .Z ( edt_scan_in_103 ) ,
    .I0 ( edt_decompressor_out_103 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_103 ) ) ;
and ( 
    .Z ( edt_scan_in_102 ) ,
    .I0 ( edt_decompressor_out_102 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_102 ) ) ;
and ( 
    .Z ( edt_scan_in_105 ) ,
    .I0 ( edt_decompressor_out_105 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_105 ) ) ;
and ( 
    .Z ( edt_scan_in_104 ) ,
    .I0 ( edt_decompressor_out_104 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_104 ) ) ;
and ( 
    .Z ( edt_scan_in_433 ) ,
    .I0 ( edt_decompressor_out_433 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_433 ) ) ;
and ( 
    .Z ( edt_scan_in_434 ) ,
    .I0 ( edt_decompressor_out_434 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_434 ) ) ;
and ( 
    .Z ( edt_scan_in_711 ) ,
    .I0 ( edt_decompressor_out_711 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_711 ) ) ;
and ( 
    .Z ( edt_scan_in_435 ) ,
    .I0 ( edt_decompressor_out_435 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_435 ) ) ;
and ( 
    .Z ( edt_scan_in_710 ) ,
    .I0 ( edt_decompressor_out_710 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_710 ) ) ;
and ( 
    .Z ( edt_scan_in_436 ) ,
    .I0 ( edt_decompressor_out_436 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_436 ) ) ;
and ( 
    .Z ( edt_scan_in_709 ) ,
    .I0 ( edt_decompressor_out_709 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_709 ) ) ;
and ( 
    .Z ( edt_scan_in_112 ) ,
    .I0 ( edt_decompressor_out_112 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_112 ) ) ;
and ( 
    .Z ( edt_scan_in_428 ) ,
    .I0 ( edt_decompressor_out_428 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_428 ) ) ;
and ( 
    .Z ( edt_scan_in_708 ) ,
    .I0 ( edt_decompressor_out_708 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_708 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_4 ) ) ;
and ( 
    .Z ( edt_scan_in_429 ) ,
    .I0 ( edt_decompressor_out_429 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_429 ) ) ;
and ( 
    .Z ( edt_scan_in_707 ) ,
    .I0 ( edt_decompressor_out_707 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_707 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N164 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_5.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N121 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1111 ) ) ;
and ( 
    .Z ( edt_scan_in_430 ) ,
    .I0 ( edt_decompressor_out_430 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_430 ) ) ;
and ( 
    .Z ( edt_scan_in_706 ) ,
    .I0 ( edt_decompressor_out_706 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_706 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1111 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_1 ) ) ;
and ( 
    .Z ( edt_scan_in_431 ) ,
    .I0 ( edt_decompressor_out_431 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_431 ) ) ;
and ( 
    .Z ( edt_scan_in_705 ) ,
    .I0 ( edt_decompressor_out_705 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_705 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N166 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_7 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N15 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n136 ) ) ;
and ( 
    .Z ( edt_scan_in_704 ) ,
    .I0 ( edt_decompressor_out_704 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_704 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n136 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_1 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N14 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n138 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n138 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_6 ) ) ;
and ( 
    .Z ( edt_scan_in_229 ) ,
    .I0 ( edt_decompressor_out_229 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_229 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N90 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n490 ) ) ;
and ( 
    .Z ( edt_scan_in_230 ) ,
    .I0 ( edt_decompressor_out_230 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_230 ) ) ;
and ( 
    .Z ( edt_scan_in_227 ) ,
    .I0 ( edt_decompressor_out_227 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_227 ) ) ;
and ( 
    .Z ( edt_scan_in_228 ) ,
    .I0 ( edt_decompressor_out_228 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_228 ) ) ;
and ( 
    .Z ( edt_scan_in_225 ) ,
    .I0 ( edt_decompressor_out_225 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_225 ) ) ;
and ( 
    .Z ( edt_scan_in_226 ) ,
    .I0 ( edt_decompressor_out_226 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_226 ) ) ;
and ( 
    .Z ( edt_scan_in_233 ) ,
    .I0 ( edt_decompressor_out_233 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_233 ) ) ;
and ( 
    .Z ( edt_scan_in_594 ) ,
    .I0 ( edt_decompressor_out_594 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_594 ) ) ;
and ( 
    .Z ( edt_scan_in_234 ) ,
    .I0 ( edt_decompressor_out_234 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_234 ) ) ;
and ( 
    .Z ( edt_scan_in_540 ) ,
    .I0 ( edt_decompressor_out_540 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_540 ) ) ;
and ( 
    .Z ( edt_scan_in_702 ) ,
    .I0 ( edt_decompressor_out_702 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_702 ) ) ;
and ( 
    .Z ( edt_scan_in_648 ) ,
    .I0 ( edt_decompressor_out_648 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_648 ) ) ;
and ( 
    .Z ( edt_scan_in_378 ) ,
    .I0 ( edt_decompressor_out_378 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_378 ) ) ;
and ( 
    .Z ( edt_scan_in_324 ) ,
    .I0 ( edt_decompressor_out_324 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_324 ) ) ;
and ( 
    .Z ( edt_scan_in_486 ) ,
    .I0 ( edt_decompressor_out_486 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_486 ) ) ;
and ( 
    .Z ( edt_scan_in_432 ) ,
    .I0 ( edt_decompressor_out_432 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_432 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N82 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n570 ) ) ;
and ( 
    .Z ( edt_scan_in_199 ) ,
    .I0 ( edt_decompressor_out_199 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_199 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N27 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1011 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1100 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_14_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1011 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N39 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n911 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n911 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_3_7 ) ) ;
and ( 
    .Z ( edt_scan_in_117 ) ,
    .I0 ( edt_decompressor_out_117 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_117 ) ) ;
and ( 
    .Z ( edt_scan_in_203 ) ,
    .I0 ( edt_decompressor_out_203 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_203 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N25 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1030 ) ) ;
and ( 
    .Z ( edt_scan_in_118 ) ,
    .I0 ( edt_decompressor_out_118 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_118 ) ) ;
and ( 
    .Z ( edt_scan_in_202 ) ,
    .I0 ( edt_decompressor_out_202 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_202 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1030 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_0 ) ) ;
and ( 
    .Z ( edt_scan_in_120 ) ,
    .I0 ( edt_decompressor_out_120 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_120 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n812 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_1 ) ) ;
and ( 
    .Z ( edt_scan_in_113 ) ,
    .I0 ( edt_decompressor_out_113 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_113 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_2 ) ) ;
and ( 
    .Z ( edt_scan_in_114 ) ,
    .I0 ( edt_decompressor_out_114 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_114 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N194 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_3.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_3 ) ) ;
and ( 
    .Z ( edt_scan_in_115 ) ,
    .I0 ( edt_decompressor_out_115 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_115 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_4 ) ) ;
and ( 
    .Z ( edt_scan_in_116 ) ,
    .I0 ( edt_decompressor_out_116 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_116 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_5 ) ) ;
and ( 
    .Z ( edt_scan_in_444 ) ,
    .I0 ( edt_decompressor_out_444 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_444 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_8_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_8_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_6 ) ) ;
and ( 
    .Z ( edt_scan_in_443 ) ,
    .I0 ( edt_decompressor_out_443 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_443 ) ) ;
and ( 
    .Z ( edt_scan_in_699 ) ,
    .I0 ( edt_decompressor_out_699 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_699 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N198 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_8_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_8_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_8_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_8_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_8_7 ) ) ;
and ( 
    .Z ( edt_scan_in_446 ) ,
    .I0 ( edt_decompressor_out_446 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_446 ) ) ;
and ( 
    .Z ( edt_scan_in_700 ) ,
    .I0 ( edt_decompressor_out_700 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_700 ) ) ;
and ( 
    .Z ( edt_scan_in_445 ) ,
    .I0 ( edt_decompressor_out_445 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_445 ) ) ;
and ( 
    .Z ( edt_scan_in_697 ) ,
    .I0 ( edt_decompressor_out_697 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_697 ) ) ;
and ( 
    .Z ( edt_scan_in_121 ) ,
    .I0 ( edt_decompressor_out_121 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_121 ) ) ;
and ( 
    .Z ( edt_scan_in_440 ) ,
    .I0 ( edt_decompressor_out_440 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_440 ) ) ;
and ( 
    .Z ( edt_scan_in_698 ) ,
    .I0 ( edt_decompressor_out_698 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_698 ) ) ;
and ( 
    .Z ( edt_scan_in_122 ) ,
    .I0 ( edt_decompressor_out_122 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_122 ) ) ;
and ( 
    .Z ( edt_scan_in_439 ) ,
    .I0 ( edt_decompressor_out_439 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_439 ) ) ;
and ( 
    .Z ( edt_scan_in_695 ) ,
    .I0 ( edt_decompressor_out_695 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_695 ) ) ;
and ( 
    .Z ( edt_scan_in_442 ) ,
    .I0 ( edt_decompressor_out_442 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_442 ) ) ;
and ( 
    .Z ( edt_scan_in_696 ) ,
    .I0 ( edt_decompressor_out_696 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_696 ) ) ;
and ( 
    .Z ( edt_scan_in_441 ) ,
    .I0 ( edt_decompressor_out_441 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_441 ) ) ;
and ( 
    .Z ( edt_scan_in_693 ) ,
    .I0 ( edt_decompressor_out_693 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_693 ) ) ;
and ( 
    .Z ( edt_scan_in_694 ) ,
    .I0 ( edt_decompressor_out_694 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_694 ) ) ;
and ( 
    .Z ( edt_scan_in_448 ) ,
    .I0 ( edt_decompressor_out_448 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_448 ) ) ;
and ( 
    .Z ( edt_scan_in_447 ) ,
    .I0 ( edt_decompressor_out_447 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_447 ) ) ;
and ( 
    .Z ( edt_scan_in_164 ) ,
    .I0 ( edt_decompressor_out_164 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_164 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n133 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_3 ) ) ;
and ( 
    .Z ( edt_scan_in_701 ) ,
    .I0 ( edt_decompressor_out_701 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_701 ) ) ;
and ( 
    .Z ( edt_scan_in_165 ) ,
    .I0 ( edt_decompressor_out_165 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_165 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N19 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n133 ) ) ;
and ( 
    .Z ( edt_scan_in_703 ) ,
    .I0 ( edt_decompressor_out_703 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_703 ) ) ;
and ( 
    .Z ( edt_scan_in_166 ) ,
    .I0 ( edt_decompressor_out_166 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_166 ) ) ;
and ( 
    .Z ( edt_scan_in_167 ) ,
    .I0 ( edt_decompressor_out_167 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_167 ) ) ;
and ( 
    .Z ( edt_scan_in_168 ) ,
    .I0 ( edt_decompressor_out_168 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_168 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n135 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_1 ) ) ;
and ( 
    .Z ( edt_scan_in_169 ) ,
    .I0 ( edt_decompressor_out_169 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_169 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N17 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n135 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n134 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_2 ) ) ;
and ( 
    .Z ( edt_scan_in_171 ) ,
    .I0 ( edt_decompressor_out_171 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_171 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N18 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n134 ) ) ;
and ( 
    .Z ( edt_scan_in_172 ) ,
    .I0 ( edt_decompressor_out_172 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_172 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n990 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_5 ) ) ;
and ( 
    .Z ( edt_scan_in_173 ) ,
    .I0 ( edt_decompressor_out_173 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_173 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N29 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n990 ) ) ;
and ( 
    .Z ( edt_scan_in_85 ) ,
    .I0 ( edt_decompressor_out_85 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_85 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n980 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_6 ) ) ;
and ( 
    .Z ( edt_scan_in_84 ) ,
    .I0 ( edt_decompressor_out_84 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_84 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N30 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n980 ) ) ;
and ( 
    .Z ( edt_scan_in_82 ) ,
    .I0 ( edt_decompressor_out_82 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_82 ) ) ;
and ( 
    .Z ( edt_scan_in_89 ) ,
    .I0 ( edt_decompressor_out_89 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_89 ) ) ;
and ( 
    .Z ( edt_scan_in_88 ) ,
    .I0 ( edt_decompressor_out_88 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_88 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N115 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1160 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N68 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_4.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1160 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N69 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_5.QT ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N111 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1200 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N70 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_6.QT ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1240 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1200 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_12_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N71 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_7_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_7_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_7_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_7_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_7_reg_7.QT ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N107 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1240 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N113 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1180 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1180 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_1 ) ) ;
and ( 
    .Z ( edt_scan_in_220 ) ,
    .I0 ( edt_decompressor_out_220 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_220 ) ) ;
and ( 
    .Z ( edt_scan_in_219 ) ,
    .I0 ( edt_decompressor_out_219 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_219 ) ) ;
and ( 
    .Z ( edt_scan_in_222 ) ,
    .I0 ( edt_decompressor_out_222 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_222 ) ) ;
and ( 
    .Z ( edt_scan_in_221 ) ,
    .I0 ( edt_decompressor_out_221 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_221 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N116 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1150 ) ) ;
and ( 
    .Z ( edt_scan_in_215 ) ,
    .I0 ( edt_decompressor_out_215 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_215 ) ) ;
and ( 
    .Z ( edt_scan_in_409 ) ,
    .I0 ( edt_decompressor_out_409 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_409 ) ) ;
and ( 
    .Z ( edt_scan_in_686 ) ,
    .I0 ( edt_decompressor_out_686 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_686 ) ) ;
and ( 
    .Z ( edt_scan_in_685 ) ,
    .I0 ( edt_decompressor_out_685 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_685 ) ) ;
and ( 
    .Z ( edt_scan_in_332 ) ,
    .I0 ( edt_decompressor_out_332 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_332 ) ) ;
and ( 
    .Z ( edt_scan_in_331 ) ,
    .I0 ( edt_decompressor_out_331 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_331 ) ) ;
and ( 
    .Z ( edt_scan_in_334 ) ,
    .I0 ( edt_decompressor_out_334 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_334 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N22 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_6.QT ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N190 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_7 ) ) ;
and ( 
    .Z ( edt_scan_in_333 ) ,
    .I0 ( edt_decompressor_out_333 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_333 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N23 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_692 ) ,
    .I0 ( edt_decompressor_out_692 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_692 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_6 ) ) ;
and ( 
    .Z ( edt_scan_in_640 ) ,
    .I0 ( edt_decompressor_out_640 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_640 ) ) ;
and ( 
    .Z ( edt_scan_in_328 ) ,
    .I0 ( edt_decompressor_out_328 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_328 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_416 ) ,
    .I0 ( edt_decompressor_out_416 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_416 ) ) ;
and ( 
    .Z ( edt_scan_in_691 ) ,
    .I0 ( edt_decompressor_out_691 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_691 ) ) ;
and ( 
    .Z ( edt_scan_in_175 ) ,
    .I0 ( edt_decompressor_out_175 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_175 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_5 ) ) ;
and ( 
    .Z ( edt_scan_in_641 ) ,
    .I0 ( edt_decompressor_out_641 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_641 ) ) ;
and ( 
    .Z ( edt_scan_in_327 ) ,
    .I0 ( edt_decompressor_out_327 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_327 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N21 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29284 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_417 ) ,
    .I0 ( edt_decompressor_out_417 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_417 ) ) ;
and ( 
    .Z ( edt_scan_in_174 ) ,
    .I0 ( edt_decompressor_out_174 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_174 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n1112 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_4 ) ) ;
and ( 
    .Z ( edt_scan_in_330 ) ,
    .I0 ( edt_decompressor_out_330 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_330 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_177 ) ,
    .I0 ( edt_decompressor_out_177 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_177 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_3 ) ) ;
and ( 
    .Z ( edt_scan_in_329 ) ,
    .I0 ( edt_decompressor_out_329 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_329 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N19 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_176 ) ,
    .I0 ( edt_decompressor_out_176 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_176 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N16 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_179 ) ,
    .I0 ( edt_decompressor_out_179 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_179 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_1_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_1_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_1_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_1_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_1_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_178 ) ,
    .I0 ( edt_decompressor_out_178 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_178 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_7_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_7_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_7_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_7_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_7_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_7_0 ) ) ;
and ( 
    .Z ( edt_scan_in_634 ) ,
    .I0 ( edt_decompressor_out_634 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_634 ) ) ;
and ( 
    .Z ( edt_scan_in_181 ) ,
    .I0 ( edt_decompressor_out_181 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_181 ) ) ;
and ( 
    .Z ( edt_scan_in_635 ) ,
    .I0 ( edt_decompressor_out_635 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_635 ) ) ;
and ( 
    .Z ( edt_scan_in_180 ) ,
    .I0 ( edt_decompressor_out_180 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_180 ) ) ;
and ( 
    .Z ( edt_scan_in_632 ) ,
    .I0 ( edt_decompressor_out_632 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_632 ) ) ;
and ( 
    .Z ( edt_scan_in_336 ) ,
    .I0 ( edt_decompressor_out_336 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_336 ) ) ;
and ( 
    .Z ( edt_scan_in_183 ) ,
    .I0 ( edt_decompressor_out_183 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_183 ) ) ;
and ( 
    .Z ( edt_scan_in_633 ) ,
    .I0 ( edt_decompressor_out_633 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_633 ) ) ;
and ( 
    .Z ( edt_scan_in_182 ) ,
    .I0 ( edt_decompressor_out_182 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_182 ) ) ;
and ( 
    .Z ( edt_scan_in_638 ) ,
    .I0 ( edt_decompressor_out_638 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_638 ) ) ;
and ( 
    .Z ( edt_scan_in_94 ) ,
    .I0 ( edt_decompressor_out_94 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_94 ) ) ;
and ( 
    .Z ( edt_scan_in_639 ) ,
    .I0 ( edt_decompressor_out_639 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_639 ) ) ;
and ( 
    .Z ( edt_scan_in_95 ) ,
    .I0 ( edt_decompressor_out_95 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_95 ) ) ;
and ( 
    .Z ( edt_scan_in_636 ) ,
    .I0 ( edt_decompressor_out_636 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_636 ) ) ;
and ( 
    .Z ( edt_scan_in_92 ) ,
    .I0 ( edt_decompressor_out_92 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_92 ) ) ;
and ( 
    .Z ( edt_scan_in_637 ) ,
    .I0 ( edt_decompressor_out_637 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_637 ) ) ;
and ( 
    .Z ( edt_scan_in_93 ) ,
    .I0 ( edt_decompressor_out_93 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_93 ) ) ;
and ( 
    .Z ( edt_scan_in_98 ) ,
    .I0 ( edt_decompressor_out_98 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_98 ) ) ;
and ( 
    .Z ( edt_scan_in_99 ) ,
    .I0 ( edt_decompressor_out_99 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_99 ) ) ;
and ( 
    .Z ( edt_scan_in_96 ) ,
    .I0 ( edt_decompressor_out_96 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_96 ) ) ;
and ( 
    .Z ( edt_scan_in_97 ) ,
    .I0 ( edt_decompressor_out_97 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_97 ) ) ;
and ( 
    .Z ( edt_scan_in_425 ) ,
    .I0 ( edt_decompressor_out_425 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_425 ) ) ;
and ( 
    .Z ( edt_scan_in_424 ) ,
    .I0 ( edt_decompressor_out_424 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_424 ) ) ;
and ( 
    .Z ( edt_scan_in_677 ) ,
    .I0 ( edt_decompressor_out_677 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_677 ) ) ;
and ( 
    .Z ( edt_scan_in_100 ) ,
    .I0 ( edt_decompressor_out_100 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_100 ) ) ;
and ( 
    .Z ( edt_scan_in_423 ) ,
    .I0 ( edt_decompressor_out_423 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_423 ) ) ;
and ( 
    .Z ( edt_scan_in_678 ) ,
    .I0 ( edt_decompressor_out_678 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_678 ) ) ;
and ( 
    .Z ( edt_scan_in_101 ) ,
    .I0 ( edt_decompressor_out_101 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_101 ) ) ;
and ( 
    .Z ( edt_scan_in_422 ) ,
    .I0 ( edt_decompressor_out_422 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_422 ) ) ;
and ( 
    .Z ( edt_scan_in_679 ) ,
    .I0 ( edt_decompressor_out_679 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_679 ) ) ;
and ( 
    .Z ( edt_scan_in_421 ) ,
    .I0 ( edt_decompressor_out_421 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_421 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n1110 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( edt_scan_in_680 ) ,
    .I0 ( edt_decompressor_out_680 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_680 ) ) ;
and ( 
    .Z ( edt_scan_in_420 ) ,
    .I0 ( edt_decompressor_out_420 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_420 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n910 ) ,
    .I0 ( n40 ) ,
    .I1 ( constant_shift_controller_i.n271 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n1012 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_4_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_4_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_4_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_4_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_4_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_4_3 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N13 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n139 ) ) ;
and ( 
    .Z ( edt_scan_in_437 ) ,
    .I0 ( edt_decompressor_out_437 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_437 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n139 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_5 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N28 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1000 ) ) ;
and ( 
    .Z ( edt_scan_in_713 ) ,
    .I0 ( edt_decompressor_out_713 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_713 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1000 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_4 ) ) ;
and ( 
    .Z ( edt_scan_in_712 ) ,
    .I0 ( edt_decompressor_out_712 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_712 ) ) ;
and ( 
    .Z ( edt_scan_in_195 ) ,
    .I0 ( edt_decompressor_out_195 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_195 ) ) ;
and ( 
    .Z ( edt_scan_in_194 ) ,
    .I0 ( edt_decompressor_out_194 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_194 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N26 ) ,
    .I0 ( constant_shift_controller_i.n261 ) ,
    .I1 ( constant_shift_controller_i.n1020 ) ) ;
and ( 
    .Z ( edt_scan_in_200 ) ,
    .I0 ( edt_decompressor_out_200 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_200 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n1020 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_2 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.N122 ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( constant_shift_controller_i.n1100 ) ) ;
and ( 
    .Z ( edt_scan_in_343 ) ,
    .I0 ( edt_decompressor_out_343 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_343 ) ) ;
and ( 
    .Z ( edt_scan_in_344 ) ,
    .I0 ( edt_decompressor_out_344 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_344 ) ) ;
and ( 
    .Z ( edt_scan_in_681 ) ,
    .I0 ( edt_decompressor_out_681 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_681 ) ) ;
and ( 
    .Z ( edt_scan_in_652 ) ,
    .I0 ( edt_decompressor_out_652 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_652 ) ) ;
and ( 
    .Z ( edt_scan_in_337 ) ,
    .I0 ( edt_decompressor_out_337 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_337 ) ) ;
and ( 
    .Z ( edt_scan_in_427 ) ,
    .I0 ( edt_decompressor_out_427 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_427 ) ) ;
and ( 
    .Z ( edt_scan_in_682 ) ,
    .I0 ( edt_decompressor_out_682 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_682 ) ) ;
and ( 
    .Z ( edt_scan_in_651 ) ,
    .I0 ( edt_decompressor_out_651 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_651 ) ) ;
and ( 
    .Z ( edt_scan_in_338 ) ,
    .I0 ( edt_decompressor_out_338 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_338 ) ) ;
and ( 
    .Z ( edt_scan_in_426 ) ,
    .I0 ( edt_decompressor_out_426 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_426 ) ) ;
and ( 
    .Z ( edt_scan_in_340 ) ,
    .I0 ( edt_decompressor_out_340 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_340 ) ) ;
and ( 
    .Z ( edt_scan_in_795 ) ,
    .I0 ( edt_decompressor_out_795 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_795 ) ) ;
and ( 
    .Z ( edt_scan_in_645 ) ,
    .I0 ( edt_decompressor_out_645 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_645 ) ) ;
and ( 
    .Z ( edt_scan_in_644 ) ,
    .I0 ( edt_decompressor_out_644 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_644 ) ) ;
and ( 
    .Z ( edt_scan_in_643 ) ,
    .I0 ( edt_decompressor_out_643 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_643 ) ) ;
and ( 
    .Z ( edt_scan_in_345 ) ,
    .I0 ( edt_decompressor_out_345 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_345 ) ) ;
and ( 
    .Z ( edt_scan_in_642 ) ,
    .I0 ( edt_decompressor_out_642 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_642 ) ) ;
and ( 
    .Z ( edt_scan_in_346 ) ,
    .I0 ( edt_decompressor_out_346 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_346 ) ) ;
and ( 
    .Z ( edt_scan_in_650 ) ,
    .I0 ( edt_decompressor_out_650 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_650 ) ) ;
and ( 
    .Z ( edt_scan_in_63 ) ,
    .I0 ( edt_decompressor_out_63 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_63 ) ) ;
and ( 
    .Z ( edt_scan_in_649 ) ,
    .I0 ( edt_decompressor_out_649 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_649 ) ) ;
and ( 
    .Z ( edt_scan_in_62 ) ,
    .I0 ( edt_decompressor_out_62 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_62 ) ) ;
and ( 
    .Z ( edt_scan_in_647 ) ,
    .I0 ( edt_decompressor_out_647 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_647 ) ) ;
and ( 
    .Z ( edt_scan_in_65 ) ,
    .I0 ( edt_decompressor_out_65 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_65 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n501 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_1 ) ) ;
and ( 
    .Z ( edt_scan_in_646 ) ,
    .I0 ( edt_decompressor_out_646 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_646 ) ) ;
and ( 
    .Z ( edt_scan_in_64 ) ,
    .I0 ( edt_decompressor_out_64 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_64 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_0 ) ) ;
and ( 
    .Z ( edt_scan_in_67 ) ,
    .I0 ( edt_decompressor_out_67 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_67 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_3 ) ) ;
and ( 
    .Z ( edt_scan_in_66 ) ,
    .I0 ( edt_decompressor_out_66 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_66 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_2 ) ) ;
and ( 
    .Z ( edt_scan_in_69 ) ,
    .I0 ( edt_decompressor_out_69 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_69 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_5 ) ) ;
and ( 
    .Z ( edt_scan_in_68 ) ,
    .I0 ( edt_decompressor_out_68 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_68 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_4 ) ) ;
and ( 
    .Z ( edt_scan_in_71 ) ,
    .I0 ( edt_decompressor_out_71 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_71 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N142 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_7 ) ) ;
and ( 
    .Z ( edt_scan_in_70 ) ,
    .I0 ( edt_decompressor_out_70 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_70 ) ) ;
and ( 
    .Z ( edt_scan_in_388 ) ,
    .I0 ( edt_decompressor_out_388 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_388 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.DI_ ) ,
    .IN ( edt_update_hfs_netlink_29285 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_1_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_1_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_1_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_1_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_1_6 ) ) ;
and ( 
    .Z ( edt_scan_in_747 ) ,
    .I0 ( edt_decompressor_out_747 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_747 ) ) ;
and ( 
    .Z ( edt_scan_in_389 ) ,
    .I0 ( edt_decompressor_out_389 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_389 ) ) ;
and ( 
    .Z ( edt_scan_in_746 ) ,
    .I0 ( edt_decompressor_out_746 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_746 ) ) ;
and ( 
    .Z ( edt_scan_in_390 ) ,
    .I0 ( edt_decompressor_out_390 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_390 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U36.AB ) ,
    .I0 ( constant_shift_controller_i.n330 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U36.CD ) ,
    .I0 ( edt_channels_in_13 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U36.ZN ) ,
    .I0 ( constant_shift_controller_i.U36.AB ) ,
    .I1 ( constant_shift_controller_i.U36.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N238 ) ,
    .IN ( constant_shift_controller_i.U36.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_745 ) ,
    .I0 ( edt_decompressor_out_745 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_745 ) ) ;
and ( 
    .Z ( edt_scan_in_391 ) ,
    .I0 ( edt_decompressor_out_391 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_391 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U37.AB ) ,
    .I0 ( edt_channels_in_6 ) ,
    .I1 ( constant_shift_controller_i.n1 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U37.CD ) ,
    .I0 ( constant_shift_controller_i.n1400 ) ,
    .I1 ( constant_shift_controller_i.n4 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U37.ZN ) ,
    .I0 ( constant_shift_controller_i.U37.AB ) ,
    .I1 ( constant_shift_controller_i.U37.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N224 ) ,
    .IN ( constant_shift_controller_i.U37.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_744 ) ,
    .I0 ( edt_decompressor_out_744 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_744 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N103 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_7 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_7.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_7.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_7.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_7.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_7.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_7.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_7.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_7.QT ) ) ;
and ( 
    .Z ( edt_scan_in_392 ) ,
    .I0 ( edt_decompressor_out_392 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_392 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U34.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_11 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U34.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n350 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U34.ZN ) ,
    .I0 ( constant_shift_controller_i.U34.AB ) ,
    .I1 ( constant_shift_controller_i.U34.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_11 ) ,
    .IN ( constant_shift_controller_i.U34.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_751 ) ,
    .I0 ( edt_decompressor_out_751 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_751 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.DI_ ) ,
    .IN ( constant_shift_controller_i.N102 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_6 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_6.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_6.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_6.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_6.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_6.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_6.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_6.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_6.QT ) ) ;
and ( 
    .Z ( edt_scan_in_393 ) ,
    .I0 ( edt_decompressor_out_393 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_393 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U35.AB ) ,
    .I0 ( constant_shift_controller_i.n310 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U35.CD ) ,
    .I0 ( edt_channels_in_14 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U35.ZN ) ,
    .I0 ( constant_shift_controller_i.U35.AB ) ,
    .I1 ( constant_shift_controller_i.U35.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N245 ) ,
    .IN ( constant_shift_controller_i.U35.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_750 ) ,
    .I0 ( edt_decompressor_out_750 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_750 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.DI_ ) ,
    .IN ( constant_shift_controller_i.N101 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_5 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_5.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_5.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_5.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_5.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_5.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_5.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_5.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_5.QT ) ) ;
and ( 
    .Z ( edt_scan_in_394 ) ,
    .I0 ( edt_decompressor_out_394 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_394 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U32.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_7 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U32.CD ) ,
    .I0 ( constant_shift_controller_i.n280 ) ,
    .I1 ( constant_shift_controller_i.n810 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U32.ZN ) ,
    .I0 ( constant_shift_controller_i.U32.AB ) ,
    .I1 ( constant_shift_controller_i.U32.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_7 ) ,
    .IN ( constant_shift_controller_i.U32.ZN ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.DI_ ) ,
    .IN ( constant_shift_controller_i.N100 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_4 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_4.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_VL_LSI_MUX21_26791.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_4.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_4.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_10 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_4.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_4.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_8 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_9 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_4.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_4.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_4.QT ) ) ;
and ( 
    .Z ( edt_scan_in_395 ) ,
    .I0 ( edt_decompressor_out_395 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_395 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U33.AB ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_9 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U33.CD ) ,
    .I0 ( constant_shift_controller_i.n3 ) ,
    .I1 ( constant_shift_controller_i.n280 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U33.ZN ) ,
    .I0 ( constant_shift_controller_i.U33.AB ) ,
    .I1 ( constant_shift_controller_i.U33.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_constant_shift_control_9 ) ,
    .IN ( constant_shift_controller_i.U33.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_748 ) ,
    .I0 ( edt_decompressor_out_748 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_748 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.DI_ ) ,
    .IN ( constant_shift_controller_i.N99 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_3 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_3.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_3.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_3.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_3.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_3.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_3.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_3.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_3.QT ) ) ;
and ( 
    .Z ( edt_scan_in_396 ) ,
    .I0 ( edt_decompressor_out_396 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_396 ) ) ;
and ( 
    .Z ( edt_scan_in_313 ) ,
    .I0 ( edt_decompressor_out_313 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_313 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.DI_ ) ,
    .IN ( constant_shift_controller_i.N98 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_2 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_2.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_2.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_2.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_2.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_2.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_2.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_2.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_2.QT ) ) ;
and ( 
    .Z ( edt_scan_in_397 ) ,
    .I0 ( edt_decompressor_out_397 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_397 ) ) ;
and ( 
    .Z ( edt_scan_in_312 ) ,
    .I0 ( edt_decompressor_out_312 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_312 ) ) ;
and ( 
    .Z ( edt_scan_in_789 ) ,
    .I0 ( edt_decompressor_out_789 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_789 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.DI_ ) ,
    .IN ( constant_shift_controller_i.N97 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_1 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_1.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_1.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_1.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_1.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_1.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_1.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_1.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_1.QT ) ) ;
and ( 
    .Z ( edt_scan_in_753 ) ,
    .I0 ( edt_decompressor_out_753 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_753 ) ) ;
and ( 
    .Z ( edt_scan_in_87 ) ,
    .I0 ( edt_decompressor_out_87 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_87 ) ) ;
and ( 
    .Z ( edt_scan_in_86 ) ,
    .I0 ( edt_decompressor_out_86 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_86 ) ) ;
and ( 
    .Z ( edt_scan_in_414 ) ,
    .I0 ( edt_decompressor_out_414 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_414 ) ) ;
and ( 
    .Z ( edt_scan_in_415 ) ,
    .I0 ( edt_decompressor_out_415 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_415 ) ) ;
and ( 
    .Z ( edt_scan_in_688 ) ,
    .I0 ( edt_decompressor_out_688 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_688 ) ) ;
and ( 
    .Z ( edt_scan_in_91 ) ,
    .I0 ( edt_decompressor_out_91 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_91 ) ) ;
and ( 
    .Z ( edt_scan_in_412 ) ,
    .I0 ( edt_decompressor_out_412 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_412 ) ) ;
and ( 
    .Z ( edt_scan_in_687 ) ,
    .I0 ( edt_decompressor_out_687 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_687 ) ) ;
and ( 
    .Z ( edt_scan_in_90 ) ,
    .I0 ( edt_decompressor_out_90 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_90 ) ) ;
and ( 
    .Z ( edt_scan_in_413 ) ,
    .I0 ( edt_decompressor_out_413 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_413 ) ) ;
and ( 
    .Z ( edt_scan_in_690 ) ,
    .I0 ( edt_decompressor_out_690 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_690 ) ) ;
and ( 
    .Z ( edt_scan_in_410 ) ,
    .I0 ( edt_decompressor_out_410 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_410 ) ) ;
and ( 
    .Z ( edt_scan_in_689 ) ,
    .I0 ( edt_decompressor_out_689 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_689 ) ) ;
and ( 
    .Z ( edt_scan_in_411 ) ,
    .I0 ( edt_decompressor_out_411 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_411 ) ) ;
and ( 
    .Z ( edt_scan_in_684 ) ,
    .I0 ( edt_decompressor_out_684 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_684 ) ) ;
and ( 
    .Z ( edt_scan_in_408 ) ,
    .I0 ( edt_decompressor_out_408 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_408 ) ) ;
and ( 
    .Z ( edt_scan_in_683 ) ,
    .I0 ( edt_decompressor_out_683 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_683 ) ) ;
and ( 
    .Z ( edt_scan_in_792 ) ,
    .I0 ( edt_decompressor_out_792 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_792 ) ) ;
and ( 
    .Z ( edt_scan_in_308 ) ,
    .I0 ( edt_decompressor_out_308 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_308 ) ) ;
and ( 
    .Z ( edt_scan_in_785 ) ,
    .I0 ( edt_decompressor_out_785 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_785 ) ) ;
and ( 
    .Z ( edt_scan_in_307 ) ,
    .I0 ( edt_decompressor_out_307 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_307 ) ) ;
and ( 
    .Z ( edt_scan_in_786 ) ,
    .I0 ( edt_decompressor_out_786 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_786 ) ) ;
and ( 
    .Z ( edt_scan_in_306 ) ,
    .I0 ( edt_decompressor_out_306 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_306 ) ) ;
and ( 
    .Z ( edt_scan_in_787 ) ,
    .I0 ( edt_decompressor_out_787 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_787 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U38.AB ) ,
    .I0 ( constant_shift_controller_i.n350 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U38.CD ) ,
    .I0 ( edt_channels_in_12 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U38.ZN ) ,
    .I0 ( constant_shift_controller_i.U38.AB ) ,
    .I1 ( constant_shift_controller_i.U38.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N230 ) ,
    .IN ( constant_shift_controller_i.U38.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_788 ) ,
    .I0 ( edt_decompressor_out_788 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_788 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U39.AB ) ,
    .I0 ( constant_shift_controller_i.n370 ) ,
    .I1 ( constant_shift_controller_i.n1040 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.U39.CD ) ,
    .I0 ( edt_channels_in_11 ) ,
    .I1 ( constant_shift_controller_i.n1050 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.U39.ZN ) ,
    .I0 ( constant_shift_controller_i.U39.AB ) ,
    .I1 ( constant_shift_controller_i.U39.CD ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.N222 ) ,
    .IN ( constant_shift_controller_i.U39.ZN ) ) ;
and ( 
    .Z ( edt_scan_in_612 ) ,
    .I0 ( edt_decompressor_out_612 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_612 ) ) ;
and ( 
    .Z ( edt_scan_in_613 ) ,
    .I0 ( edt_decompressor_out_613 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_613 ) ) ;
and ( 
    .Z ( edt_scan_in_614 ) ,
    .I0 ( edt_decompressor_out_614 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_614 ) ) ;
and ( 
    .Z ( edt_scan_in_615 ) ,
    .I0 ( edt_decompressor_out_615 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_615 ) ) ;
and ( 
    .Z ( edt_scan_in_793 ) ,
    .I0 ( edt_decompressor_out_793 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_793 ) ) ;
and ( 
    .Z ( edt_scan_in_539 ) ,
    .I0 ( edt_decompressor_out_539 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_539 ) ) ;
and ( 
    .Z ( edt_scan_in_616 ) ,
    .I0 ( edt_decompressor_out_616 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_616 ) ) ;
and ( 
    .Z ( edt_scan_in_315 ) ,
    .I0 ( edt_decompressor_out_315 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_315 ) ) ;
and ( 
    .Z ( edt_scan_in_794 ) ,
    .I0 ( edt_decompressor_out_794 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_794 ) ) ;
and ( 
    .Z ( edt_scan_in_72 ) ,
    .I0 ( edt_decompressor_out_72 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_72 ) ) ;
and ( 
    .Z ( edt_scan_in_538 ) ,
    .I0 ( edt_decompressor_out_538 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_538 ) ) ;
and ( 
    .Z ( edt_scan_in_617 ) ,
    .I0 ( edt_decompressor_out_617 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_617 ) ) ;
and ( 
    .Z ( edt_scan_in_314 ) ,
    .I0 ( edt_decompressor_out_314 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_314 ) ) ;
and ( 
    .Z ( edt_scan_in_73 ) ,
    .I0 ( edt_decompressor_out_73 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_73 ) ) ;
and ( 
    .Z ( edt_scan_in_74 ) ,
    .I0 ( edt_decompressor_out_74 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_74 ) ) ;
and ( 
    .Z ( edt_scan_in_75 ) ,
    .I0 ( edt_decompressor_out_75 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_75 ) ) ;
and ( 
    .Z ( edt_scan_in_76 ) ,
    .I0 ( edt_decompressor_out_76 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_76 ) ) ;
and ( 
    .Z ( edt_scan_in_77 ) ,
    .I0 ( edt_decompressor_out_77 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_77 ) ) ;
and ( 
    .Z ( edt_scan_in_533 ) ,
    .I0 ( edt_decompressor_out_533 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_533 ) ) ;
and ( 
    .Z ( edt_scan_in_78 ) ,
    .I0 ( edt_decompressor_out_78 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_78 ) ) ;
and ( 
    .Z ( edt_scan_in_532 ) ,
    .I0 ( edt_decompressor_out_532 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_532 ) ) ;
and ( 
    .Z ( edt_scan_in_79 ) ,
    .I0 ( edt_decompressor_out_79 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_79 ) ) ;
and ( 
    .Z ( edt_scan_in_531 ) ,
    .I0 ( edt_decompressor_out_531 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_531 ) ) ;
and ( 
    .Z ( edt_scan_in_80 ) ,
    .I0 ( edt_decompressor_out_80 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_80 ) ) ;
and ( 
    .Z ( edt_scan_in_537 ) ,
    .I0 ( edt_decompressor_out_537 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_537 ) ) ;
and ( 
    .Z ( edt_scan_in_736 ) ,
    .I0 ( edt_decompressor_out_736 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_736 ) ) ;
and ( 
    .Z ( edt_scan_in_536 ) ,
    .I0 ( edt_decompressor_out_536 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_536 ) ) ;
and ( 
    .Z ( edt_scan_in_398 ) ,
    .I0 ( edt_decompressor_out_398 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_398 ) ) ;
and ( 
    .Z ( edt_scan_in_737 ) ,
    .I0 ( edt_decompressor_out_737 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_737 ) ) ;
and ( 
    .Z ( edt_scan_in_535 ) ,
    .I0 ( edt_decompressor_out_535 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_535 ) ) ;
and ( 
    .Z ( edt_scan_in_401 ) ,
    .I0 ( edt_decompressor_out_401 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_401 ) ) ;
and ( 
    .Z ( edt_scan_in_734 ) ,
    .I0 ( edt_decompressor_out_734 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_734 ) ) ;
and ( 
    .Z ( edt_scan_in_50 ) ,
    .I0 ( edt_decompressor_out_50 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_50 ) ) ;
and ( 
    .Z ( edt_scan_in_534 ) ,
    .I0 ( edt_decompressor_out_534 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_534 ) ) ;
and ( 
    .Z ( edt_scan_in_400 ) ,
    .I0 ( edt_decompressor_out_400 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_400 ) ) ;
and ( 
    .Z ( edt_scan_in_735 ) ,
    .I0 ( edt_decompressor_out_735 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_735 ) ) ;
and ( 
    .Z ( edt_scan_in_47 ) ,
    .I0 ( edt_decompressor_out_47 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_47 ) ) ;
and ( 
    .Z ( edt_scan_in_403 ) ,
    .I0 ( edt_decompressor_out_403 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_403 ) ) ;
and ( 
    .Z ( edt_scan_in_740 ) ,
    .I0 ( edt_decompressor_out_740 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_740 ) ) ;
and ( 
    .Z ( edt_scan_in_48 ) ,
    .I0 ( edt_decompressor_out_48 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_48 ) ) ;
and ( 
    .Z ( edt_scan_in_402 ) ,
    .I0 ( edt_decompressor_out_402 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_402 ) ) ;
and ( 
    .Z ( edt_scan_in_741 ) ,
    .I0 ( edt_decompressor_out_741 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_741 ) ) ;
and ( 
    .Z ( edt_scan_in_45 ) ,
    .I0 ( edt_decompressor_out_45 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_45 ) ) ;
and ( 
    .Z ( edt_scan_in_405 ) ,
    .I0 ( edt_decompressor_out_405 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_405 ) ) ;
and ( 
    .Z ( edt_scan_in_738 ) ,
    .I0 ( edt_decompressor_out_738 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_738 ) ) ;
and ( 
    .Z ( edt_scan_in_46 ) ,
    .I0 ( edt_decompressor_out_46 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_46 ) ) ;
and ( 
    .Z ( edt_scan_in_404 ) ,
    .I0 ( edt_decompressor_out_404 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_404 ) ) ;
and ( 
    .Z ( edt_scan_in_739 ) ,
    .I0 ( edt_decompressor_out_739 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_739 ) ) ;
and ( 
    .Z ( edt_scan_in_43 ) ,
    .I0 ( edt_decompressor_out_43 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_43 ) ) ;
and ( 
    .Z ( edt_scan_in_407 ) ,
    .I0 ( edt_decompressor_out_407 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_407 ) ) ;
and ( 
    .Z ( edt_scan_in_44 ) ,
    .I0 ( edt_decompressor_out_44 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_44 ) ) ;
and ( 
    .Z ( edt_scan_in_322 ) ,
    .I0 ( edt_decompressor_out_322 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_322 ) ) ;
and ( 
    .Z ( edt_scan_in_406 ) ,
    .I0 ( edt_decompressor_out_406 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_406 ) ) ;
and ( 
    .Z ( edt_scan_in_41 ) ,
    .I0 ( edt_decompressor_out_41 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_41 ) ) ;
and ( 
    .Z ( edt_scan_in_323 ) ,
    .I0 ( edt_decompressor_out_323 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_323 ) ) ;
and ( 
    .Z ( edt_scan_in_780 ) ,
    .I0 ( edt_decompressor_out_780 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_780 ) ) ;
and ( 
    .Z ( edt_scan_in_742 ) ,
    .I0 ( edt_decompressor_out_742 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_742 ) ) ;
and ( 
    .Z ( edt_scan_in_42 ) ,
    .I0 ( edt_decompressor_out_42 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_42 ) ) ;
and ( 
    .Z ( edt_scan_in_631 ) ,
    .I0 ( edt_decompressor_out_631 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_631 ) ) ;
and ( 
    .Z ( edt_scan_in_320 ) ,
    .I0 ( edt_decompressor_out_320 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_320 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_0.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_0.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_0.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_0.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_0.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_0 ) ) ;
and ( 
    .Z ( edt_scan_in_779 ) ,
    .I0 ( edt_decompressor_out_779 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_779 ) ) ;
and ( 
    .Z ( edt_scan_in_743 ) ,
    .I0 ( edt_decompressor_out_743 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_743 ) ) ;
and ( 
    .Z ( edt_scan_in_630 ) ,
    .I0 ( edt_decompressor_out_630 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_630 ) ) ;
and ( 
    .Z ( edt_scan_in_321 ) ,
    .I0 ( edt_decompressor_out_321 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_321 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_1.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_1.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_1.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_1.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_1.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_1.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_1 ) ) ;
and ( 
    .Z ( edt_scan_in_782 ) ,
    .I0 ( edt_decompressor_out_782 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_782 ) ) ;
and ( 
    .Z ( edt_scan_in_318 ) ,
    .I0 ( edt_decompressor_out_318 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_318 ) ) ;
and ( 
    .Z ( edt_scan_in_673 ) ,
    .I0 ( edt_decompressor_out_673 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_673 ) ) ;
and ( 
    .Z ( edt_scan_in_419 ) ,
    .I0 ( edt_decompressor_out_419 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_419 ) ) ;
and ( 
    .Z ( edt_scan_in_674 ) ,
    .I0 ( edt_decompressor_out_674 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_674 ) ) ;
and ( 
    .Z ( edt_scan_in_418 ) ,
    .I0 ( edt_decompressor_out_418 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_418 ) ) ;
and ( 
    .Z ( edt_scan_in_675 ) ,
    .I0 ( edt_decompressor_out_675 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_675 ) ) ;
and ( 
    .Z ( edt_scan_in_676 ) ,
    .I0 ( edt_decompressor_out_676 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_676 ) ) ;
and ( 
    .Z ( edt_scan_in_341 ) ,
    .I0 ( edt_decompressor_out_341 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_341 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n1 ) ,
    .I0 ( n40 ) ,
    .I1 ( n54 ) ) ;
and ( 
    .Z ( edt_scan_in_342 ) ,
    .I0 ( edt_decompressor_out_342 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_342 ) ) ;
and ( 
    .Z ( edt_scan_in_319 ) ,
    .I0 ( edt_decompressor_out_319 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_319 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_4 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_3.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_3.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_3.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_3.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_3.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_3.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_3 ) ) ;
and ( 
    .Z ( edt_scan_in_776 ) ,
    .I0 ( edt_decompressor_out_776 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_776 ) ) ;
and ( 
    .Z ( edt_scan_in_316 ) ,
    .I0 ( edt_decompressor_out_316 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_316 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.CDNI_ ) ,
    .IN ( constant_shift_controller_i.n511 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_4.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_4.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_4.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_4.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_4.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_4.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_4 ) ) ;
and ( 
    .Z ( edt_scan_in_775 ) ,
    .I0 ( edt_decompressor_out_775 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_775 ) ) ;
and ( 
    .Z ( edt_scan_in_317 ) ,
    .I0 ( edt_decompressor_out_317 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_317 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_6 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_5.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_5.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_5.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_5.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_5.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_5.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_5 ) ) ;
and ( 
    .Z ( edt_scan_in_778 ) ,
    .I0 ( edt_decompressor_out_778 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_778 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_7 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_6.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_6.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_6.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_6.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_6.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_6.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_6 ) ) ;
and ( 
    .Z ( edt_scan_in_777 ) ,
    .I0 ( edt_decompressor_out_777 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_777 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_7.DI_ ) ,
    .IN ( constant_shift_controller_i.N222 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_7.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_7.udp1.I0 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_7.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_7.DI_ ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_7 ) ) ;
and ( 
    .Z ( edt_scan_in_623 ) ,
    .I0 ( edt_decompressor_out_623 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_623 ) ) ;
and ( 
    .Z ( edt_scan_in_622 ) ,
    .I0 ( edt_decompressor_out_622 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_622 ) ) ;
and ( 
    .Z ( edt_scan_in_625 ) ,
    .I0 ( edt_decompressor_out_625 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_625 ) ) ;
and ( 
    .Z ( edt_scan_in_624 ) ,
    .I0 ( edt_decompressor_out_624 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_624 ) ) ;
and ( 
    .Z ( edt_scan_in_784 ) ,
    .I0 ( edt_decompressor_out_784 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_784 ) ) ;
and ( 
    .Z ( edt_scan_in_549 ) ,
    .I0 ( edt_decompressor_out_549 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_549 ) ) ;
and ( 
    .Z ( edt_scan_in_627 ) ,
    .I0 ( edt_decompressor_out_627 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_627 ) ) ;
and ( 
    .Z ( edt_scan_in_325 ) ,
    .I0 ( edt_decompressor_out_325 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_325 ) ) ;
and ( 
    .Z ( edt_scan_in_783 ) ,
    .I0 ( edt_decompressor_out_783 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_783 ) ) ;
and ( 
    .Z ( edt_scan_in_550 ) ,
    .I0 ( edt_decompressor_out_550 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_550 ) ) ;
and ( 
    .Z ( edt_scan_in_626 ) ,
    .I0 ( edt_decompressor_out_626 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_626 ) ) ;
and ( 
    .Z ( edt_scan_in_326 ) ,
    .I0 ( edt_decompressor_out_326 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_326 ) ) ;
and ( 
    .Z ( edt_scan_in_629 ) ,
    .I0 ( edt_decompressor_out_629 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_629 ) ) ;
and ( 
    .Z ( edt_scan_in_628 ) ,
    .I0 ( edt_decompressor_out_628 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_628 ) ) ;
and ( 
    .Z ( edt_scan_in_543 ) ,
    .I0 ( edt_decompressor_out_543 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_543 ) ) ;
and ( 
    .Z ( edt_scan_in_544 ) ,
    .I0 ( edt_decompressor_out_544 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_544 ) ) ;
and ( 
    .Z ( edt_scan_in_541 ) ,
    .I0 ( edt_decompressor_out_541 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_541 ) ) ;
and ( 
    .Z ( edt_scan_in_542 ) ,
    .I0 ( edt_decompressor_out_542 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_542 ) ) ;
and ( 
    .Z ( edt_scan_in_547 ) ,
    .I0 ( edt_decompressor_out_547 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_547 ) ) ;
and ( 
    .Z ( edt_scan_in_369 ) ,
    .I0 ( edt_decompressor_out_369 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_369 ) ) ;
and ( 
    .Z ( edt_scan_in_725 ) ,
    .I0 ( edt_decompressor_out_725 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_725 ) ) ;
and ( 
    .Z ( edt_scan_in_548 ) ,
    .I0 ( edt_decompressor_out_548 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_548 ) ) ;
and ( 
    .Z ( edt_scan_in_370 ) ,
    .I0 ( edt_decompressor_out_370 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_370 ) ) ;
and ( 
    .Z ( edt_scan_in_724 ) ,
    .I0 ( edt_decompressor_out_724 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_724 ) ) ;
and ( 
    .Z ( edt_scan_in_61 ) ,
    .I0 ( edt_decompressor_out_61 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_61 ) ) ;
and ( 
    .Z ( edt_scan_in_545 ) ,
    .I0 ( edt_decompressor_out_545 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_545 ) ) ;
and ( 
    .Z ( edt_scan_in_367 ) ,
    .I0 ( edt_decompressor_out_367 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_367 ) ) ;
and ( 
    .Z ( edt_scan_in_727 ) ,
    .I0 ( edt_decompressor_out_727 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_727 ) ) ;
and ( 
    .Z ( edt_scan_in_546 ) ,
    .I0 ( edt_decompressor_out_546 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_546 ) ) ;
and ( 
    .Z ( edt_scan_in_368 ) ,
    .I0 ( edt_decompressor_out_368 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_368 ) ) ;
and ( 
    .Z ( edt_scan_in_726 ) ,
    .I0 ( edt_decompressor_out_726 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_726 ) ) ;
and ( 
    .Z ( edt_scan_in_59 ) ,
    .I0 ( edt_decompressor_out_59 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_59 ) ) ;
and ( 
    .Z ( edt_scan_in_373 ) ,
    .I0 ( edt_decompressor_out_373 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_373 ) ) ;
and ( 
    .Z ( edt_scan_in_729 ) ,
    .I0 ( edt_decompressor_out_729 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_729 ) ) ;
and ( 
    .Z ( edt_scan_in_58 ) ,
    .I0 ( edt_decompressor_out_58 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_58 ) ) ;
and ( 
    .Z ( edt_scan_in_374 ) ,
    .I0 ( edt_decompressor_out_374 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_374 ) ) ;
and ( 
    .Z ( edt_scan_in_728 ) ,
    .I0 ( edt_decompressor_out_728 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_728 ) ) ;
and ( 
    .Z ( edt_scan_in_57 ) ,
    .I0 ( edt_decompressor_out_57 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_57 ) ) ;
and ( 
    .Z ( edt_scan_in_371 ) ,
    .I0 ( edt_decompressor_out_371 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_371 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n1050 ) ,
    .I0 ( n43 ) ,
    .I1 ( n54 ) ) ;
and ( 
    .Z ( edt_scan_in_731 ) ,
    .I0 ( edt_decompressor_out_731 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_731 ) ) ;
and ( 
    .Z ( edt_scan_in_56 ) ,
    .I0 ( edt_decompressor_out_56 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_56 ) ) ;
and ( 
    .Z ( edt_scan_in_372 ) ,
    .I0 ( edt_decompressor_out_372 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_372 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n4 ) ,
    .I0 ( n43 ) ,
    .I1 ( n54 ) ) ;
and ( 
    .Z ( edt_scan_in_730 ) ,
    .I0 ( edt_decompressor_out_730 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_730 ) ) ;
and ( 
    .Z ( edt_scan_in_55 ) ,
    .I0 ( edt_decompressor_out_55 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_55 ) ) ;
and ( 
    .Z ( edt_scan_in_733 ) ,
    .I0 ( edt_decompressor_out_733 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_733 ) ) ;
and ( 
    .Z ( edt_scan_in_53 ) ,
    .I0 ( edt_decompressor_out_53 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_53 ) ) ;
and ( 
    .Z ( edt_scan_in_287 ) ,
    .I0 ( edt_decompressor_out_287 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_287 ) ) ;
and ( 
    .Z ( edt_scan_in_732 ) ,
    .I0 ( edt_decompressor_out_732 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_732 ) ) ;
and ( 
    .Z ( edt_scan_in_52 ) ,
    .I0 ( edt_decompressor_out_52 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_52 ) ) ;
and ( 
    .Z ( edt_scan_in_286 ) ,
    .I0 ( edt_decompressor_out_286 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_286 ) ) ;
and ( 
    .Z ( edt_scan_in_375 ) ,
    .I0 ( edt_decompressor_out_375 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_375 ) ) ;
and ( 
    .Z ( edt_scan_in_51 ) ,
    .I0 ( edt_decompressor_out_51 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_51 ) ) ;
and ( 
    .Z ( edt_scan_in_289 ) ,
    .I0 ( edt_decompressor_out_289 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_289 ) ) ;
and ( 
    .Z ( edt_scan_in_376 ) ,
    .I0 ( edt_decompressor_out_376 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_376 ) ) ;
and ( 
    .Z ( edt_scan_in_288 ) ,
    .I0 ( edt_decompressor_out_288 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_288 ) ) ;
and ( 
    .Z ( edt_scan_in_291 ) ,
    .I0 ( edt_decompressor_out_291 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_291 ) ) ;
and ( 
    .Z ( edt_scan_in_290 ) ,
    .I0 ( edt_decompressor_out_290 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_290 ) ) ;
and ( 
    .Z ( edt_scan_in_293 ) ,
    .I0 ( edt_decompressor_out_293 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_293 ) ) ;
nand ( 
    .Z ( constant_shift_controller_i.n1040 ) ,
    .I0 ( n40 ) ,
    .I1 ( n54 ) ) ;
and ( 
    .Z ( edt_scan_in_292 ) ,
    .I0 ( edt_decompressor_out_292 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_292 ) ) ;
and ( 
    .Z ( edt_scan_in_600 ) ,
    .I0 ( edt_decompressor_out_600 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_600 ) ) ;
and ( 
    .Z ( edt_scan_in_295 ) ,
    .I0 ( edt_decompressor_out_295 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_295 ) ) ;
and ( 
    .Z ( edt_scan_in_601 ) ,
    .I0 ( edt_decompressor_out_601 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_601 ) ) ;
and ( 
    .Z ( edt_scan_in_598 ) ,
    .I0 ( edt_decompressor_out_598 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_598 ) ) ;
and ( 
    .Z ( edt_scan_in_599 ) ,
    .I0 ( edt_decompressor_out_599 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_599 ) ) ;
and ( 
    .Z ( edt_scan_in_519 ) ,
    .I0 ( edt_decompressor_out_519 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_519 ) ) ;
and ( 
    .Z ( edt_scan_in_596 ) ,
    .I0 ( edt_decompressor_out_596 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_596 ) ) ;
and ( 
    .Z ( edt_scan_in_518 ) ,
    .I0 ( edt_decompressor_out_518 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_518 ) ) ;
and ( 
    .Z ( edt_scan_in_620 ) ,
    .I0 ( edt_decompressor_out_620 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_620 ) ) ;
and ( 
    .Z ( edt_scan_in_311 ) ,
    .I0 ( edt_decompressor_out_311 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_311 ) ) ;
and ( 
    .Z ( edt_scan_in_790 ) ,
    .I0 ( edt_decompressor_out_790 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_790 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.DI_ ) ,
    .IN ( constant_shift_controller_i.N96 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_0 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_0.QT ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_16 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_17 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_18 ) ,
    .A ( GND ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_VL_LSI_MUX21_24108.I0 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_0.QT ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.DI_ ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.ED ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_0.E_ ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.CD_ ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_18 ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_0.ED ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_hold_reg_11_reg_0.U6.I2 ( 
    .I0 ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_16 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.Q1 ) ,
    .S ( constant_shift_controller_i.control_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_17 ) ) ;
DFF constant_shift_controller_i.control_hold_reg_11_reg_0.U6.I3 ( 
    .CK ( constant_shift_controller_i.control_hold_reg_11_reg_0.CPI_ ) ,
    .D ( constant_shift_controller_i.control_hold_reg_11_reg_0.U6.Q1 ) ,
    .Q ( constant_shift_controller_i.control_hold_reg_11_reg_0.QT ) ) ;
and ( 
    .Z ( edt_scan_in_752 ) ,
    .I0 ( edt_decompressor_out_752 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_752 ) ) ;
and ( 
    .Z ( edt_scan_in_621 ) ,
    .I0 ( edt_decompressor_out_621 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_621 ) ) ;
and ( 
    .Z ( edt_scan_in_310 ) ,
    .I0 ( edt_decompressor_out_310 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_310 ) ) ;
and ( 
    .Z ( edt_scan_in_791 ) ,
    .I0 ( edt_decompressor_out_791 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_791 ) ) ;
and ( 
    .Z ( edt_scan_in_309 ) ,
    .I0 ( edt_decompressor_out_309 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_309 ) ) ;
and ( 
    .Z ( edt_scan_in_597 ) ,
    .I0 ( edt_decompressor_out_597 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_597 ) ) ;
and ( 
    .Z ( edt_scan_in_593 ) ,
    .I0 ( edt_decompressor_out_593 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_593 ) ) ;
and ( 
    .Z ( edt_scan_in_595 ) ,
    .I0 ( edt_decompressor_out_595 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_595 ) ) ;
and ( 
    .Z ( edt_scan_in_591 ) ,
    .I0 ( edt_decompressor_out_591 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_591 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.DI_ ) ,
    .IN ( n54 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.CPI_ ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.CDNI_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_3 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.CD ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.CD_ ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_reg_2.CD ) ) ;
and ( 
    .Z ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.D_1 ) ,
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_2.DI_ ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.CD_ ) ) ;
MUX21 constant_shift_controller_i.control_shift_reg_11_reg_2.U5.I2 ( 
    .I0 ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.D_1 ) ,
    .I1 ( constant_shift_controller_i.control_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.Q1 ) ,
    .S ( constant_shift_controller_i.control_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF constant_shift_controller_i.control_shift_reg_11_reg_2.U5.I3 ( 
    .CK ( constant_shift_controller_i.control_shift_reg_11_reg_2.CPI_ ) ,
    .D ( constant_shift_controller_i.control_shift_reg_11_reg_2.U5.Q1 ) ,
    .Q ( constant_shift_controller_i.control_shift_reg_11_2 ) ) ;
and ( 
    .Z ( edt_scan_in_781 ) ,
    .I0 ( edt_decompressor_out_781 ) ,
    .I1 ( constant_shift_controller_i.bias_inputs_781 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n7 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_0_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n311 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n320 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n331 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n340 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n351 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_2_6 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n360 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_10_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n371 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n381 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_4_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n391 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_12_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n401 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_11_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n410 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n421 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_3_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n431 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_8_5 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n461 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_7 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n441 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_6_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n451 ) ,
    .IN ( constant_shift_controller_i.control_hold_reg_7_0 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n471 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_13_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n481 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_2_4 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n491 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_5_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n501 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_1_2 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n511 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_11_5 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I17 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I20 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I18 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I22 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I26 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I28 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I30 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n261 ) ,
    .IN ( constant_shift_controller_i.n160 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n271 ) ,
    .IN ( constant_shift_controller_i.n160 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n280 ) ,
    .IN ( constant_shift_controller_i.n271 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n5 ) ,
    .IN ( constant_shift_controller_i.control_shift_reg_9_3 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2821 ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I22 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.CTS_lsi_ss_clk_delay2761 ) ,
    .IN ( constant_shift_controller_i.net_LSI_EDT_CLOCK_power_clock_gate_G2B2I28 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC16.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n231 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC16.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n240 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC16.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_2 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_2 ) ,
    .I0 ( constant_shift_controller_i.PIC16.AB ) ,
    .I1 ( constant_shift_controller_i.PIC16.CD ) ,
    .I2 ( constant_shift_controller_i.PIC16.EF ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC17.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n200 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC17.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n210 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC17.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_3 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_3 ) ,
    .I0 ( constant_shift_controller_i.PIC17.AB ) ,
    .I1 ( constant_shift_controller_i.PIC17.CD ) ,
    .I2 ( constant_shift_controller_i.PIC17.EF ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC18.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n260 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC18.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n270 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC18.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_1 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_1 ) ,
    .I0 ( constant_shift_controller_i.PIC18.AB ) ,
    .I1 ( constant_shift_controller_i.PIC18.CD ) ,
    .I2 ( constant_shift_controller_i.PIC18.EF ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC19.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n1010 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC19.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n1270 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC19.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_6 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_6 ) ,
    .I0 ( constant_shift_controller_i.PIC19.AB ) ,
    .I1 ( constant_shift_controller_i.PIC19.CD ) ,
    .I2 ( constant_shift_controller_i.PIC19.EF ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC20.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n1400 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC20.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n1510 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC20.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_5 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_5 ) ,
    .I0 ( constant_shift_controller_i.PIC20.AB ) ,
    .I1 ( constant_shift_controller_i.PIC20.CD ) ,
    .I2 ( constant_shift_controller_i.PIC20.EF ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n201 ) ,
    .IN ( edt_shift_const_en ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n160 ) ,
    .IN ( constant_shift_controller_i.n171 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n171 ) ,
    .IN ( constant_shift_controller_i.n232 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n181 ) ,
    .IN ( constant_shift_controller_i.n191 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n191 ) ,
    .IN ( constant_shift_controller_i.n241 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n130 ) ,
    .IN ( constant_shift_controller_i.n140 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n140 ) ,
    .IN ( constant_shift_controller_i.n211 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n211 ) ,
    .IN ( constant_shift_controller_i.n151 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n151 ) ,
    .IN ( constant_shift_controller_i.n2 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n220 ) ,
    .IN ( edt_channels_in_0 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n232 ) ,
    .IN ( constant_shift_controller_i.n181 ) ) ;
not ( 
    .O1 ( constant_shift_controller_i.n241 ) ,
    .IN ( constant_shift_controller_i.n201 ) ) ;
buf ( 
    .O1 ( constant_shift_controller_i.n2 ) ,
    .IN ( constant_shift_controller_i.n220 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC15.AB ) ,
    .I0 ( constant_shift_controller_i.n910 ) ,
    .I1 ( constant_shift_controller_i.n170 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC15.CD ) ,
    .I0 ( constant_shift_controller_i.n1110 ) ,
    .I1 ( constant_shift_controller_i.n180 ) ) ;
or ( 
    .Z ( constant_shift_controller_i.PIC15.EF ) ,
    .I0 ( constant_shift_controller_i.n271 ) ,
    .I1 ( edt_channels_in_4 ) ) ;
and ( 
    .Z ( edt_channels_out_from_constant_shift_control_4 ) ,
    .I0 ( constant_shift_controller_i.PIC15.AB ) ,
    .I1 ( constant_shift_controller_i.PIC15.CD ) ,
    .I2 ( constant_shift_controller_i.PIC15.EF ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_19 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n152 ) ) ;
xor ( 
    .Z ( xor_decoder.n39 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_encoded_masks_76 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_36 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_decoder.n37 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_2 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_3 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_19 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n48 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_8 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n144 ) ) ;
xor ( 
    .Z ( xor_decoder.n190 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_encoded_masks_4 ) ) ;
xor ( 
    .Z ( xor_decoder.n136 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_encoded_masks_138 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_12 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_33 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n38 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_29 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.n36 ) ) ;
xor ( 
    .Z ( xor_decoder.U283.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_encoded_masks_50 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_40 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.U283.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_12 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n135 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_7 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoder.n102 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_encoded_masks_28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_12 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n188 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_24 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n137 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_4 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoder.n33 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_encoded_masks_73 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_34 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.n32 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_41 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n60 ) ) ;
xor ( 
    .Z ( xor_decoder.n137 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_encoded_masks_133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_18 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n102 ) ) ;
xor ( 
    .Z ( xor_decoder.n96 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_encoded_masks_26 ) ) ;
xor ( 
    .Z ( xor_decoder.n188 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_encoded_masks_6 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_50 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n122 ) ) ;
xor ( 
    .Z ( xor_decoder.n127 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_encoded_masks_149 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_11 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n36 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_42 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n58 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_16 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_decoder.n47 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_16 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_decoder.n99 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_11 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n101 ) ) ;
xor ( 
    .Z ( xor_decoder.n115 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_encoded_masks_18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_11 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n193 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_51 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.n121 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_10 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.n130 ) ) ;
xor ( 
    .Z ( xor_decoder.n31 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_encoded_masks_76 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_5 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_21 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n17 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_26 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n37 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_43 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.n56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_23 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n52 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_17 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n52 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_15 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_decoder.n146 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_17 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n104 ) ) ;
xor ( 
    .Z ( xor_decoder.n98 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_encoded_masks_23 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_18 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n115 ) ) ;
xor ( 
    .Z ( xor_decoder.n186 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_encoded_masks_5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_52 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_decoder.n120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_37 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_decoder.n188 ) ) ;
xor ( 
    .Z ( xor_decoder.n122 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_encoded_masks_146 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_6 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoder.n17 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_encoded_masks_84 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_25 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.n32 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_22 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.n42 ) ) ;
xor ( 
    .Z ( xor_decoder.n151 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_encoded_masks_129 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_15 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_decoder.n94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_12 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n96 ) ) ;
xor ( 
    .Z ( xor_decoder.n113 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_encoded_masks_18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_14 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n195 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_46 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_decoder.n124 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_36 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_decoder.n194 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_11 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n127 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_51 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.n134 ) ) ;
xor ( 
    .Z ( xor_decoder.n99 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_encoded_masks_29 ) ) ;
xor ( 
    .Z ( xor_decoder.n104 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_encoded_masks_26 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_19 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n113 ) ) ;
xor ( 
    .Z ( xor_decoder.n195 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_encoded_masks_9 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_2 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_47 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_decoder.n121 ) ) ;
xor ( 
    .Z ( xor_decoder.n124 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_encoded_masks_143 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_52 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_decoder.n133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_14 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n103 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_0 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_1 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_13 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_decoder.n190 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_29 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.n140 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_48 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n122 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_12 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n122 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_9 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_decoder.n131 ) ) ;
xor ( 
    .Z ( xor_decoder.n94 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_encoded_masks_25 ) ) ;
xor ( 
    .Z ( xor_decoder.n101 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_encoded_masks_29 ) ) ;
xor ( 
    .Z ( xor_decoder.U572.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_encoded_masks_11 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_20 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.U572.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_30 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_decoder.n131 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_49 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n123 ) ) ;
xor ( 
    .Z ( xor_decoder.n129 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_encoded_masks_149 ) ) ;
xor ( 
    .Z ( xor_decoder.n119 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_encoded_masks_140 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_13 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_decoder.n98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_10 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.n104 ) ) ;
xor ( 
    .Z ( xor_decoder.n108 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_encoded_masks_14 ) ) ;
xor ( 
    .Z ( xor_decoder.n131 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_encoded_masks_133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_45 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n186 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_13 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_decoder.n124 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_7 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_26 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n102 ) ) ;
xor ( 
    .Z ( xor_decoder.n103 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_encoded_masks_29 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_21 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_26 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n141 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_46 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_decoder.n190 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_8 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n131 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_25 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.n97 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_25 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.n136 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_47 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_decoder.n187 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_44 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n120 ) ) ;
xor ( 
    .Z ( xor_decoder.n93 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_encoded_masks_20 ) ) ;
xor ( 
    .Z ( xor_decoder.n193 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_encoded_masks_9 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_28 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n137 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_15 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_decoder.n55 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_48 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n188 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_45 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_44 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n186 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_5 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_9 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_decoder.n105 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_10 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n196 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_27 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n142 ) ) ;
xor ( 
    .Z ( xor_decoder.n60 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_encoded_masks_59 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_49 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n189 ) ) ;
xor ( 
    .Z ( xor_decoder.n57 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_encoded_masks_56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_43 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n187 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_6 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoder.n85 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_encoded_masks_33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_16 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_decoder.n60 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_4 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_11 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n62 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_42 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n189 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_22 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.n68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_51 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.n82 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_12 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_5 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_17 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n65 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_50 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n188 ) ) ;
xor ( 
    .Z ( xor_decoder.n62 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_encoded_masks_59 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_41 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n191 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_23 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_4 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_52 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_decoder.n81 ) ) ;
xor ( 
    .Z ( xor_decoder.n83 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_encoded_masks_36 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_6 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoder.n63 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_encoded_masks_58 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_51 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_decoder.n187 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_10 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.n65 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_40 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n185 ) ) ;
xor ( 
    .Z ( xor_decoder.n130 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_encoded_masks_146 ) ) ;
xor ( 
    .Z ( xor_decoder.n69 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_encoded_masks_44 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_50 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n135 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_4 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_11 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n88 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_7 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_16 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_decoder.n112 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_18 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n63 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_52 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_decoder.n186 ) ) ;
xor ( 
    .Z ( xor_decoder.n64 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_encoded_masks_59 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_3 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_0 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_21 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_32 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_decoder.n95 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_50 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n83 ) ) ;
xor ( 
    .Z ( xor_decoder.n81 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_encoded_masks_35 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_8 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n92 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_34 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.n162 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_3 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_22 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.n3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_45 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_17 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n117 ) ) ;
xor ( 
    .Z ( xor_decoder.n61 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_encoded_masks_58 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_53 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n185 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_13 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_decoder.n59 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_39 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n192 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_1 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_31 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n101 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_48 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_14 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n90 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_9 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_decoder.n92 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_33 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n168 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_39 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n178 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_23 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n13 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_44 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_33 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n12 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_19 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n61 ) ) ;
xor ( 
    .Z ( xor_decoder.n59 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_encoded_masks_53 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_38 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_decoder.n193 ) ) ;
xor ( 
    .Z ( xor_decoder.U374.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_encoded_masks_41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_20 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.U374.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_30 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_decoder.n92 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_49 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n84 ) ) ;
xor ( 
    .Z ( xor_decoder.n90 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_encoded_masks_39 ) ) ;
xor ( 
    .Z ( xor_decoder.n80 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_encoded_masks_30 ) ) ;
xor ( 
    .Z ( xor_decoder.n4 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_encoded_masks_94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_43 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.n4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_34 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.n6 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_12 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n57 ) ) ;
xor ( 
    .Z ( xor_decoder.n74 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_encoded_masks_48 ) ) ;
xor ( 
    .Z ( xor_decoder.n92 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_encoded_masks_23 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_46 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_decoder.n85 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_13 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_decoder.n85 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_0 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_25 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.n162 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_21 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_42 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n6 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_35 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.n5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_19 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n74 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_2 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_47 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_decoder.n82 ) ) ;
xor ( 
    .Z ( xor_decoder.n91 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_encoded_masks_36 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_38 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_decoder.n166 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_26 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n167 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_1 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_49 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n6 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_36 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_decoder.n11 ) ) ;
xor ( 
    .Z ( xor_decoder.n76 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_encoded_masks_48 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_29 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.n101 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_37 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_decoder.n161 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_27 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n168 ) ) ;
xor ( 
    .Z ( xor_decoder.n153 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_encoded_masks_129 ) ) ;
xor ( 
    .Z ( xor_decoder.U44.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_encoded_masks_91 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_20 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.U44.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_48 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_37 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_decoder.n5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_18 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n76 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_28 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n98 ) ) ;
xor ( 
    .Z ( xor_decoder.n24 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_encoded_masks_88 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_36 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_decoder.n167 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_4 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_28 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n163 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_45 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n172 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_10 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.n156 ) ) ;
xor ( 
    .Z ( xor_decoder.n9 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_encoded_masks_98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_5 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_47 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_decoder.n4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_3 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_38 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_decoder.n10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_27 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n103 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_18 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n24 ) ) ;
xor ( 
    .Z ( xor_decoder.n18 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_encoded_masks_86 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_35 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.n161 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_50 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n44 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_29 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.n166 ) ) ;
xor ( 
    .Z ( xor_decoder.n42 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_encoded_masks_65 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_44 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n172 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_19 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n9 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_6 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_46 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_decoder.n7 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_39 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n152 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_39 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n9 ) ) ;
xor ( 
    .Z ( xor_decoder.n65 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_encoded_masks_56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_16 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_decoder.n21 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_11 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n23 ) ) ;
xor ( 
    .Z ( xor_decoder.n88 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_encoded_masks_39 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_22 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.n29 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_41 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n164 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_51 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.n43 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_2 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_14 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n51 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_47 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_decoder.n173 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_10 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.n52 ) ) ;
xor ( 
    .Z ( xor_decoder.n11 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_encoded_masks_98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_51 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.n147 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_41 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n151 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_3 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_14 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n64 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_0 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_17 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n26 ) ) ;
xor ( 
    .Z ( xor_decoder.n20 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_encoded_masks_83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_10 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.n91 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_23 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n39 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_28 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n59 ) ) ;
xor ( 
    .Z ( xor_decoder.U811.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_encoded_masks_110 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_40 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.U811.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_52 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_decoder.n42 ) ) ;
xor ( 
    .Z ( xor_decoder.n157 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_encoded_masks_113 ) ) ;
xor ( 
    .Z ( xor_decoder.n47 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_encoded_masks_69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_46 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_decoder.n176 ) ) ;
xor ( 
    .Z ( xor_decoder.n49 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_encoded_masks_69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_18 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n11 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_52 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_decoder.n146 ) ) ;
xor ( 
    .Z ( xor_decoder.U745.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_encoded_masks_120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_40 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.U745.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n55 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_encoded_masks_55 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_1 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_12 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_24 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_27 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n64 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_3 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_5 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_30 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_decoder.n157 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_15 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_decoder.n42 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_41 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n177 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_0 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_4 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_43 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.n147 ) ) ;
xor ( 
    .Z ( xor_decoder.U110.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_encoded_masks_81 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_20 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.U110.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n25 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_encoded_masks_89 ) ) ;
xor ( 
    .Z ( xor_decoder.n32 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_encoded_masks_78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_51 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.n95 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_2 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_39 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n165 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_6 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_31 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n166 ) ) ;
xor ( 
    .Z ( xor_decoder.n46 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_encoded_masks_63 ) ) ;
xor ( 
    .Z ( xor_decoder.U877.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_encoded_masks_100 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_40 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.U877.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n52 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_encoded_masks_66 ) ) ;
xor ( 
    .Z ( xor_decoder.n155 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_encoded_masks_129 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_50 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n148 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_42 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n149 ) ) ;
xor ( 
    .Z ( xor_decoder.n22 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_encoded_masks_88 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_13 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_decoder.n20 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_1 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_52 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_decoder.n94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_29 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.n62 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_7 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_32 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_decoder.n160 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_12 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n44 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_43 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.n173 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_9 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_decoder.n53 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_13 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_decoder.n150 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_48 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n148 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_41 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n8 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_45 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n146 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_19 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n22 ) ) ;
xor ( 
    .Z ( xor_decoder.n16 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_encoded_masks_85 ) ) ;
xor ( 
    .Z ( xor_decoder.U176.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_encoded_masks_71 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_20 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.U176.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_30 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_decoder.n53 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_8 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n40 ) ) ;
xor ( 
    .Z ( xor_decoder.n51 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_encoded_masks_69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_42 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n175 ) ) ;
xor ( 
    .Z ( xor_decoder.n41 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_encoded_masks_60 ) ) ;
xor ( 
    .Z ( xor_decoder.n146 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_encoded_masks_125 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_49 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n149 ) ) ;
xor ( 
    .Z ( xor_decoder.U19.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_encoded_masks_90 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_40 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.U19.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_44 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n146 ) ) ;
xor ( 
    .Z ( xor_decoder.n109 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_encoded_masks_16 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_14 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n25 ) ) ;
xor ( 
    .Z ( xor_decoder.n30 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_encoded_masks_74 ) ) ;
xor ( 
    .Z ( xor_decoder.n53 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_encoded_masks_53 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_13 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_decoder.n46 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_7 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_14 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n155 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_46 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_decoder.n150 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_11 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n114 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_21 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_32 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_decoder.n56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_8 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n53 ) ) ;
xor ( 
    .Z ( xor_decoder.n148 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_encoded_masks_126 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_47 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_decoder.n147 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_31 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_41 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n125 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_31 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n62 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_5 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_11 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n153 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_32 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_decoder.n4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_5 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoder.U613.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_encoded_masks_140 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_40 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.U613.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_33 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n129 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_34 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.n58 ) ) ;
xor ( 
    .Z ( xor_decoder.n44 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_encoded_masks_66 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_6 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoder.n150 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_encoded_masks_123 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_6 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_43 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.n108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_43 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.n121 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_34 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.n123 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_45 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_15 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_decoder.n16 ) ) ;
xor ( 
    .Z ( xor_decoder.n35 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_encoded_masks_78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_33 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n64 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_11 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n49 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_12 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n148 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_5 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_7 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_42 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n110 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_0 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_42 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n123 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_28 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n190 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_31 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n127 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_44 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n133 ) ) ;
xor ( 
    .Z ( xor_decoder.n21 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_encoded_masks_89 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_19 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n35 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_6 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_8 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n105 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_41 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n112 ) ) ;
xor ( 
    .Z ( xor_decoder.n196 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_encoded_masks_6 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_38 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_decoder.n127 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_29 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_decoder.n193 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_32 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_decoder.n121 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_43 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.n134 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_48 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n44 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_51 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.n4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_38 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_decoder.n153 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_4 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoder.U547.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_encoded_masks_10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_40 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.U547.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_37 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_decoder.n122 ) ) ;
xor ( 
    .Z ( xor_decoder.n118 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_encoded_masks_143 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_42 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n136 ) ) ;
xor ( 
    .Z ( xor_decoder.n23 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_encoded_masks_89 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_49 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n45 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_52 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_decoder.n3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_37 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_decoder.n148 ) ) ;
xor ( 
    .Z ( xor_decoder.n112 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_encoded_masks_19 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_50 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_47 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_decoder.n108 ) ) ;
xor ( 
    .Z ( xor_decoder.n184 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_encoded_masks_0 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_17 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n182 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_3 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_30 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_decoder.n118 ) ) ;
xor ( 
    .Z ( xor_decoder.n187 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_encoded_masks_4 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_49 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n136 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_10 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.n26 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_9 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_decoder.n1 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_15 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_decoder.n107 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_51 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.n108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_46 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_decoder.n111 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_16 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_decoder.n177 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_39 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n126 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_29 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.n127 ) ) ;
xor ( 
    .Z ( xor_decoder.U969.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_encoded_masks_1 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_20 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.U969.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_48 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n135 ) ) ;
xor ( 
    .Z ( xor_decoder.n107 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_encoded_masks_15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_52 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_decoder.n107 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_45 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n107 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_2 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_47 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_decoder.n134 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_7 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_14 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n116 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_44 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n107 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_27 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n129 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_46 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_decoder.n137 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_8 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n1 ) ) ;
xor ( 
    .Z ( xor_decoder.n116 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_encoded_masks_19 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_19 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n178 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_36 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_decoder.n128 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_28 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n124 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_33 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n181 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_13 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_decoder.n111 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_48 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n109 ) ) ;
xor ( 
    .Z ( xor_decoder.n178 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_encoded_masks_108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_35 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.n122 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_34 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_decoder.n189 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_45 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n81 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_34 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.n175 ) ) ;
xor ( 
    .Z ( xor_decoder.n111 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_encoded_masks_13 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_49 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n110 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_18 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n180 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_5 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_35 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n188 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_25 ) ,
    .I0 ( xor_encoded_masks_5 ) ,
    .I1 ( xor_decoder.n189 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_44 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n81 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_33 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n90 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_31 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n179 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_12 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n109 ) ) ;
xor ( 
    .Z ( xor_decoder.n180 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_encoded_masks_108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_6 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_32 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_decoder.n187 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_47 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_decoder.n69 ) ) ;
xor ( 
    .Z ( xor_decoder.n189 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_encoded_masks_8 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_43 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.n82 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_34 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.n84 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_45 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_32 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_decoder.n173 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_3 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_21 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n173 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_51 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.n69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_33 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n195 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_46 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_decoder.n72 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_27 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n195 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_41 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n138 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_42 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n84 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_35 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.n83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_44 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_37 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_decoder.n174 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_13 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_decoder.n163 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_4 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_39 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n113 ) ) ;
xor ( 
    .Z ( xor_decoder.n72 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_encoded_masks_43 ) ) ;
xor ( 
    .Z ( xor_decoder.n173 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_encoded_masks_104 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_52 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_decoder.n68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_30 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_decoder.n183 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_49 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n71 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_26 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n194 ) ) ;
xor ( 
    .Z ( xor_decoder.U679.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_encoded_masks_130 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_40 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.U679.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_41 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n86 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_36 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_decoder.n89 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_47 ) ,
    .I0 ( xor_encoded_masks_27 ) ,
    .I1 ( xor_decoder.n95 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_38 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_decoder.n179 ) ) ;
xor ( 
    .Z ( xor_decoder.n168 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_encoded_masks_119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_50 ) ,
    .I0 ( xor_encoded_masks_93 ) ,
    .I1 ( xor_decoder.n5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_12 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n70 ) ) ;
xor ( 
    .Z ( xor_decoder.U902.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_encoded_masks_101 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_20 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.U902.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_9 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_decoder.n66 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_31 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n193 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_48 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n70 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_22 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_decoder.n186 ) ) ;
xor ( 
    .Z ( xor_decoder.U415.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_encoded_masks_30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_40 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.U415.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n79 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_encoded_masks_33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_46 ) ,
    .I0 ( xor_encoded_masks_21 ) ,
    .I1 ( xor_decoder.n98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_35 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.n174 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_17 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n13 ) ) ;
xor ( 
    .Z ( xor_decoder.n77 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_encoded_masks_49 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_1 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoder.n54 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_encoded_masks_50 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_2 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_43 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.n69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_21 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n187 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_3 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_30 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_decoder.n79 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_49 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n97 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_36 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_decoder.n180 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_16 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_decoder.n8 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_10 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.n13 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_26 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n11 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_13 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_decoder.n72 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_7 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoder.n183 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_encoded_masks_3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_42 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n71 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_24 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n190 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_39 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n87 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_31 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n88 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_48 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n96 ) ) ;
xor ( 
    .Z ( xor_decoder.n8 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_encoded_masks_99 ) ) ;
xor ( 
    .Z ( xor_decoder.n10 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_encoded_masks_99 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_25 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_decoder.n6 ) ) ;
xor ( 
    .Z ( xor_decoder.n68 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_encoded_masks_45 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_8 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n66 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_45 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_23 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n196 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_38 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_decoder.n88 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_32 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_decoder.n82 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_50 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n96 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_19 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n165 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_37 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_decoder.n18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_15 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_decoder.n3 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_11 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_28 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n7 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_14 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n77 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_44 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_37 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_decoder.n83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_4 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoder.n165 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_encoded_masks_118 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_38 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_decoder.n23 ) ) ;
xor ( 
    .Z ( xor_decoder.n3 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_encoded_masks_95 ) ) ;
xor ( 
    .Z ( xor_decoder.n5 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_encoded_masks_96 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_27 ) ,
    .I0 ( xor_encoded_masks_90 ) ,
    .I1 ( xor_decoder.n12 ) ) ;
xor ( 
    .Z ( xor_decoder.n73 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_encoded_masks_49 ) ) ;
xor ( 
    .Z ( xor_decoder.U836.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_encoded_masks_111 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_20 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.U836.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_51 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.n160 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_14 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n12 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_9 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_decoder.n14 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_2 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_15 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_decoder.n68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_29 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.n88 ) ) ;
xor ( 
    .Z ( xor_decoder.n170 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_encoded_masks_103 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_41 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n47 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_1 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoder.n167 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_encoded_masks_118 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_52 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_decoder.n159 ) ) ;
xor ( 
    .Z ( xor_decoder.n12 ) ,
    .I0 ( xor_encoded_masks_95 ) ,
    .I1 ( xor_encoded_masks_99 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_21 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n134 ) ) ;
xor ( 
    .Z ( xor_decoder.n2 ) ,
    .I0 ( xor_encoded_masks_91 ) ,
    .I1 ( xor_encoded_masks_90 ) ) ;
xor ( 
    .Z ( xor_decoder.n144 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_encoded_masks_123 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_29 ) ,
    .I0 ( xor_encoded_masks_96 ) ,
    .I1 ( xor_decoder.n10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_17 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_41 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n73 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_5 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_2 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_30 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_decoder.n170 ) ) ;
xor ( 
    .Z ( xor_decoder.U217.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_encoded_masks_60 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_40 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.U217.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_21 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n160 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_33 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n51 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_18 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n167 ) ) ;
xor ( 
    .Z ( xor_decoder.U85.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_encoded_masks_80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_40 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.U85.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_13 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_decoder.n7 ) ) ;
xor ( 
    .Z ( xor_decoder.n134 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_encoded_masks_134 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_0 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_decoder.n2 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_30 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_decoder.n144 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_30 ) ,
    .I0 ( xor_encoded_masks_97 ) ,
    .I1 ( xor_decoder.n1 ) ) ;
xor ( 
    .Z ( xor_decoder.n149 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_encoded_masks_128 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_16 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_decoder.n73 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_4 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoder.U349.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_encoded_masks_40 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_40 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.U349.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n38 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_encoded_masks_79 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_6 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_50 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_43 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.n43 ) ) ;
xor ( 
    .Z ( xor_decoder.n160 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_encoded_masks_114 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_34 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.n45 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_16 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_decoder.n164 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_52 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_decoder.n55 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_41 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n21 ) ) ;
xor ( 
    .Z ( xor_decoder.n7 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_encoded_masks_93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_23 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n143 ) ) ;
xor ( 
    .Z ( xor_decoder.n13 ) ,
    .I0 ( xor_encoded_masks_94 ) ,
    .I1 ( xor_encoded_masks_96 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_31 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n153 ) ) ;
xor ( 
    .Z ( xor_decoder.n1 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_encoded_masks_93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_24 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n150 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_50 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n70 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_13 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_decoder.n33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_7 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_4 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_42 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n45 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_23 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n169 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_31 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n49 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_17 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n169 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_51 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.n56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_39 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n22 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_12 ) ,
    .I0 ( xor_encoded_masks_98 ) ,
    .I1 ( xor_decoder.n5 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_22 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.n133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_32 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_decoder.n147 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_23 ) ,
    .I0 ( xor_encoded_masks_128 ) ,
    .I1 ( xor_decoder.n156 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_8 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n27 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_49 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n32 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_45 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n42 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_22 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.n159 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_32 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_decoder.n43 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_15 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_decoder.n159 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_50 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n57 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_3 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_19 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n139 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_33 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n155 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_22 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.n146 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_9 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_decoder.n27 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_48 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_43 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.n95 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_44 ) ,
    .I0 ( xor_encoded_masks_68 ) ,
    .I1 ( xor_decoder.n42 ) ) ;
xor ( 
    .Z ( xor_decoder.n162 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_encoded_masks_118 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_37 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_decoder.n44 ) ) ;
xor ( 
    .Z ( xor_decoder.n164 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_encoded_masks_119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_4 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_9 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_decoder.n157 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_44 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n16 ) ) ;
xor ( 
    .Z ( xor_decoder.n139 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_encoded_masks_138 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_7 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_34 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.n149 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_28 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n150 ) ) ;
xor ( 
    .Z ( xor_decoder.n34 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_encoded_masks_79 ) ) ;
xor ( 
    .Z ( xor_decoder.n15 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_encoded_masks_80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_47 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_decoder.n30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_42 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n97 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_47 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_decoder.n43 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_24 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n163 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_38 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_decoder.n49 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_14 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n168 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_49 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n58 ) ) ;
xor ( 
    .Z ( xor_decoder.n145 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_encoded_masks_120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_45 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n16 ) ) ;
xor ( 
    .Z ( xor_decoder.U704.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_encoded_masks_131 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_20 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.U704.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_8 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n14 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_35 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.n148 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_27 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n155 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_15 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_decoder.n29 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_0 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_46 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_decoder.n33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_46 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_decoder.n46 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_35 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.n44 ) ) ;
xor ( 
    .Z ( xor_decoder.n159 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_encoded_masks_115 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_48 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n57 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_0 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_42 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n19 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_1 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_36 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_decoder.n154 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_26 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n154 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_5 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoder.n29 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_encoded_masks_75 ) ) ;
xor ( 
    .Z ( xor_decoder.n26 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_encoded_masks_86 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_45 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n29 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_36 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_decoder.n50 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_47 ) ,
    .I0 ( xor_encoded_masks_57 ) ,
    .I1 ( xor_decoder.n56 ) ) ;
xor ( 
    .Z ( xor_decoder.n156 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_encoded_masks_126 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_43 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.n17 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_25 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.n149 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_6 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_14 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n38 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_44 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n29 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_46 ) ,
    .I0 ( xor_encoded_masks_51 ) ,
    .I1 ( xor_decoder.n59 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_5 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoder.n6 ) ,
    .I0 ( xor_encoded_masks_92 ) ,
    .I1 ( xor_encoded_masks_98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_31 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n140 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_18 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n37 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_43 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.n30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_45 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n55 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_6 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_18 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n141 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_9_24 ) ,
    .I0 ( xor_encoded_masks_99 ) ,
    .I1 ( xor_decoder.n7 ) ) ;
xor ( 
    .Z ( xor_decoder.n97 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_encoded_masks_28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_32 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_decoder.n134 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_26 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n128 ) ) ;
xor ( 
    .Z ( xor_decoder.n37 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_encoded_masks_78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_42 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n32 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_44 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n55 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_7 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoder.n141 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_encoded_masks_138 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_24 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n98 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_33 ) ,
    .I0 ( xor_encoded_masks_13 ) ,
    .I1 ( xor_decoder.n116 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_25 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.n123 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_15 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_decoder.n120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_17 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n39 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_8 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n157 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_23 ) ,
    .I0 ( xor_encoded_masks_28 ) ,
    .I1 ( xor_decoder.n104 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_34 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.n110 ) ) ;
xor ( 
    .Z ( xor_decoder.n110 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_encoded_masks_18 ) ) ;
xor ( 
    .Z ( xor_decoder.n123 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_encoded_masks_148 ) ) ;
xor ( 
    .Z ( xor_decoder.n125 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_encoded_masks_149 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_16 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_decoder.n34 ) ) ;
xor ( 
    .Z ( xor_decoder.n40 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_encoded_masks_63 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_21 ) ,
    .I0 ( xor_encoded_masks_129 ) ,
    .I1 ( xor_decoder.n147 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_22 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.n94 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_31 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n114 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_24 ) ,
    .I0 ( xor_encoded_masks_19 ) ,
    .I1 ( xor_decoder.n111 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_24 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n124 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_16 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_decoder.n125 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_3 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_30 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_decoder.n40 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_29 ) ,
    .I0 ( xor_encoded_masks_126 ) ,
    .I1 ( xor_decoder.n153 ) ) ;
xor ( 
    .Z ( xor_decoder.n147 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_encoded_masks_124 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_21 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n95 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_32 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_decoder.n108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_26 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n115 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_23 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n130 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_17 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n130 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_51 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.n30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_39 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n48 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_2 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_10 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.n117 ) ) ;
xor ( 
    .Z ( xor_decoder.n95 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_encoded_masks_24 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_37 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_decoder.n109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_25 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.n110 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_37 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_decoder.n135 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_11 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n179 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_22 ) ,
    .I0 ( xor_encoded_masks_146 ) ,
    .I1 ( xor_decoder.n120 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_15 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_decoder.n186 ) ) ;
xor ( 
    .Z ( xor_decoder.n128 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_encoded_masks_148 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_52 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_decoder.n29 ) ) ;
xor ( 
    .Z ( xor_decoder.n114 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_encoded_masks_19 ) ) ;
xor ( 
    .Z ( xor_decoder.U506.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_encoded_masks_21 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_20 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.U506.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_38 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_decoder.n114 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_28 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n111 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_38 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_decoder.n140 ) ) ;
xor ( 
    .Z ( xor_decoder.n174 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_encoded_masks_106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_21 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n121 ) ) ;
xor ( 
    .Z ( xor_decoder.n191 ) ,
    .I0 ( xor_encoded_masks_6 ) ,
    .I1 ( xor_encoded_masks_9 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_18 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n128 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_0 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_1 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_35 ) ,
    .I0 ( xor_encoded_masks_15 ) ,
    .I1 ( xor_decoder.n109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_27 ) ,
    .I0 ( xor_encoded_masks_10 ) ,
    .I1 ( xor_decoder.n116 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_39 ) ,
    .I0 ( xor_encoded_masks_139 ) ,
    .I1 ( xor_decoder.n139 ) ) ;
xor ( 
    .Z ( xor_decoder.n121 ) ,
    .I0 ( xor_encoded_masks_142 ) ,
    .I1 ( xor_encoded_masks_144 ) ) ;
xor ( 
    .Z ( xor_decoder.n126 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_encoded_masks_148 ) ) ;
xor ( 
    .Z ( xor_decoder.n117 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_encoded_masks_16 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_19 ) ,
    .I0 ( xor_encoded_masks_20 ) ,
    .I1 ( xor_decoder.n100 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_36 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_decoder.n115 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_2 ) ,
    .I0 ( xor_encoded_masks_14 ) ,
    .I1 ( xor_decoder.n106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_3 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_6 ) ,
    .I0 ( xor_encoded_masks_8 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoder.U638.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_144 ) ,
    .I1 ( xor_encoded_masks_141 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_20 ) ,
    .I0 ( xor_encoded_masks_145 ) ,
    .I1 ( xor_decoder.U638.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_19 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n126 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_33 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n103 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_9 ) ,
    .I0 ( xor_encoded_masks_141 ) ,
    .I1 ( xor_decoder.n118 ) ) ;
xor ( 
    .Z ( xor_decoder.n100 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_encoded_masks_28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_29 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.n114 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_33 ) ,
    .I0 ( xor_encoded_masks_133 ) ,
    .I1 ( xor_decoder.n142 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_13 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_decoder.n176 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_5 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_1 ) ,
    .I0 ( xor_encoded_masks_143 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_34 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.n97 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_26 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n180 ) ) ;
xor ( 
    .Z ( xor_decoder.n106 ) ,
    .I0 ( xor_encoded_masks_11 ) ,
    .I1 ( xor_encoded_masks_10 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_34 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_decoder.n136 ) ) ;
xor ( 
    .Z ( xor_decoder.n181 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_encoded_masks_109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_8 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n183 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_25 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.n175 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_7 ) ,
    .I0 ( xor_encoded_masks_149 ) ,
    .I1 ( xor_decoder.n119 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_35 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.n135 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_12 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n174 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_21 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n56 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_7 ) ,
    .I0 ( xor_encoded_masks_9 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_18 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n194 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_26 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n89 ) ) ;
xor ( 
    .Z ( xor_decoder.n175 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_encoded_masks_108 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_8 ) ,
    .I0 ( xor_encoded_masks_140 ) ,
    .I1 ( xor_decoder.n118 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_36 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_decoder.n141 ) ) ;
xor ( 
    .Z ( xor_decoder.n176 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_encoded_masks_103 ) ) ;
xor ( 
    .Z ( xor_decoder.n56 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_encoded_masks_54 ) ) ;
xor ( 
    .Z ( xor_decoder.n171 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_encoded_masks_100 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_37 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_decoder.n70 ) ) ;
xor ( 
    .Z ( xor_decoder.n192 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_encoded_masks_8 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_25 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.n84 ) ) ;
xor ( 
    .Z ( xor_decoder.n89 ) ,
    .I0 ( xor_encoded_masks_37 ) ,
    .I1 ( xor_encoded_masks_38 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_24 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n176 ) ) ;
xor ( 
    .Z ( xor_decoder.n105 ) ,
    .I0 ( xor_encoded_masks_12 ) ,
    .I1 ( xor_encoded_masks_13 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_15 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_decoder.n172 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_23 ) ,
    .I0 ( xor_encoded_masks_58 ) ,
    .I1 ( xor_decoder.n65 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_9 ) ,
    .I0 ( xor_encoded_masks_1 ) ,
    .I1 ( xor_decoder.n183 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_38 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_decoder.n75 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_19 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_decoder.n192 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_30 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_decoder.n66 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_28 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n85 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_18 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n89 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_2 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoder.n158 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_encoded_masks_110 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_30 ) ,
    .I0 ( xor_encoded_masks_17 ) ,
    .I1 ( xor_decoder.n105 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_7 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoder.n177 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_encoded_masks_109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_22 ) ,
    .I0 ( xor_encoded_masks_56 ) ,
    .I1 ( xor_decoder.n55 ) ) ;
xor ( 
    .Z ( xor_decoder.n182 ) ,
    .I0 ( xor_encoded_masks_104 ) ,
    .I1 ( xor_encoded_masks_106 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_39 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n74 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_1 ) ,
    .I0 ( xor_encoded_masks_3 ) ,
    .I1 ( xor_decoder.n184 ) ) ;
xor ( 
    .Z ( xor_decoder.n66 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_encoded_masks_43 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_27 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n90 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_16 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_decoder.n86 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_29 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.n179 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_9 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_decoder.n170 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_8 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n79 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_14 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n181 ) ) ;
xor ( 
    .Z ( xor_decoder.n58 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_encoded_masks_58 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_0 ) ,
    .I0 ( xor_encoded_masks_102 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_3 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_16 ) ,
    .I0 ( xor_encoded_masks_2 ) ,
    .I1 ( xor_decoder.n191 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_14_14 ) ,
    .I0 ( xor_encoded_masks_148 ) ,
    .I1 ( xor_decoder.n129 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_2 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_23 ) ,
    .I0 ( xor_encoded_masks_38 ) ,
    .I1 ( xor_decoder.n91 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_17 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n91 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_28 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n176 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_23 ) ,
    .I0 ( xor_encoded_masks_18 ) ,
    .I1 ( xor_decoder.n117 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_9 ) ,
    .I0 ( xor_encoded_masks_31 ) ,
    .I1 ( xor_decoder.n79 ) ) ;
xor ( 
    .Z ( xor_decoder.n172 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_encoded_masks_105 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_24 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n59 ) ) ;
xor ( 
    .Z ( xor_decoder.n179 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_encoded_masks_109 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_33 ) ,
    .I0 ( xor_encoded_masks_43 ) ,
    .I1 ( xor_decoder.n77 ) ) ;
xor ( 
    .Z ( xor_decoder.n185 ) ,
    .I0 ( xor_encoded_masks_0 ) ,
    .I1 ( xor_encoded_masks_6 ) ) ;
xor ( 
    .Z ( xor_decoder.n120 ) ,
    .I0 ( xor_encoded_masks_147 ) ,
    .I1 ( xor_encoded_masks_145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_29 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.n75 ) ) ;
xor ( 
    .Z ( xor_decoder.U481.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_encoded_masks_20 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_40 ) ,
    .I0 ( xor_encoded_masks_26 ) ,
    .I1 ( xor_decoder.U481.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_22 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_decoder.n81 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_1 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_decoder.n80 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_27 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n181 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_42 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n162 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_48 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n174 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_52 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_decoder.n16 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_1_22 ) ,
    .I0 ( xor_encoded_masks_16 ) ,
    .I1 ( xor_decoder.n107 ) ) ;
xor ( 
    .Z ( xor_decoder.n67 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_encoded_masks_40 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_26 ) ,
    .I0 ( xor_encoded_masks_50 ) ,
    .I1 ( xor_decoder.n63 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_10 ) ,
    .I0 ( xor_encoded_masks_105 ) ,
    .I1 ( xor_decoder.n182 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_34 ) ,
    .I0 ( xor_encoded_masks_46 ) ,
    .I1 ( xor_decoder.n71 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_0_17 ) ,
    .I0 ( xor_encoded_masks_4 ) ,
    .I1 ( xor_decoder.n185 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_28 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n72 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_41 ) ,
    .I0 ( xor_encoded_masks_23 ) ,
    .I1 ( xor_decoder.n99 ) ) ;
xor ( 
    .Z ( xor_decoder.n84 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_encoded_masks_38 ) ) ;
xor ( 
    .Z ( xor_decoder.U440.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_34 ) ,
    .I1 ( xor_encoded_masks_31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_20 ) ,
    .I0 ( xor_encoded_masks_35 ) ,
    .I1 ( xor_decoder.U440.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_43 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.n160 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_49 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n175 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_51 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.n17 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_0 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_decoder.n67 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_25 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.n58 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_35 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.n70 ) ) ;
xor ( 
    .Z ( xor_decoder.n194 ) ,
    .I0 ( xor_encoded_masks_7 ) ,
    .I1 ( xor_encoded_masks_8 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_27 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n77 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_39 ) ,
    .I0 ( xor_encoded_masks_29 ) ,
    .I1 ( xor_decoder.n100 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_24 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n85 ) ) ;
xor ( 
    .Z ( xor_decoder.n87 ) ,
    .I0 ( xor_encoded_masks_33 ) ,
    .I1 ( xor_encoded_masks_38 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_2 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_6 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoder.n78 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_encoded_masks_46 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_36 ) ,
    .I0 ( xor_encoded_masks_44 ) ,
    .I1 ( xor_decoder.n76 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_26 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n76 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_3 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.n93 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_19 ) ,
    .I0 ( xor_encoded_masks_30 ) ,
    .I1 ( xor_decoder.n87 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_29 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.n23 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_5 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_10 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.n78 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_25 ) ,
    .I0 ( xor_encoded_masks_45 ) ,
    .I1 ( xor_decoder.n71 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_37 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_decoder.n96 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_46 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_decoder.n163 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_49 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n19 ) ) ;
xor ( 
    .Z ( xor_decoder.n75 ) ,
    .I0 ( xor_encoded_masks_47 ) ,
    .I1 ( xor_encoded_masks_49 ) ) ;
xor ( 
    .Z ( xor_decoder.n71 ) ,
    .I0 ( xor_encoded_masks_42 ) ,
    .I1 ( xor_encoded_masks_48 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_38 ) ,
    .I0 ( xor_encoded_masks_22 ) ,
    .I1 ( xor_decoder.n101 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_21 ) ,
    .I0 ( xor_encoded_masks_39 ) ,
    .I1 ( xor_decoder.n82 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_23 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n182 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_47 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_decoder.n160 ) ) ;
xor ( 
    .Z ( xor_decoder.n163 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_encoded_masks_113 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_15 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_decoder.n133 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_48 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_11 ) ,
    .I0 ( xor_encoded_masks_40 ) ,
    .I1 ( xor_decoder.n75 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_31 ) ,
    .I0 ( xor_encoded_masks_48 ) ,
    .I1 ( xor_decoder.n75 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_24 ) ,
    .I0 ( xor_encoded_masks_49 ) ,
    .I1 ( xor_decoder.n72 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_35 ) ,
    .I0 ( xor_encoded_masks_25 ) ,
    .I1 ( xor_decoder.n96 ) ) ;
xor ( 
    .Z ( xor_decoder.n19 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_encoded_masks_88 ) ) ;
xor ( 
    .Z ( xor_decoder.n82 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_encoded_masks_34 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_22 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.n172 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_44 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n159 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_26 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n50 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_12 ) ,
    .I0 ( xor_encoded_masks_118 ) ,
    .I1 ( xor_decoder.n161 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_5 ) ,
    .I0 ( xor_encoded_masks_107 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_32 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_decoder.n17 ) ) ;
xor ( 
    .Z ( xor_decoder.n138 ) ,
    .I0 ( xor_encoded_masks_136 ) ,
    .I1 ( xor_encoded_masks_139 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_50 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n18 ) ) ;
xor ( 
    .Z ( xor_decoder.n135 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_encoded_masks_136 ) ) ;
xor ( 
    .Z ( xor_decoder.n154 ) ,
    .I0 ( xor_encoded_masks_127 ) ,
    .I1 ( xor_encoded_masks_128 ) ) ;
xor ( 
    .Z ( xor_decoder.n70 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_encoded_masks_46 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_4_32 ) ,
    .I0 ( xor_encoded_masks_41 ) ,
    .I1 ( xor_decoder.n69 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_9 ) ,
    .I0 ( xor_encoded_masks_61 ) ,
    .I1 ( xor_decoder.n40 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_2_36 ) ,
    .I0 ( xor_encoded_masks_24 ) ,
    .I1 ( xor_decoder.n102 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_24 ) ,
    .I0 ( xor_encoded_masks_89 ) ,
    .I1 ( xor_decoder.n20 ) ) ;
xor ( 
    .Z ( xor_decoder.U151.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_encoded_masks_70 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_40 ) ,
    .I0 ( xor_encoded_masks_76 ) ,
    .I1 ( xor_decoder.U151.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_45 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n159 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_25 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.n45 ) ) ;
xor ( 
    .Z ( xor_decoder.n161 ) ,
    .I0 ( xor_encoded_masks_111 ) ,
    .I1 ( xor_encoded_masks_116 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_1 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_6 ) ,
    .I0 ( xor_encoded_masks_108 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_31 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n23 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_16 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_decoder.n138 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_4 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.n15 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_11 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n140 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_18 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n154 ) ) ;
xor ( 
    .Z ( xor_decoder.n28 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_encoded_masks_70 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_23 ) ,
    .I0 ( xor_encoded_masks_88 ) ,
    .I1 ( xor_decoder.n26 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_41 ) ,
    .I0 ( xor_encoded_masks_73 ) ,
    .I1 ( xor_decoder.n34 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_3_15 ) ,
    .I0 ( xor_encoded_masks_32 ) ,
    .I1 ( xor_decoder.n81 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_30 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_decoder.n27 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_4 ) ,
    .I0 ( xor_encoded_masks_116 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoder.n45 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_encoded_masks_68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_11 ) ,
    .I0 ( xor_encoded_masks_110 ) ,
    .I1 ( xor_decoder.n166 ) ) ;
xor ( 
    .Z ( xor_decoder.U242.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_encoded_masks_61 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_20 ) ,
    .I0 ( xor_encoded_masks_65 ) ,
    .I1 ( xor_decoder.U242.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_7 ) ,
    .I0 ( xor_encoded_masks_109 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_30 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_decoder.n14 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_17 ) ,
    .I0 ( xor_encoded_masks_130 ) ,
    .I1 ( xor_decoder.n143 ) ) ;
xor ( 
    .Z ( xor_decoder.n140 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_encoded_masks_139 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_16 ) ,
    .I0 ( xor_encoded_masks_122 ) ,
    .I1 ( xor_decoder.n151 ) ) ;
xor ( 
    .Z ( xor_decoder.U308.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_encoded_masks_51 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_20 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.U308.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_22 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.n16 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_39 ) ,
    .I0 ( xor_encoded_masks_79 ) ,
    .I1 ( xor_decoder.n35 ) ) ;
xor ( 
    .Z ( xor_decoder.n86 ) ,
    .I0 ( xor_encoded_masks_36 ) ,
    .I1 ( xor_encoded_masks_39 ) ) ;
xor ( 
    .Z ( xor_decoder.n27 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_encoded_masks_73 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_35 ) ,
    .I0 ( xor_encoded_masks_55 ) ,
    .I1 ( xor_decoder.n57 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_50 ) ,
    .I0 ( xor_encoded_masks_113 ) ,
    .I1 ( xor_decoder.n161 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_24 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n46 ) ) ;
xor ( 
    .Z ( xor_decoder.n166 ) ,
    .I0 ( xor_encoded_masks_117 ) ,
    .I1 ( xor_encoded_masks_119 ) ) ;
xor ( 
    .Z ( xor_decoder.n43 ) ,
    .I0 ( xor_encoded_masks_62 ) ,
    .I1 ( xor_encoded_masks_64 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_8 ) ,
    .I0 ( xor_encoded_masks_100 ) ,
    .I1 ( xor_decoder.n170 ) ) ;
xor ( 
    .Z ( xor_decoder.n14 ) ,
    .I0 ( xor_encoded_masks_82 ) ,
    .I1 ( xor_encoded_masks_83 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_13 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_decoder.n137 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_10 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_decoder.n143 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_17 ) ,
    .I0 ( xor_encoded_masks_120 ) ,
    .I1 ( xor_decoder.n156 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_1 ) ,
    .I0 ( xor_encoded_masks_53 ) ,
    .I1 ( xor_decoder.n54 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_28 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n20 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_3 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_32 ) ,
    .I0 ( xor_encoded_masks_71 ) ,
    .I1 ( xor_decoder.n30 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_36 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_decoder.n63 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_48 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n161 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_2 ) ,
    .I0 ( xor_encoded_masks_64 ) ,
    .I1 ( xor_decoder.n41 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_10 ) ,
    .I0 ( xor_encoded_masks_115 ) ,
    .I1 ( xor_decoder.n169 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_21 ) ,
    .I0 ( xor_encoded_masks_69 ) ,
    .I1 ( xor_decoder.n43 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_4 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.n171 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_36 ) ,
    .I0 ( xor_encoded_masks_84 ) ,
    .I1 ( xor_decoder.n24 ) ) ;
xor ( 
    .Z ( xor_decoder.n142 ) ,
    .I0 ( xor_encoded_masks_135 ) ,
    .I1 ( xor_encoded_masks_139 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_47 ) ,
    .I0 ( xor_encoded_masks_87 ) ,
    .I1 ( xor_decoder.n17 ) ) ;
xor ( 
    .Z ( xor_decoder.n143 ) ,
    .I0 ( xor_encoded_masks_134 ) ,
    .I1 ( xor_encoded_masks_136 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_1 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_decoder.n145 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_10 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.n39 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_27 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n25 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_37 ) ,
    .I0 ( xor_encoded_masks_74 ) ,
    .I1 ( xor_decoder.n31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_31 ) ,
    .I0 ( xor_encoded_masks_78 ) ,
    .I1 ( xor_decoder.n36 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_37 ) ,
    .I0 ( xor_encoded_masks_54 ) ,
    .I1 ( xor_decoder.n57 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_49 ) ,
    .I0 ( xor_encoded_masks_119 ) ,
    .I1 ( xor_decoder.n162 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_29 ) ,
    .I0 ( xor_encoded_masks_66 ) ,
    .I1 ( xor_decoder.n49 ) ) ;
xor ( 
    .Z ( xor_decoder.n169 ) ,
    .I0 ( xor_encoded_masks_114 ) ,
    .I1 ( xor_encoded_masks_116 ) ) ;
xor ( 
    .Z ( xor_decoder.n50 ) ,
    .I0 ( xor_encoded_masks_67 ) ,
    .I1 ( xor_encoded_masks_68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_50 ) ,
    .I0 ( xor_encoded_masks_103 ) ,
    .I1 ( xor_decoder.n174 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_35 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.n18 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_14 ) ,
    .I0 ( xor_encoded_masks_138 ) ,
    .I1 ( xor_decoder.n142 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_46 ) ,
    .I0 ( xor_encoded_masks_81 ) ,
    .I1 ( xor_decoder.n20 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_13_0 ) ,
    .I0 ( xor_encoded_masks_132 ) ,
    .I1 ( xor_decoder.n132 ) ) ;
xor ( 
    .Z ( xor_decoder.U770.SYNTEST_VL_xor_28002_299 ) ,
    .I0 ( xor_encoded_masks_124 ) ,
    .I1 ( xor_encoded_masks_121 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_20 ) ,
    .I0 ( xor_encoded_masks_125 ) ,
    .I1 ( xor_decoder.U770.SYNTEST_VL_xor_28002_299 ) ) ;
xor ( 
    .Z ( xor_decoder.n36 ) ,
    .I0 ( xor_encoded_masks_77 ) ,
    .I1 ( xor_encoded_masks_79 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_26 ) ,
    .I0 ( xor_encoded_masks_80 ) ,
    .I1 ( xor_decoder.n24 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_38 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_decoder.n36 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_28 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n33 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_38 ) ,
    .I0 ( xor_encoded_masks_52 ) ,
    .I1 ( xor_decoder.n62 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_28 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n46 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_11_0 ) ,
    .I0 ( xor_encoded_masks_112 ) ,
    .I1 ( xor_decoder.n158 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_18 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_decoder.n50 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_51 ) ,
    .I0 ( xor_encoded_masks_106 ) ,
    .I1 ( xor_decoder.n173 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_34 ) ,
    .I0 ( xor_encoded_masks_86 ) ,
    .I1 ( xor_decoder.n19 ) ) ;
xor ( 
    .Z ( xor_decoder.n133 ) ,
    .I0 ( xor_encoded_masks_137 ) ,
    .I1 ( xor_encoded_masks_135 ) ) ;
xor ( 
    .Z ( xor_decoder.n132 ) ,
    .I0 ( xor_encoded_masks_131 ) ,
    .I1 ( xor_encoded_masks_130 ) ) ;
xor ( 
    .Z ( xor_decoder.n152 ) ,
    .I0 ( xor_encoded_masks_123 ) ,
    .I1 ( xor_encoded_masks_128 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_0 ) ,
    .I0 ( xor_encoded_masks_72 ) ,
    .I1 ( xor_decoder.n28 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_25 ) ,
    .I0 ( xor_encoded_masks_85 ) ,
    .I1 ( xor_decoder.n19 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_35 ) ,
    .I0 ( xor_encoded_masks_75 ) ,
    .I1 ( xor_decoder.n31 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_7_27 ) ,
    .I0 ( xor_encoded_masks_70 ) ,
    .I1 ( xor_decoder.n38 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_5_39 ) ,
    .I0 ( xor_encoded_masks_59 ) ,
    .I1 ( xor_decoder.n61 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_6_27 ) ,
    .I0 ( xor_encoded_masks_60 ) ,
    .I1 ( xor_decoder.n51 ) ) ;
xor ( 
    .Z ( xor_decoder.n48 ) ,
    .I0 ( xor_encoded_masks_63 ) ,
    .I1 ( xor_encoded_masks_68 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_10_52 ) ,
    .I0 ( xor_encoded_masks_101 ) ,
    .I1 ( xor_decoder.n172 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_8_33 ) ,
    .I0 ( xor_encoded_masks_83 ) ,
    .I1 ( xor_decoder.n25 ) ) ;
xor ( 
    .Z ( xor_decoded_masks_12_9 ) ,
    .I0 ( xor_encoded_masks_121 ) ,
    .I1 ( xor_decoder.n144 ) ) ;
or ( 
    .Z ( config0_decoder9.U52.AB ) ,
    .I0 ( config0_decoder9.n40 ) ,
    .I1 ( masks_hold_reg_7_4 ) ) ;
and ( 
    .Z ( config0_decoder9.U52.ZN ) ,
    .I0 ( config0_decoder9.U52.AB ) ,
    .I1 ( config0_decoder9.n52 ) ) ;
not ( 
    .O1 ( config0_decoder9.n1 ) ,
    .IN ( config0_decoder9.U52.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U76.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n56 ) ) ;
and ( 
    .Z ( config0_decoder9.U76.ZN ) ,
    .I0 ( config0_decoder9.U76.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_4 ) ,
    .IN ( config0_decoder9.U76.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n50 ) ,
    .I0 ( config0_decoder9.n40 ) ,
    .I1 ( masks_hold_reg_7_4 ) ) ;
or ( 
    .Z ( config0_decoder9.U17.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n53 ) ) ;
and ( 
    .Z ( config0_decoder9.U17.ZN ) ,
    .I0 ( config0_decoder9.U17.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_0 ) ,
    .IN ( config0_decoder9.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U37.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n47 ) ) ;
and ( 
    .Z ( config0_decoder9.U37.ZN ) ,
    .I0 ( config0_decoder9.U37.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_12 ) ,
    .IN ( config0_decoder9.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U87.AB ) ,
    .I0 ( config0_decoder9.n57 ) ,
    .I1 ( config0_decoder9.n54 ) ) ;
and ( 
    .Z ( config0_decoder9.U87.ZN ) ,
    .I0 ( config0_decoder9.U87.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_50 ) ,
    .IN ( config0_decoder9.U87.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n49 ) ,
    .I0 ( config0_decoder9.n46 ) ,
    .I1 ( masks_hold_reg_7_1 ) ) ;
or ( 
    .Z ( config0_decoder9.U47.AB ) ,
    .I0 ( config0_decoder9.n56 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U47.ZN ) ,
    .I0 ( config0_decoder9.U47.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_35 ) ,
    .IN ( config0_decoder9.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U77.AB ) ,
    .I0 ( config0_decoder9.n50 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U77.ZN ) ,
    .I0 ( config0_decoder9.U77.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_45 ) ,
    .IN ( config0_decoder9.U77.ZN ) ) ;
nor ( 
    .Z ( config0_decoder9.n37 ) ,
    .I0 ( config0_decoder9.n36 ) ,
    .I1 ( masks_hold_reg_7_6 ) ) ;
nand ( 
    .Z ( config0_decoder9.n58 ) ,
    .I0 ( config0_decoder9.n40 ) ,
    .I1 ( config0_decoder9.n39 ) ) ;
or ( 
    .Z ( config0_decoder9.U34.AB ) ,
    .I0 ( config0_decoder9.n54 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U34.ZN ) ,
    .I0 ( config0_decoder9.U34.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_34 ) ,
    .IN ( config0_decoder9.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U3.AB ) ,
    .I0 ( config0_decoder9.n50 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U3.ZN ) ,
    .I0 ( config0_decoder9.U3.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_30 ) ,
    .IN ( config0_decoder9.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U86.AB ) ,
    .I0 ( config0_decoder9.n57 ) ,
    .I1 ( config0_decoder9.n56 ) ) ;
and ( 
    .Z ( config0_decoder9.U86.ZN ) ,
    .I0 ( config0_decoder9.U86.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_52 ) ,
    .IN ( config0_decoder9.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n44 ) ,
    .I0 ( config0_decoder9.n37 ) ,
    .I1 ( masks_hold_reg_7_1 ) ) ;
or ( 
    .Z ( config0_decoder9.U46.AB ) ,
    .I0 ( config0_decoder9.n54 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U46.ZN ) ,
    .I0 ( config0_decoder9.U46.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_17 ) ,
    .IN ( config0_decoder9.U46.ZN ) ) ;
not ( 
    .O1 ( config0_decoder9.n36 ) ,
    .IN ( masks_hold_reg_7_5 ) ) ;
not ( 
    .O1 ( config0_decoder9.n41 ) ,
    .IN ( masks_hold_reg_7_2 ) ) ;
nor ( 
    .Z ( config0_decoder9.n52 ) ,
    .I0 ( config0_decoder9.n45 ) ,
    .I1 ( config0_decoder9.n36 ) ) ;
or ( 
    .Z ( config0_decoder9.U38.AB ) ,
    .I0 ( config0_decoder9.n54 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U38.ZN ) ,
    .I0 ( config0_decoder9.U38.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_18 ) ,
    .IN ( config0_decoder9.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U35.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U35.ZN ) ,
    .I0 ( config0_decoder9.U35.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_26 ) ,
    .IN ( config0_decoder9.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U2.AB ) ,
    .I0 ( config0_decoder9.n53 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U2.ZN ) ,
    .I0 ( config0_decoder9.U2.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_31 ) ,
    .IN ( config0_decoder9.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U81.AB ) ,
    .I0 ( config0_decoder9.n60 ) ,
    .I1 ( config0_decoder9.n59 ) ) ;
and ( 
    .Z ( config0_decoder9.U81.ZN ) ,
    .I0 ( config0_decoder9.U81.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_8 ) ,
    .IN ( config0_decoder9.U81.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n63 ) ,
    .I0 ( masks_hold_reg_7_2 ) ,
    .I1 ( config0_decoder9.n42 ) ) ;
or ( 
    .Z ( config0_decoder9.U49.AB ) ,
    .I0 ( config0_decoder9.n60 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U49.ZN ) ,
    .I0 ( config0_decoder9.U49.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_39 ) ,
    .IN ( config0_decoder9.U49.ZN ) ) ;
not ( 
    .O1 ( config0_decoder9.n45 ) ,
    .IN ( masks_hold_reg_7_6 ) ) ;
nor ( 
    .Z ( config0_decoder9.n42 ) ,
    .I0 ( config0_decoder9.n39 ) ,
    .I1 ( masks_hold_reg_7_3 ) ) ;
nand ( 
    .Z ( config0_decoder9.n55 ) ,
    .I0 ( config0_decoder9.n52 ) ,
    .I1 ( config0_decoder9.n51 ) ) ;
or ( 
    .Z ( config0_decoder9.U39.AB ) ,
    .I0 ( config0_decoder9.n50 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U39.ZN ) ,
    .I0 ( config0_decoder9.U39.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_29 ) ,
    .IN ( config0_decoder9.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U32.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n59 ) ) ;
and ( 
    .Z ( config0_decoder9.U32.ZN ) ,
    .I0 ( config0_decoder9.U32.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_10 ) ,
    .IN ( config0_decoder9.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U29.AB ) ,
    .I0 ( config0_decoder9.n60 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U29.ZN ) ,
    .I0 ( config0_decoder9.U29.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_24 ) ,
    .IN ( config0_decoder9.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U80.AB ) ,
    .I0 ( config0_decoder9.n60 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U80.ZN ) ,
    .I0 ( config0_decoder9.U80.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_40 ) ,
    .IN ( config0_decoder9.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U48.AB ) ,
    .I0 ( config0_decoder9.n47 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U48.ZN ) ,
    .I0 ( config0_decoder9.U48.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_27 ) ,
    .IN ( config0_decoder9.U48.ZN ) ) ;
nor ( 
    .Z ( config0_decoder9.n35 ) ,
    .I0 ( masks_hold_reg_7_5 ) ,
    .I1 ( masks_hold_reg_7_6 ) ) ;
or ( 
    .Z ( config0_decoder9.U13.AB ) ,
    .I0 ( config0_decoder9.n60 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U13.ZN ) ,
    .I0 ( config0_decoder9.U13.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_23 ) ,
    .IN ( config0_decoder9.U13.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U33.AB ) ,
    .I0 ( config0_decoder9.n53 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U33.ZN ) ,
    .I0 ( config0_decoder9.U33.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_16 ) ,
    .IN ( config0_decoder9.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U28.AB ) ,
    .I0 ( config0_decoder9.n53 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U28.ZN ) ,
    .I0 ( config0_decoder9.U28.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_32 ) ,
    .IN ( config0_decoder9.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U83.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U83.ZN ) ,
    .I0 ( config0_decoder9.U83.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_41 ) ,
    .IN ( config0_decoder9.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U50.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n62 ) ) ;
and ( 
    .Z ( config0_decoder9.U50.ZN ) ,
    .I0 ( config0_decoder9.U50.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_9 ) ,
    .IN ( config0_decoder9.U50.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U30.AB ) ,
    .I0 ( config0_decoder9.n56 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U30.ZN ) ,
    .I0 ( config0_decoder9.U30.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_36 ) ,
    .IN ( config0_decoder9.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U22.AB ) ,
    .I0 ( config0_decoder9.n56 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U22.ZN ) ,
    .I0 ( config0_decoder9.U22.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_20 ) ,
    .IN ( config0_decoder9.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U82.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U82.ZN ) ,
    .I0 ( config0_decoder9.U82.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_42 ) ,
    .IN ( config0_decoder9.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U51.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n50 ) ) ;
and ( 
    .Z ( config0_decoder9.U51.ZN ) ,
    .I0 ( config0_decoder9.U51.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_13 ) ,
    .IN ( config0_decoder9.U51.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U41.AB ) ,
    .I0 ( config0_decoder9.n63 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U41.ZN ) ,
    .I0 ( config0_decoder9.U41.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_25 ) ,
    .IN ( config0_decoder9.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U78.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n54 ) ) ;
and ( 
    .Z ( config0_decoder9.U78.ZN ) ,
    .I0 ( config0_decoder9.U78.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_1 ) ,
    .IN ( config0_decoder9.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U31.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n50 ) ) ;
and ( 
    .Z ( config0_decoder9.U31.ZN ) ,
    .I0 ( config0_decoder9.U31.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_14 ) ,
    .IN ( config0_decoder9.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U21.AB ) ,
    .I0 ( config0_decoder9.n55 ) ,
    .I1 ( config0_decoder9.n54 ) ) ;
and ( 
    .Z ( config0_decoder9.U21.ZN ) ,
    .I0 ( config0_decoder9.U21.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_49 ) ,
    .IN ( config0_decoder9.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n48 ) ,
    .I0 ( config0_decoder9.n46 ) ,
    .I1 ( config0_decoder9.n51 ) ) ;
or ( 
    .Z ( config0_decoder9.U40.AB ) ,
    .I0 ( config0_decoder9.n54 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U40.ZN ) ,
    .I0 ( config0_decoder9.U40.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_33 ) ,
    .IN ( config0_decoder9.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U79.AB ) ,
    .I0 ( config0_decoder9.n55 ) ,
    .I1 ( config0_decoder9.n53 ) ) ;
and ( 
    .Z ( config0_decoder9.U79.ZN ) ,
    .I0 ( config0_decoder9.U79.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_47 ) ,
    .IN ( config0_decoder9.U79.ZN ) ) ;
not ( 
    .O1 ( config0_decoder9.n39 ) ,
    .IN ( masks_hold_reg_7_4 ) ) ;
or ( 
    .Z ( config0_decoder9.U69.AB ) ,
    .I0 ( config0_decoder9.n49 ) ,
    .I1 ( config0_decoder9.n47 ) ) ;
and ( 
    .Z ( config0_decoder9.U69.ZN ) ,
    .I0 ( config0_decoder9.U69.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_44 ) ,
    .IN ( config0_decoder9.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U20.AB ) ,
    .I0 ( config0_decoder9.n57 ) ,
    .I1 ( config0_decoder9.n53 ) ) ;
and ( 
    .Z ( config0_decoder9.U20.ZN ) ,
    .I0 ( config0_decoder9.U20.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_48 ) ,
    .IN ( config0_decoder9.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n60 ) ,
    .I0 ( config0_decoder9.n42 ) ,
    .I1 ( config0_decoder9.n41 ) ) ;
or ( 
    .Z ( config0_decoder9.U4.AB ) ,
    .I0 ( config0_decoder9.n58 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U4.ZN ) ,
    .I0 ( config0_decoder9.U4.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_22 ) ,
    .IN ( config0_decoder9.U4.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n56 ) ,
    .I0 ( config0_decoder9.n41 ) ,
    .I1 ( config0_decoder9.n39 ) ,
    .I2 ( masks_hold_reg_7_3 ) ) ;
or ( 
    .Z ( config0_decoder9.U43.AB ) ,
    .I0 ( config0_decoder9.n58 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U43.ZN ) ,
    .I0 ( config0_decoder9.U43.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_21 ) ,
    .IN ( config0_decoder9.U43.ZN ) ) ;
and ( 
    .Z ( config0_decoder9.n40 ) ,
    .I0 ( masks_hold_reg_7_3 ) ,
    .I1 ( masks_hold_reg_7_2 ) ) ;
nor ( 
    .Z ( config0_decoder9.n46 ) ,
    .I0 ( config0_decoder9.n45 ) ,
    .I1 ( masks_hold_reg_7_5 ) ) ;
not ( 
    .O1 ( config0_decoder9.n51 ) ,
    .IN ( masks_hold_reg_7_1 ) ) ;
or ( 
    .Z ( config0_decoder9.U14.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n58 ) ) ;
and ( 
    .Z ( config0_decoder9.U14.ZN ) ,
    .I0 ( config0_decoder9.U14.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_5 ) ,
    .IN ( config0_decoder9.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n53 ) ,
    .I0 ( config0_decoder9.n38 ) ,
    .I1 ( config0_decoder9.n41 ) ) ;
nand ( 
    .Z ( config0_decoder9.n62 ) ,
    .I0 ( config0_decoder9.n35 ) ,
    .I1 ( config0_decoder9.n51 ) ) ;
nand ( 
    .Z ( config0_decoder9.n47 ) ,
    .I0 ( masks_hold_reg_7_4 ) ,
    .I1 ( config0_decoder9.n41 ) ,
    .I2 ( masks_hold_reg_7_3 ) ) ;
or ( 
    .Z ( config0_decoder9.U42.AB ) ,
    .I0 ( config0_decoder9.n58 ) ,
    .I1 ( config0_decoder9.n48 ) ) ;
and ( 
    .Z ( config0_decoder9.U42.ZN ) ,
    .I0 ( config0_decoder9.U42.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_37 ) ,
    .IN ( config0_decoder9.U42.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U70.AB ) ,
    .I0 ( config0_decoder9.n50 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U70.ZN ) ,
    .I0 ( config0_decoder9.U70.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_46 ) ,
    .IN ( config0_decoder9.U70.ZN ) ) ;
nor ( 
    .Z ( config0_decoder9.n38 ) ,
    .I0 ( masks_hold_reg_7_3 ) ,
    .I1 ( masks_hold_reg_7_4 ) ) ;
or ( 
    .Z ( config0_decoder9.U18.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n56 ) ) ;
and ( 
    .Z ( config0_decoder9.U18.ZN ) ,
    .I0 ( config0_decoder9.U18.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_3 ) ,
    .IN ( config0_decoder9.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U15.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n60 ) ) ;
and ( 
    .Z ( config0_decoder9.U15.ZN ) ,
    .I0 ( config0_decoder9.U15.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_7 ) ,
    .IN ( config0_decoder9.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n43 ) ,
    .I0 ( config0_decoder9.n37 ) ,
    .I1 ( config0_decoder9.n51 ) ) ;
or ( 
    .Z ( config0_decoder9.U85.AB ) ,
    .I0 ( config0_decoder9.n48 ) ,
    .I1 ( config0_decoder9.n47 ) ) ;
and ( 
    .Z ( config0_decoder9.U85.ZN ) ,
    .I0 ( config0_decoder9.U85.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_43 ) ,
    .IN ( config0_decoder9.U85.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n59 ) ,
    .I0 ( masks_hold_reg_7_1 ) ,
    .I1 ( config0_decoder9.n35 ) ) ;
or ( 
    .Z ( config0_decoder9.U45.AB ) ,
    .I0 ( config0_decoder9.n62 ) ,
    .I1 ( config0_decoder9.n47 ) ) ;
and ( 
    .Z ( config0_decoder9.U45.ZN ) ,
    .I0 ( config0_decoder9.U45.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_11 ) ,
    .IN ( config0_decoder9.U45.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U71.AB ) ,
    .I0 ( config0_decoder9.n56 ) ,
    .I1 ( config0_decoder9.n55 ) ) ;
and ( 
    .Z ( config0_decoder9.U71.ZN ) ,
    .I0 ( config0_decoder9.U71.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_51 ) ,
    .IN ( config0_decoder9.U71.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n57 ) ,
    .I0 ( masks_hold_reg_7_1 ) ,
    .I1 ( config0_decoder9.n52 ) ) ;
or ( 
    .Z ( config0_decoder9.U19.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n54 ) ) ;
and ( 
    .Z ( config0_decoder9.U19.ZN ) ,
    .I0 ( config0_decoder9.U19.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_2 ) ,
    .IN ( config0_decoder9.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U16.AB ) ,
    .I0 ( config0_decoder9.n59 ) ,
    .I1 ( config0_decoder9.n58 ) ) ;
and ( 
    .Z ( config0_decoder9.U16.ZN ) ,
    .I0 ( config0_decoder9.U16.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_6 ) ,
    .IN ( config0_decoder9.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U36.AB ) ,
    .I0 ( config0_decoder9.n58 ) ,
    .I1 ( config0_decoder9.n49 ) ) ;
and ( 
    .Z ( config0_decoder9.U36.ZN ) ,
    .I0 ( config0_decoder9.U36.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_38 ) ,
    .IN ( config0_decoder9.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U1.AB ) ,
    .I0 ( config0_decoder9.n47 ) ,
    .I1 ( config0_decoder9.n44 ) ) ;
and ( 
    .Z ( config0_decoder9.U1.ZN ) ,
    .I0 ( config0_decoder9.U1.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_28 ) ,
    .IN ( config0_decoder9.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder9.U84.AB ) ,
    .I0 ( config0_decoder9.n56 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U84.ZN ) ,
    .I0 ( config0_decoder9.U84.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_19 ) ,
    .IN ( config0_decoder9.U84.ZN ) ) ;
nand ( 
    .Z ( config0_decoder9.n54 ) ,
    .I0 ( config0_decoder9.n38 ) ,
    .I1 ( masks_hold_reg_7_2 ) ) ;
or ( 
    .Z ( config0_decoder9.U44.AB ) ,
    .I0 ( config0_decoder9.n53 ) ,
    .I1 ( config0_decoder9.n43 ) ) ;
and ( 
    .Z ( config0_decoder9.U44.ZN ) ,
    .I0 ( config0_decoder9.U44.AB ) ,
    .I1 ( config0_decoder9.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_8_15 ) ,
    .IN ( config0_decoder9.U44.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U28.AB ) ,
    .I0 ( config0_decoder8.n40 ) ,
    .I1 ( masks_hold_reg_6_3 ) ) ;
and ( 
    .Z ( config0_decoder8.U28.ZN ) ,
    .I0 ( config0_decoder8.U28.AB ) ,
    .I1 ( config0_decoder8.n52 ) ) ;
not ( 
    .O1 ( config0_decoder8.n1 ) ,
    .IN ( config0_decoder8.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U76.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n47 ) ) ;
and ( 
    .Z ( config0_decoder8.U76.ZN ) ,
    .I0 ( config0_decoder8.U76.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_11 ) ,
    .IN ( config0_decoder8.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U60.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n59 ) ) ;
and ( 
    .Z ( config0_decoder8.U60.ZN ) ,
    .I0 ( config0_decoder8.U60.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_10 ) ,
    .IN ( config0_decoder8.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U17.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n54 ) ) ;
and ( 
    .Z ( config0_decoder8.U17.ZN ) ,
    .I0 ( config0_decoder8.U17.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_2 ) ,
    .IN ( config0_decoder8.U17.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n57 ) ,
    .I0 ( masks_hold_reg_6_0 ) ,
    .I1 ( config0_decoder8.n52 ) ) ;
or ( 
    .Z ( config0_decoder8.U87.AB ) ,
    .I0 ( config0_decoder8.n57 ) ,
    .I1 ( config0_decoder8.n54 ) ) ;
and ( 
    .Z ( config0_decoder8.U87.ZN ) ,
    .I0 ( config0_decoder8.U87.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_50 ) ,
    .IN ( config0_decoder8.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U57.AB ) ,
    .I0 ( config0_decoder8.n56 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U57.ZN ) ,
    .I0 ( config0_decoder8.U57.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_36 ) ,
    .IN ( config0_decoder8.U57.ZN ) ) ;
not ( 
    .O1 ( config0_decoder8.n36 ) ,
    .IN ( masks_hold_reg_6_4 ) ) ;
or ( 
    .Z ( config0_decoder8.U77.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U77.ZN ) ,
    .I0 ( config0_decoder8.U77.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_41 ) ,
    .IN ( config0_decoder8.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U67.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n47 ) ) ;
and ( 
    .Z ( config0_decoder8.U67.ZN ) ,
    .I0 ( config0_decoder8.U67.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_12 ) ,
    .IN ( config0_decoder8.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U10.AB ) ,
    .I0 ( config0_decoder8.n50 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U10.ZN ) ,
    .I0 ( config0_decoder8.U10.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_30 ) ,
    .IN ( config0_decoder8.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n44 ) ,
    .I0 ( config0_decoder8.n37 ) ,
    .I1 ( masks_hold_reg_6_0 ) ) ;
or ( 
    .Z ( config0_decoder8.U26.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n56 ) ) ;
and ( 
    .Z ( config0_decoder8.U26.ZN ) ,
    .I0 ( config0_decoder8.U26.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_3 ) ,
    .IN ( config0_decoder8.U26.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n43 ) ,
    .I0 ( config0_decoder8.n37 ) ,
    .I1 ( config0_decoder8.n51 ) ) ;
or ( 
    .Z ( config0_decoder8.U86.AB ) ,
    .I0 ( config0_decoder8.n57 ) ,
    .I1 ( config0_decoder8.n56 ) ) ;
and ( 
    .Z ( config0_decoder8.U86.ZN ) ,
    .I0 ( config0_decoder8.U86.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_52 ) ,
    .IN ( config0_decoder8.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U58.AB ) ,
    .I0 ( config0_decoder8.n56 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U58.ZN ) ,
    .I0 ( config0_decoder8.U58.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_20 ) ,
    .IN ( config0_decoder8.U58.ZN ) ) ;
not ( 
    .O1 ( config0_decoder8.n45 ) ,
    .IN ( masks_hold_reg_6_5 ) ) ;
or ( 
    .Z ( config0_decoder8.U74.AB ) ,
    .I0 ( config0_decoder8.n58 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U74.ZN ) ,
    .I0 ( config0_decoder8.U74.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_21 ) ,
    .IN ( config0_decoder8.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U66.AB ) ,
    .I0 ( config0_decoder8.n60 ) ,
    .I1 ( config0_decoder8.n59 ) ) ;
and ( 
    .Z ( config0_decoder8.U66.ZN ) ,
    .I0 ( config0_decoder8.U66.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_8 ) ,
    .IN ( config0_decoder8.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U11.AB ) ,
    .I0 ( config0_decoder8.n53 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U11.ZN ) ,
    .I0 ( config0_decoder8.U11.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_31 ) ,
    .IN ( config0_decoder8.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder8.n35 ) ,
    .I0 ( masks_hold_reg_6_4 ) ,
    .I1 ( masks_hold_reg_6_5 ) ) ;
nand ( 
    .Z ( config0_decoder8.n63 ) ,
    .I0 ( masks_hold_reg_6_1 ) ,
    .I1 ( config0_decoder8.n42 ) ) ;
or ( 
    .Z ( config0_decoder8.U25.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n58 ) ) ;
and ( 
    .Z ( config0_decoder8.U25.ZN ) ,
    .I0 ( config0_decoder8.U25.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_6 ) ,
    .IN ( config0_decoder8.U25.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n62 ) ,
    .I0 ( config0_decoder8.n35 ) ,
    .I1 ( config0_decoder8.n51 ) ) ;
or ( 
    .Z ( config0_decoder8.U81.AB ) ,
    .I0 ( config0_decoder8.n60 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U81.ZN ) ,
    .I0 ( config0_decoder8.U81.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_23 ) ,
    .IN ( config0_decoder8.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U59.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n50 ) ) ;
and ( 
    .Z ( config0_decoder8.U59.ZN ) ,
    .I0 ( config0_decoder8.U59.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_14 ) ,
    .IN ( config0_decoder8.U59.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U49.AB ) ,
    .I0 ( config0_decoder8.n50 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U49.ZN ) ,
    .I0 ( config0_decoder8.U49.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_46 ) ,
    .IN ( config0_decoder8.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U75.AB ) ,
    .I0 ( config0_decoder8.n53 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U75.ZN ) ,
    .I0 ( config0_decoder8.U75.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_15 ) ,
    .IN ( config0_decoder8.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U65.AB ) ,
    .I0 ( config0_decoder8.n58 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U65.ZN ) ,
    .I0 ( config0_decoder8.U65.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_22 ) ,
    .IN ( config0_decoder8.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U12.AB ) ,
    .I0 ( config0_decoder8.n53 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U12.ZN ) ,
    .I0 ( config0_decoder8.U12.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_16 ) ,
    .IN ( config0_decoder8.U12.ZN ) ) ;
nor ( 
    .Z ( config0_decoder8.n37 ) ,
    .I0 ( config0_decoder8.n36 ) ,
    .I1 ( masks_hold_reg_6_5 ) ) ;
nand ( 
    .Z ( config0_decoder8.n54 ) ,
    .I0 ( config0_decoder8.n38 ) ,
    .I1 ( masks_hold_reg_6_1 ) ) ;
nand ( 
    .Z ( config0_decoder8.n56 ) ,
    .I0 ( config0_decoder8.n41 ) ,
    .I1 ( config0_decoder8.n39 ) ,
    .I2 ( masks_hold_reg_6_2 ) ) ;
or ( 
    .Z ( config0_decoder8.U80.AB ) ,
    .I0 ( config0_decoder8.n60 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U80.ZN ) ,
    .I0 ( config0_decoder8.U80.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_39 ) ,
    .IN ( config0_decoder8.U80.ZN ) ) ;
and ( 
    .Z ( config0_decoder8.n40 ) ,
    .I0 ( masks_hold_reg_6_2 ) ,
    .I1 ( masks_hold_reg_6_1 ) ) ;
or ( 
    .Z ( config0_decoder8.U64.AB ) ,
    .I0 ( config0_decoder8.n58 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U64.ZN ) ,
    .I0 ( config0_decoder8.U64.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_38 ) ,
    .IN ( config0_decoder8.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U13.AB ) ,
    .I0 ( config0_decoder8.n54 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U13.ZN ) ,
    .I0 ( config0_decoder8.U13.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_18 ) ,
    .IN ( config0_decoder8.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n49 ) ,
    .I0 ( config0_decoder8.n46 ) ,
    .I1 ( masks_hold_reg_6_0 ) ) ;
or ( 
    .Z ( config0_decoder8.U83.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n50 ) ) ;
and ( 
    .Z ( config0_decoder8.U83.ZN ) ,
    .I0 ( config0_decoder8.U83.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_13 ) ,
    .IN ( config0_decoder8.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U50.AB ) ,
    .I0 ( config0_decoder8.n49 ) ,
    .I1 ( config0_decoder8.n47 ) ) ;
and ( 
    .Z ( config0_decoder8.U50.ZN ) ,
    .I0 ( config0_decoder8.U50.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_44 ) ,
    .IN ( config0_decoder8.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n47 ) ,
    .I0 ( masks_hold_reg_6_3 ) ,
    .I1 ( config0_decoder8.n41 ) ,
    .I2 ( masks_hold_reg_6_2 ) ) ;
or ( 
    .Z ( config0_decoder8.U82.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n62 ) ) ;
and ( 
    .Z ( config0_decoder8.U82.ZN ) ,
    .I0 ( config0_decoder8.U82.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_9 ) ,
    .IN ( config0_decoder8.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U51.AB ) ,
    .I0 ( config0_decoder8.n50 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U51.ZN ) ,
    .I0 ( config0_decoder8.U51.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_45 ) ,
    .IN ( config0_decoder8.U51.ZN ) ) ;
not ( 
    .O1 ( config0_decoder8.n51 ) ,
    .IN ( masks_hold_reg_6_0 ) ) ;
or ( 
    .Z ( config0_decoder8.U78.AB ) ,
    .I0 ( config0_decoder8.n47 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U78.ZN ) ,
    .I0 ( config0_decoder8.U78.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_27 ) ,
    .IN ( config0_decoder8.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n59 ) ,
    .I0 ( masks_hold_reg_6_0 ) ,
    .I1 ( config0_decoder8.n35 ) ) ;
nand ( 
    .Z ( config0_decoder8.n60 ) ,
    .I0 ( config0_decoder8.n42 ) ,
    .I1 ( config0_decoder8.n41 ) ) ;
or ( 
    .Z ( config0_decoder8.U52.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n58 ) ) ;
and ( 
    .Z ( config0_decoder8.U52.ZN ) ,
    .I0 ( config0_decoder8.U52.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_5 ) ,
    .IN ( config0_decoder8.U52.ZN ) ) ;
nor ( 
    .Z ( config0_decoder8.n38 ) ,
    .I0 ( masks_hold_reg_6_2 ) ,
    .I1 ( masks_hold_reg_6_3 ) ) ;
or ( 
    .Z ( config0_decoder8.U79.AB ) ,
    .I0 ( config0_decoder8.n56 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U79.ZN ) ,
    .I0 ( config0_decoder8.U79.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_35 ) ,
    .IN ( config0_decoder8.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U72.AB ) ,
    .I0 ( config0_decoder8.n58 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U72.ZN ) ,
    .I0 ( config0_decoder8.U72.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_37 ) ,
    .IN ( config0_decoder8.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U69.AB ) ,
    .I0 ( config0_decoder8.n50 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U69.ZN ) ,
    .I0 ( config0_decoder8.U69.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_29 ) ,
    .IN ( config0_decoder8.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U20.AB ) ,
    .I0 ( config0_decoder8.n56 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U20.ZN ) ,
    .I0 ( config0_decoder8.U20.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_19 ) ,
    .IN ( config0_decoder8.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U9.AB ) ,
    .I0 ( config0_decoder8.n47 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U9.ZN ) ,
    .I0 ( config0_decoder8.U9.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_28 ) ,
    .IN ( config0_decoder8.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n53 ) ,
    .I0 ( config0_decoder8.n38 ) ,
    .I1 ( config0_decoder8.n41 ) ) ;
or ( 
    .Z ( config0_decoder8.U53.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n54 ) ) ;
and ( 
    .Z ( config0_decoder8.U53.ZN ) ,
    .I0 ( config0_decoder8.U53.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_1 ) ,
    .IN ( config0_decoder8.U53.ZN ) ) ;
nor ( 
    .Z ( config0_decoder8.n42 ) ,
    .I0 ( config0_decoder8.n39 ) ,
    .I1 ( masks_hold_reg_6_2 ) ) ;
or ( 
    .Z ( config0_decoder8.U73.AB ) ,
    .I0 ( config0_decoder8.n54 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U73.ZN ) ,
    .I0 ( config0_decoder8.U73.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_17 ) ,
    .IN ( config0_decoder8.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U68.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U68.ZN ) ,
    .I0 ( config0_decoder8.U68.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_42 ) ,
    .IN ( config0_decoder8.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U63.AB ) ,
    .I0 ( config0_decoder8.n54 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U63.ZN ) ,
    .I0 ( config0_decoder8.U63.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_34 ) ,
    .IN ( config0_decoder8.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U14.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n56 ) ) ;
and ( 
    .Z ( config0_decoder8.U14.ZN ) ,
    .I0 ( config0_decoder8.U14.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_4 ) ,
    .IN ( config0_decoder8.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n55 ) ,
    .I0 ( config0_decoder8.n52 ) ,
    .I1 ( config0_decoder8.n51 ) ) ;
nor ( 
    .Z ( config0_decoder8.n52 ) ,
    .I0 ( config0_decoder8.n45 ) ,
    .I1 ( config0_decoder8.n36 ) ) ;
or ( 
    .Z ( config0_decoder8.U54.AB ) ,
    .I0 ( config0_decoder8.n55 ) ,
    .I1 ( config0_decoder8.n53 ) ) ;
and ( 
    .Z ( config0_decoder8.U54.ZN ) ,
    .I0 ( config0_decoder8.U54.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_47 ) ,
    .IN ( config0_decoder8.U54.ZN ) ) ;
nor ( 
    .Z ( config0_decoder8.n46 ) ,
    .I0 ( config0_decoder8.n45 ) ,
    .I1 ( masks_hold_reg_6_4 ) ) ;
or ( 
    .Z ( config0_decoder8.U70.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n43 ) ) ;
and ( 
    .Z ( config0_decoder8.U70.ZN ) ,
    .I0 ( config0_decoder8.U70.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_25 ) ,
    .IN ( config0_decoder8.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U62.AB ) ,
    .I0 ( config0_decoder8.n63 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U62.ZN ) ,
    .I0 ( config0_decoder8.U62.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_26 ) ,
    .IN ( config0_decoder8.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U18.AB ) ,
    .I0 ( config0_decoder8.n57 ) ,
    .I1 ( config0_decoder8.n53 ) ) ;
and ( 
    .Z ( config0_decoder8.U18.ZN ) ,
    .I0 ( config0_decoder8.U18.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_48 ) ,
    .IN ( config0_decoder8.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U15.AB ) ,
    .I0 ( config0_decoder8.n62 ) ,
    .I1 ( config0_decoder8.n60 ) ) ;
and ( 
    .Z ( config0_decoder8.U15.ZN ) ,
    .I0 ( config0_decoder8.U15.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_7 ) ,
    .IN ( config0_decoder8.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n58 ) ,
    .I0 ( config0_decoder8.n40 ) ,
    .I1 ( config0_decoder8.n39 ) ) ;
or ( 
    .Z ( config0_decoder8.U85.AB ) ,
    .I0 ( config0_decoder8.n56 ) ,
    .I1 ( config0_decoder8.n55 ) ) ;
and ( 
    .Z ( config0_decoder8.U85.ZN ) ,
    .I0 ( config0_decoder8.U85.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_51 ) ,
    .IN ( config0_decoder8.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U55.AB ) ,
    .I0 ( config0_decoder8.n60 ) ,
    .I1 ( config0_decoder8.n44 ) ) ;
and ( 
    .Z ( config0_decoder8.U55.ZN ) ,
    .I0 ( config0_decoder8.U55.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_24 ) ,
    .IN ( config0_decoder8.U55.ZN ) ) ;
not ( 
    .O1 ( config0_decoder8.n39 ) ,
    .IN ( masks_hold_reg_6_3 ) ) ;
or ( 
    .Z ( config0_decoder8.U71.AB ) ,
    .I0 ( config0_decoder8.n54 ) ,
    .I1 ( config0_decoder8.n48 ) ) ;
and ( 
    .Z ( config0_decoder8.U71.ZN ) ,
    .I0 ( config0_decoder8.U71.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_33 ) ,
    .IN ( config0_decoder8.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U61.AB ) ,
    .I0 ( config0_decoder8.n60 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U61.ZN ) ,
    .I0 ( config0_decoder8.U61.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_40 ) ,
    .IN ( config0_decoder8.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U19.AB ) ,
    .I0 ( config0_decoder8.n55 ) ,
    .I1 ( config0_decoder8.n54 ) ) ;
and ( 
    .Z ( config0_decoder8.U19.ZN ) ,
    .I0 ( config0_decoder8.U19.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_49 ) ,
    .IN ( config0_decoder8.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U16.AB ) ,
    .I0 ( config0_decoder8.n59 ) ,
    .I1 ( config0_decoder8.n53 ) ) ;
and ( 
    .Z ( config0_decoder8.U16.ZN ) ,
    .I0 ( config0_decoder8.U16.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_0 ) ,
    .IN ( config0_decoder8.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder8.n50 ) ,
    .I0 ( config0_decoder8.n40 ) ,
    .I1 ( masks_hold_reg_6_3 ) ) ;
nand ( 
    .Z ( config0_decoder8.n48 ) ,
    .I0 ( config0_decoder8.n46 ) ,
    .I1 ( config0_decoder8.n51 ) ) ;
or ( 
    .Z ( config0_decoder8.U84.AB ) ,
    .I0 ( config0_decoder8.n48 ) ,
    .I1 ( config0_decoder8.n47 ) ) ;
and ( 
    .Z ( config0_decoder8.U84.ZN ) ,
    .I0 ( config0_decoder8.U84.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_43 ) ,
    .IN ( config0_decoder8.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder8.U56.AB ) ,
    .I0 ( config0_decoder8.n53 ) ,
    .I1 ( config0_decoder8.n49 ) ) ;
and ( 
    .Z ( config0_decoder8.U56.ZN ) ,
    .I0 ( config0_decoder8.U56.AB ) ,
    .I1 ( config0_decoder8.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_7_32 ) ,
    .IN ( config0_decoder8.U56.ZN ) ) ;
not ( 
    .O1 ( config0_decoder8.n41 ) ,
    .IN ( masks_hold_reg_6_1 ) ) ;
or ( 
    .Z ( config0_decoder3.U55.AB ) ,
    .I0 ( config0_decoder3.n40 ) ,
    .I1 ( masks_hold_reg_2_9 ) ) ;
and ( 
    .Z ( config0_decoder3.U55.ZN ) ,
    .I0 ( config0_decoder3.U55.AB ) ,
    .I1 ( config0_decoder3.n52 ) ) ;
not ( 
    .O1 ( config0_decoder3.n1 ) ,
    .IN ( config0_decoder3.U55.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U44.AB ) ,
    .I0 ( config0_decoder3.n58 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U44.ZN ) ,
    .I0 ( config0_decoder3.U44.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_37 ) ,
    .IN ( config0_decoder3.U44.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U76.AB ) ,
    .I0 ( config0_decoder3.n50 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U76.ZN ) ,
    .I0 ( config0_decoder3.U76.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_46 ) ,
    .IN ( config0_decoder3.U76.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n44 ) ,
    .I0 ( config0_decoder3.n37 ) ,
    .I1 ( n86 ) ) ;
or ( 
    .Z ( config0_decoder3.U17.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n58 ) ) ;
and ( 
    .Z ( config0_decoder3.U17.ZN ) ,
    .I0 ( config0_decoder3.U17.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_6 ) ,
    .IN ( config0_decoder3.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U37.AB ) ,
    .I0 ( config0_decoder3.n58 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U37.ZN ) ,
    .I0 ( config0_decoder3.U37.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_38 ) ,
    .IN ( config0_decoder3.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U87.AB ) ,
    .I0 ( config0_decoder3.n57 ) ,
    .I1 ( config0_decoder3.n54 ) ) ;
and ( 
    .Z ( config0_decoder3.U87.ZN ) ,
    .I0 ( config0_decoder3.U87.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_50 ) ,
    .IN ( config0_decoder3.U87.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n59 ) ,
    .I0 ( n86 ) ,
    .I1 ( config0_decoder3.n35 ) ) ;
or ( 
    .Z ( config0_decoder3.U47.AB ) ,
    .I0 ( config0_decoder3.n53 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U47.ZN ) ,
    .I0 ( config0_decoder3.U47.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_15 ) ,
    .IN ( config0_decoder3.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U77.AB ) ,
    .I0 ( config0_decoder3.n49 ) ,
    .I1 ( config0_decoder3.n47 ) ) ;
and ( 
    .Z ( config0_decoder3.U77.ZN ) ,
    .I0 ( config0_decoder3.U77.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_44 ) ,
    .IN ( config0_decoder3.U77.ZN ) ) ;
nor ( 
    .Z ( config0_decoder3.n42 ) ,
    .I0 ( config0_decoder3.n39 ) ,
    .I1 ( masks_hold_reg_2_8 ) ) ;
nand ( 
    .Z ( config0_decoder3.n62 ) ,
    .I0 ( config0_decoder3.n35 ) ,
    .I1 ( config0_decoder3.n51 ) ) ;
or ( 
    .Z ( config0_decoder3.U34.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n50 ) ) ;
and ( 
    .Z ( config0_decoder3.U34.ZN ) ,
    .I0 ( config0_decoder3.U34.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_14 ) ,
    .IN ( config0_decoder3.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U3.AB ) ,
    .I0 ( config0_decoder3.n53 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U3.ZN ) ,
    .I0 ( config0_decoder3.U3.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_31 ) ,
    .IN ( config0_decoder3.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U86.AB ) ,
    .I0 ( config0_decoder3.n57 ) ,
    .I1 ( config0_decoder3.n56 ) ) ;
and ( 
    .Z ( config0_decoder3.U86.ZN ) ,
    .I0 ( config0_decoder3.U86.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_52 ) ,
    .IN ( config0_decoder3.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n47 ) ,
    .I0 ( masks_hold_reg_2_9 ) ,
    .I1 ( config0_decoder3.n41 ) ,
    .I2 ( masks_hold_reg_2_8 ) ) ;
or ( 
    .Z ( config0_decoder3.U46.AB ) ,
    .I0 ( config0_decoder3.n54 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U46.ZN ) ,
    .I0 ( config0_decoder3.U46.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_17 ) ,
    .IN ( config0_decoder3.U46.ZN ) ) ;
not ( 
    .O1 ( config0_decoder3.n36 ) ,
    .IN ( masks_hold_reg_2_10 ) ) ;
nor ( 
    .Z ( config0_decoder3.n38 ) ,
    .I0 ( masks_hold_reg_2_8 ) ,
    .I1 ( masks_hold_reg_2_9 ) ) ;
nand ( 
    .Z ( config0_decoder3.n53 ) ,
    .I0 ( config0_decoder3.n38 ) ,
    .I1 ( config0_decoder3.n41 ) ) ;
or ( 
    .Z ( config0_decoder3.U38.AB ) ,
    .I0 ( config0_decoder3.n54 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U38.ZN ) ,
    .I0 ( config0_decoder3.U38.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_18 ) ,
    .IN ( config0_decoder3.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U35.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U35.ZN ) ,
    .I0 ( config0_decoder3.U35.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_26 ) ,
    .IN ( config0_decoder3.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U2.AB ) ,
    .I0 ( config0_decoder3.n50 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U2.ZN ) ,
    .I0 ( config0_decoder3.U2.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_30 ) ,
    .IN ( config0_decoder3.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U81.AB ) ,
    .I0 ( config0_decoder3.n60 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U81.ZN ) ,
    .I0 ( config0_decoder3.U81.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_40 ) ,
    .IN ( config0_decoder3.U81.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n49 ) ,
    .I0 ( config0_decoder3.n46 ) ,
    .I1 ( n86 ) ) ;
or ( 
    .Z ( config0_decoder3.U49.AB ) ,
    .I0 ( config0_decoder3.n47 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U49.ZN ) ,
    .I0 ( config0_decoder3.U49.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_27 ) ,
    .IN ( config0_decoder3.U49.ZN ) ) ;
not ( 
    .O1 ( config0_decoder3.n45 ) ,
    .IN ( masks_hold_reg_1_0 ) ) ;
nand ( 
    .Z ( config0_decoder3.n50 ) ,
    .I0 ( config0_decoder3.n40 ) ,
    .I1 ( masks_hold_reg_2_9 ) ) ;
nand ( 
    .Z ( config0_decoder3.n60 ) ,
    .I0 ( config0_decoder3.n42 ) ,
    .I1 ( config0_decoder3.n41 ) ) ;
or ( 
    .Z ( config0_decoder3.U39.AB ) ,
    .I0 ( config0_decoder3.n60 ) ,
    .I1 ( config0_decoder3.n59 ) ) ;
and ( 
    .Z ( config0_decoder3.U39.ZN ) ,
    .I0 ( config0_decoder3.U39.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_8 ) ,
    .IN ( config0_decoder3.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U32.AB ) ,
    .I0 ( config0_decoder3.n56 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U32.ZN ) ,
    .I0 ( config0_decoder3.U32.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_36 ) ,
    .IN ( config0_decoder3.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U29.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n58 ) ) ;
and ( 
    .Z ( config0_decoder3.U29.ZN ) ,
    .I0 ( config0_decoder3.U29.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_5 ) ,
    .IN ( config0_decoder3.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U80.AB ) ,
    .I0 ( config0_decoder3.n55 ) ,
    .I1 ( config0_decoder3.n53 ) ) ;
and ( 
    .Z ( config0_decoder3.U80.ZN ) ,
    .I0 ( config0_decoder3.U80.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_47 ) ,
    .IN ( config0_decoder3.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U48.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n47 ) ) ;
and ( 
    .Z ( config0_decoder3.U48.ZN ) ,
    .I0 ( config0_decoder3.U48.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_11 ) ,
    .IN ( config0_decoder3.U48.ZN ) ) ;
not ( 
    .O1 ( config0_decoder3.n51 ) ,
    .IN ( n86 ) ) ;
nand ( 
    .Z ( config0_decoder3.n58 ) ,
    .I0 ( config0_decoder3.n40 ) ,
    .I1 ( config0_decoder3.n39 ) ) ;
or ( 
    .Z ( config0_decoder3.U33.AB ) ,
    .I0 ( config0_decoder3.n53 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U33.ZN ) ,
    .I0 ( config0_decoder3.U33.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_16 ) ,
    .IN ( config0_decoder3.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U28.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n59 ) ) ;
and ( 
    .Z ( config0_decoder3.U28.ZN ) ,
    .I0 ( config0_decoder3.U28.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_10 ) ,
    .IN ( config0_decoder3.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U83.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U83.ZN ) ,
    .I0 ( config0_decoder3.U83.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_41 ) ,
    .IN ( config0_decoder3.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U50.AB ) ,
    .I0 ( config0_decoder3.n56 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U50.ZN ) ,
    .I0 ( config0_decoder3.U50.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_35 ) ,
    .IN ( config0_decoder3.U50.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U30.AB ) ,
    .I0 ( config0_decoder3.n60 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U30.ZN ) ,
    .I0 ( config0_decoder3.U30.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_24 ) ,
    .IN ( config0_decoder3.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U22.AB ) ,
    .I0 ( config0_decoder3.n55 ) ,
    .I1 ( config0_decoder3.n54 ) ) ;
and ( 
    .Z ( config0_decoder3.U22.ZN ) ,
    .I0 ( config0_decoder3.U22.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_49 ) ,
    .IN ( config0_decoder3.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U82.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U82.ZN ) ,
    .I0 ( config0_decoder3.U82.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_42 ) ,
    .IN ( config0_decoder3.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U51.AB ) ,
    .I0 ( config0_decoder3.n60 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U51.ZN ) ,
    .I0 ( config0_decoder3.U51.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_39 ) ,
    .IN ( config0_decoder3.U51.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U41.AB ) ,
    .I0 ( config0_decoder3.n50 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U41.ZN ) ,
    .I0 ( config0_decoder3.U41.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_29 ) ,
    .IN ( config0_decoder3.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U78.AB ) ,
    .I0 ( config0_decoder3.n50 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U78.ZN ) ,
    .I0 ( config0_decoder3.U78.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_45 ) ,
    .IN ( config0_decoder3.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U31.AB ) ,
    .I0 ( config0_decoder3.n53 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U31.ZN ) ,
    .I0 ( config0_decoder3.U31.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_32 ) ,
    .IN ( config0_decoder3.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U21.AB ) ,
    .I0 ( config0_decoder3.n57 ) ,
    .I1 ( config0_decoder3.n53 ) ) ;
and ( 
    .Z ( config0_decoder3.U21.ZN ) ,
    .I0 ( config0_decoder3.U21.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_48 ) ,
    .IN ( config0_decoder3.U21.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U5.AB ) ,
    .I0 ( config0_decoder3.n60 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U5.ZN ) ,
    .I0 ( config0_decoder3.U5.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_23 ) ,
    .IN ( config0_decoder3.U5.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U52.AB ) ,
    .I0 ( config0_decoder3.n56 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U52.ZN ) ,
    .I0 ( config0_decoder3.U52.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_19 ) ,
    .IN ( config0_decoder3.U52.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U40.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n47 ) ) ;
and ( 
    .Z ( config0_decoder3.U40.ZN ) ,
    .I0 ( config0_decoder3.U40.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_12 ) ,
    .IN ( config0_decoder3.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U79.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n54 ) ) ;
and ( 
    .Z ( config0_decoder3.U79.ZN ) ,
    .I0 ( config0_decoder3.U79.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_1 ) ,
    .IN ( config0_decoder3.U79.ZN ) ) ;
nor ( 
    .Z ( config0_decoder3.n37 ) ,
    .I0 ( config0_decoder3.n36 ) ,
    .I1 ( masks_hold_reg_1_0 ) ) ;
nor ( 
    .Z ( config0_decoder3.n35 ) ,
    .I0 ( masks_hold_reg_2_10 ) ,
    .I1 ( masks_hold_reg_1_0 ) ) ;
or ( 
    .Z ( config0_decoder3.U20.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n54 ) ) ;
and ( 
    .Z ( config0_decoder3.U20.ZN ) ,
    .I0 ( config0_decoder3.U20.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_2 ) ,
    .IN ( config0_decoder3.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n43 ) ,
    .I0 ( config0_decoder3.n37 ) ,
    .I1 ( config0_decoder3.n51 ) ) ;
or ( 
    .Z ( config0_decoder3.U4.AB ) ,
    .I0 ( config0_decoder3.n58 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U4.ZN ) ,
    .I0 ( config0_decoder3.U4.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_22 ) ,
    .IN ( config0_decoder3.U4.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U53.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n62 ) ) ;
and ( 
    .Z ( config0_decoder3.U53.ZN ) ,
    .I0 ( config0_decoder3.U53.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_9 ) ,
    .IN ( config0_decoder3.U53.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U43.AB ) ,
    .I0 ( config0_decoder3.n54 ) ,
    .I1 ( config0_decoder3.n48 ) ) ;
and ( 
    .Z ( config0_decoder3.U43.ZN ) ,
    .I0 ( config0_decoder3.U43.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_33 ) ,
    .IN ( config0_decoder3.U43.ZN ) ) ;
and ( 
    .Z ( config0_decoder3.n40 ) ,
    .I0 ( masks_hold_reg_2_8 ) ,
    .I1 ( masks_hold_reg_2_7 ) ) ;
not ( 
    .O1 ( config0_decoder3.n41 ) ,
    .IN ( masks_hold_reg_2_7 ) ) ;
nand ( 
    .Z ( config0_decoder3.n63 ) ,
    .I0 ( masks_hold_reg_2_7 ) ,
    .I1 ( config0_decoder3.n42 ) ) ;
nor ( 
    .Z ( config0_decoder3.n52 ) ,
    .I0 ( config0_decoder3.n45 ) ,
    .I1 ( config0_decoder3.n36 ) ) ;
nand ( 
    .Z ( config0_decoder3.n48 ) ,
    .I0 ( config0_decoder3.n46 ) ,
    .I1 ( config0_decoder3.n51 ) ) ;
or ( 
    .Z ( config0_decoder3.U7.AB ) ,
    .I0 ( config0_decoder3.n56 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U7.ZN ) ,
    .I0 ( config0_decoder3.U7.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_20 ) ,
    .IN ( config0_decoder3.U7.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U54.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n50 ) ) ;
and ( 
    .Z ( config0_decoder3.U54.ZN ) ,
    .I0 ( config0_decoder3.U54.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_13 ) ,
    .IN ( config0_decoder3.U54.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U42.AB ) ,
    .I0 ( config0_decoder3.n63 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U42.ZN ) ,
    .I0 ( config0_decoder3.U42.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_25 ) ,
    .IN ( config0_decoder3.U42.ZN ) ) ;
not ( 
    .O1 ( config0_decoder3.n39 ) ,
    .IN ( masks_hold_reg_2_9 ) ) ;
nand ( 
    .Z ( config0_decoder3.n54 ) ,
    .I0 ( config0_decoder3.n38 ) ,
    .I1 ( masks_hold_reg_2_7 ) ) ;
or ( 
    .Z ( config0_decoder3.U18.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n53 ) ) ;
and ( 
    .Z ( config0_decoder3.U18.ZN ) ,
    .I0 ( config0_decoder3.U18.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_0 ) ,
    .IN ( config0_decoder3.U18.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n55 ) ,
    .I0 ( config0_decoder3.n52 ) ,
    .I1 ( config0_decoder3.n51 ) ) ;
or ( 
    .Z ( config0_decoder3.U6.AB ) ,
    .I0 ( config0_decoder3.n59 ) ,
    .I1 ( config0_decoder3.n56 ) ) ;
and ( 
    .Z ( config0_decoder3.U6.ZN ) ,
    .I0 ( config0_decoder3.U6.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_4 ) ,
    .IN ( config0_decoder3.U6.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U85.AB ) ,
    .I0 ( config0_decoder3.n56 ) ,
    .I1 ( config0_decoder3.n55 ) ) ;
and ( 
    .Z ( config0_decoder3.U85.ZN ) ,
    .I0 ( config0_decoder3.U85.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_51 ) ,
    .IN ( config0_decoder3.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U45.AB ) ,
    .I0 ( config0_decoder3.n58 ) ,
    .I1 ( config0_decoder3.n43 ) ) ;
and ( 
    .Z ( config0_decoder3.U45.ZN ) ,
    .I0 ( config0_decoder3.U45.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_21 ) ,
    .IN ( config0_decoder3.U45.ZN ) ) ;
nor ( 
    .Z ( config0_decoder3.n46 ) ,
    .I0 ( config0_decoder3.n45 ) ,
    .I1 ( masks_hold_reg_2_10 ) ) ;
nand ( 
    .Z ( config0_decoder3.n57 ) ,
    .I0 ( n86 ) ,
    .I1 ( config0_decoder3.n52 ) ) ;
or ( 
    .Z ( config0_decoder3.U19.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n56 ) ) ;
and ( 
    .Z ( config0_decoder3.U19.ZN ) ,
    .I0 ( config0_decoder3.U19.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_3 ) ,
    .IN ( config0_decoder3.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U16.AB ) ,
    .I0 ( config0_decoder3.n62 ) ,
    .I1 ( config0_decoder3.n60 ) ) ;
and ( 
    .Z ( config0_decoder3.U16.ZN ) ,
    .I0 ( config0_decoder3.U16.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_7 ) ,
    .IN ( config0_decoder3.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U36.AB ) ,
    .I0 ( config0_decoder3.n54 ) ,
    .I1 ( config0_decoder3.n49 ) ) ;
and ( 
    .Z ( config0_decoder3.U36.ZN ) ,
    .I0 ( config0_decoder3.U36.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_34 ) ,
    .IN ( config0_decoder3.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U1.AB ) ,
    .I0 ( config0_decoder3.n47 ) ,
    .I1 ( config0_decoder3.n44 ) ) ;
and ( 
    .Z ( config0_decoder3.U1.ZN ) ,
    .I0 ( config0_decoder3.U1.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_28 ) ,
    .IN ( config0_decoder3.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder3.U84.AB ) ,
    .I0 ( config0_decoder3.n48 ) ,
    .I1 ( config0_decoder3.n47 ) ) ;
and ( 
    .Z ( config0_decoder3.U84.ZN ) ,
    .I0 ( config0_decoder3.U84.AB ) ,
    .I1 ( config0_decoder3.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_2_43 ) ,
    .IN ( config0_decoder3.U84.ZN ) ) ;
nand ( 
    .Z ( config0_decoder3.n56 ) ,
    .I0 ( config0_decoder3.n41 ) ,
    .I1 ( config0_decoder3.n39 ) ,
    .I2 ( masks_hold_reg_2_8 ) ) ;
or ( 
    .Z ( config0_decoder2.U54.AB ) ,
    .I0 ( config0_decoder2.n29 ) ,
    .I1 ( masks_hold_reg_1_8 ) ) ;
and ( 
    .Z ( config0_decoder2.U54.ZN ) ,
    .I0 ( config0_decoder2.U54.AB ) ,
    .I1 ( config0_decoder2.n17 ) ) ;
not ( 
    .O1 ( config0_decoder2.n1 ) ,
    .IN ( config0_decoder2.U54.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n22 ) ,
    .I0 ( masks_hold_reg_1_8 ) ,
    .I1 ( config0_decoder2.n28 ) ,
    .I2 ( masks_hold_reg_1_7 ) ) ;
or ( 
    .Z ( config0_decoder2.U44.AB ) ,
    .I0 ( config0_decoder2.n15 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U44.ZN ) ,
    .I0 ( config0_decoder2.U44.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_17 ) ,
    .IN ( config0_decoder2.U44.ZN ) ) ;
not ( 
    .O1 ( config0_decoder2.n30 ) ,
    .IN ( masks_hold_reg_1_8 ) ) ;
nand ( 
    .Z ( config0_decoder2.n25 ) ,
    .I0 ( config0_decoder2.n32 ) ,
    .I1 ( masks_hold_reg_1_5 ) ) ;
or ( 
    .Z ( config0_decoder2.U17.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n11 ) ) ;
and ( 
    .Z ( config0_decoder2.U17.ZN ) ,
    .I0 ( config0_decoder2.U17.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_6 ) ,
    .IN ( config0_decoder2.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U37.AB ) ,
    .I0 ( config0_decoder2.n9 ) ,
    .I1 ( config0_decoder2.n10 ) ) ;
and ( 
    .Z ( config0_decoder2.U37.ZN ) ,
    .I0 ( config0_decoder2.U37.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_8 ) ,
    .IN ( config0_decoder2.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U87.AB ) ,
    .I0 ( config0_decoder2.n12 ) ,
    .I1 ( config0_decoder2.n15 ) ) ;
and ( 
    .Z ( config0_decoder2.U87.ZN ) ,
    .I0 ( config0_decoder2.U87.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_50 ) ,
    .IN ( config0_decoder2.U87.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n10 ) ,
    .I0 ( masks_hold_reg_1_5 ) ,
    .I1 ( config0_decoder2.n34 ) ) ;
or ( 
    .Z ( config0_decoder2.U47.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n22 ) ) ;
and ( 
    .Z ( config0_decoder2.U47.ZN ) ,
    .I0 ( config0_decoder2.U47.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_11 ) ,
    .IN ( config0_decoder2.U47.ZN ) ) ;
not ( 
    .O1 ( config0_decoder2.n33 ) ,
    .IN ( masks_hold_reg_1_9 ) ) ;
nor ( 
    .Z ( config0_decoder2.n32 ) ,
    .I0 ( config0_decoder2.n33 ) ,
    .I1 ( masks_hold_reg_1_10 ) ) ;
nand ( 
    .Z ( config0_decoder2.n16 ) ,
    .I0 ( config0_decoder2.n31 ) ,
    .I1 ( config0_decoder2.n28 ) ) ;
or ( 
    .Z ( config0_decoder2.U34.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U34.ZN ) ,
    .I0 ( config0_decoder2.U34.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_26 ) ,
    .IN ( config0_decoder2.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U3.AB ) ,
    .I0 ( config0_decoder2.n16 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U3.ZN ) ,
    .I0 ( config0_decoder2.U3.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_31 ) ,
    .IN ( config0_decoder2.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U86.AB ) ,
    .I0 ( config0_decoder2.n12 ) ,
    .I1 ( config0_decoder2.n13 ) ) ;
and ( 
    .Z ( config0_decoder2.U86.ZN ) ,
    .I0 ( config0_decoder2.U86.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_52 ) ,
    .IN ( config0_decoder2.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n15 ) ,
    .I0 ( config0_decoder2.n31 ) ,
    .I1 ( masks_hold_reg_1_6 ) ) ;
or ( 
    .Z ( config0_decoder2.U46.AB ) ,
    .I0 ( config0_decoder2.n11 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U46.ZN ) ,
    .I0 ( config0_decoder2.U46.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_21 ) ,
    .IN ( config0_decoder2.U46.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U74.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n15 ) ) ;
and ( 
    .Z ( config0_decoder2.U74.ZN ) ,
    .I0 ( config0_decoder2.U74.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_1 ) ,
    .IN ( config0_decoder2.U74.ZN ) ) ;
not ( 
    .O1 ( config0_decoder2.n18 ) ,
    .IN ( masks_hold_reg_1_5 ) ) ;
nand ( 
    .Z ( config0_decoder2.n9 ) ,
    .I0 ( config0_decoder2.n27 ) ,
    .I1 ( config0_decoder2.n28 ) ) ;
or ( 
    .Z ( config0_decoder2.U38.AB ) ,
    .I0 ( config0_decoder2.n11 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U38.ZN ) ,
    .I0 ( config0_decoder2.U38.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_22 ) ,
    .IN ( config0_decoder2.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U35.AB ) ,
    .I0 ( config0_decoder2.n15 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U35.ZN ) ,
    .I0 ( config0_decoder2.U35.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_34 ) ,
    .IN ( config0_decoder2.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U2.AB ) ,
    .I0 ( config0_decoder2.n19 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U2.ZN ) ,
    .I0 ( config0_decoder2.U2.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_30 ) ,
    .IN ( config0_decoder2.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U81.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n11 ) ) ;
and ( 
    .Z ( config0_decoder2.U81.ZN ) ,
    .I0 ( config0_decoder2.U81.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_5 ) ,
    .IN ( config0_decoder2.U81.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n20 ) ,
    .I0 ( config0_decoder2.n23 ) ,
    .I1 ( masks_hold_reg_1_5 ) ) ;
or ( 
    .Z ( config0_decoder2.U49.AB ) ,
    .I0 ( config0_decoder2.n13 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U49.ZN ) ,
    .I0 ( config0_decoder2.U49.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_35 ) ,
    .IN ( config0_decoder2.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U75.AB ) ,
    .I0 ( config0_decoder2.n13 ) ,
    .I1 ( config0_decoder2.n14 ) ) ;
and ( 
    .Z ( config0_decoder2.U75.ZN ) ,
    .I0 ( config0_decoder2.U75.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_51 ) ,
    .IN ( config0_decoder2.U75.ZN ) ) ;
nor ( 
    .Z ( config0_decoder2.n31 ) ,
    .I0 ( masks_hold_reg_1_7 ) ,
    .I1 ( masks_hold_reg_1_8 ) ) ;
nand ( 
    .Z ( config0_decoder2.n11 ) ,
    .I0 ( config0_decoder2.n29 ) ,
    .I1 ( config0_decoder2.n30 ) ) ;
or ( 
    .Z ( config0_decoder2.U39.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n22 ) ) ;
and ( 
    .Z ( config0_decoder2.U39.ZN ) ,
    .I0 ( config0_decoder2.U39.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_12 ) ,
    .IN ( config0_decoder2.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U32.AB ) ,
    .I0 ( config0_decoder2.n13 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U32.ZN ) ,
    .I0 ( config0_decoder2.U32.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_20 ) ,
    .IN ( config0_decoder2.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U29.AB ) ,
    .I0 ( config0_decoder2.n9 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U29.ZN ) ,
    .I0 ( config0_decoder2.U29.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_24 ) ,
    .IN ( config0_decoder2.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U80.AB ) ,
    .I0 ( config0_decoder2.n19 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U80.ZN ) ,
    .I0 ( config0_decoder2.U80.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_45 ) ,
    .IN ( config0_decoder2.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U48.AB ) ,
    .I0 ( config0_decoder2.n22 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U48.ZN ) ,
    .I0 ( config0_decoder2.U48.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_27 ) ,
    .IN ( config0_decoder2.U48.ZN ) ) ;
nor ( 
    .Z ( config0_decoder2.n34 ) ,
    .I0 ( masks_hold_reg_1_9 ) ,
    .I1 ( masks_hold_reg_1_10 ) ) ;
nor ( 
    .Z ( config0_decoder2.n17 ) ,
    .I0 ( config0_decoder2.n24 ) ,
    .I1 ( config0_decoder2.n33 ) ) ;
or ( 
    .Z ( config0_decoder2.U33.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n10 ) ) ;
and ( 
    .Z ( config0_decoder2.U33.ZN ) ,
    .I0 ( config0_decoder2.U33.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_10 ) ,
    .IN ( config0_decoder2.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U28.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n19 ) ) ;
and ( 
    .Z ( config0_decoder2.U28.ZN ) ,
    .I0 ( config0_decoder2.U28.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_14 ) ,
    .IN ( config0_decoder2.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U83.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U83.ZN ) ,
    .I0 ( config0_decoder2.U83.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_42 ) ,
    .IN ( config0_decoder2.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U50.AB ) ,
    .I0 ( config0_decoder2.n9 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U50.ZN ) ,
    .I0 ( config0_decoder2.U50.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_39 ) ,
    .IN ( config0_decoder2.U50.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U30.AB ) ,
    .I0 ( config0_decoder2.n16 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U30.ZN ) ,
    .I0 ( config0_decoder2.U30.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_32 ) ,
    .IN ( config0_decoder2.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U22.AB ) ,
    .I0 ( config0_decoder2.n14 ) ,
    .I1 ( config0_decoder2.n15 ) ) ;
and ( 
    .Z ( config0_decoder2.U22.ZN ) ,
    .I0 ( config0_decoder2.U22.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_49 ) ,
    .IN ( config0_decoder2.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U82.AB ) ,
    .I0 ( config0_decoder2.n9 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U82.ZN ) ,
    .I0 ( config0_decoder2.U82.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_40 ) ,
    .IN ( config0_decoder2.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U51.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n7 ) ) ;
and ( 
    .Z ( config0_decoder2.U51.ZN ) ,
    .I0 ( config0_decoder2.U51.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_9 ) ,
    .IN ( config0_decoder2.U51.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U41.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U41.ZN ) ,
    .I0 ( config0_decoder2.U41.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_25 ) ,
    .IN ( config0_decoder2.U41.ZN ) ) ;
not ( 
    .O1 ( config0_decoder2.n24 ) ,
    .IN ( masks_hold_reg_1_10 ) ) ;
or ( 
    .Z ( config0_decoder2.U31.AB ) ,
    .I0 ( config0_decoder2.n13 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U31.ZN ) ,
    .I0 ( config0_decoder2.U31.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_36 ) ,
    .IN ( config0_decoder2.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U21.AB ) ,
    .I0 ( config0_decoder2.n12 ) ,
    .I1 ( config0_decoder2.n16 ) ) ;
and ( 
    .Z ( config0_decoder2.U21.ZN ) ,
    .I0 ( config0_decoder2.U21.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_48 ) ,
    .IN ( config0_decoder2.U21.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U5.AB ) ,
    .I0 ( config0_decoder2.n15 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U5.ZN ) ,
    .I0 ( config0_decoder2.U5.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_18 ) ,
    .IN ( config0_decoder2.U5.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U52.AB ) ,
    .I0 ( config0_decoder2.n9 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U52.ZN ) ,
    .I0 ( config0_decoder2.U52.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_23 ) ,
    .IN ( config0_decoder2.U52.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U40.AB ) ,
    .I0 ( config0_decoder2.n19 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U40.ZN ) ,
    .I0 ( config0_decoder2.U40.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_29 ) ,
    .IN ( config0_decoder2.U40.ZN ) ) ;
and ( 
    .Z ( config0_decoder2.n29 ) ,
    .I0 ( masks_hold_reg_1_7 ) ,
    .I1 ( masks_hold_reg_1_6 ) ) ;
or ( 
    .Z ( config0_decoder2.U72.AB ) ,
    .I0 ( config0_decoder2.n14 ) ,
    .I1 ( config0_decoder2.n16 ) ) ;
and ( 
    .Z ( config0_decoder2.U72.ZN ) ,
    .I0 ( config0_decoder2.U72.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_47 ) ,
    .IN ( config0_decoder2.U72.ZN ) ) ;
nor ( 
    .Z ( config0_decoder2.n23 ) ,
    .I0 ( config0_decoder2.n24 ) ,
    .I1 ( masks_hold_reg_1_9 ) ) ;
or ( 
    .Z ( config0_decoder2.U20.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n15 ) ) ;
and ( 
    .Z ( config0_decoder2.U20.ZN ) ,
    .I0 ( config0_decoder2.U20.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_2 ) ,
    .IN ( config0_decoder2.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n26 ) ,
    .I0 ( config0_decoder2.n32 ) ,
    .I1 ( config0_decoder2.n18 ) ) ;
or ( 
    .Z ( config0_decoder2.U4.AB ) ,
    .I0 ( config0_decoder2.n16 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U4.ZN ) ,
    .I0 ( config0_decoder2.U4.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_16 ) ,
    .IN ( config0_decoder2.U4.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U53.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n19 ) ) ;
and ( 
    .Z ( config0_decoder2.U53.ZN ) ,
    .I0 ( config0_decoder2.U53.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_13 ) ,
    .IN ( config0_decoder2.U53.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U43.AB ) ,
    .I0 ( config0_decoder2.n11 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U43.ZN ) ,
    .I0 ( config0_decoder2.U43.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_37 ) ,
    .IN ( config0_decoder2.U43.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U73.AB ) ,
    .I0 ( config0_decoder2.n19 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U73.ZN ) ,
    .I0 ( config0_decoder2.U73.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_46 ) ,
    .IN ( config0_decoder2.U73.ZN ) ) ;
nor ( 
    .Z ( config0_decoder2.n27 ) ,
    .I0 ( config0_decoder2.n30 ) ,
    .I1 ( masks_hold_reg_1_7 ) ) ;
nand ( 
    .Z ( config0_decoder2.n12 ) ,
    .I0 ( masks_hold_reg_1_5 ) ,
    .I1 ( config0_decoder2.n17 ) ) ;
nand ( 
    .Z ( config0_decoder2.n14 ) ,
    .I0 ( config0_decoder2.n17 ) ,
    .I1 ( config0_decoder2.n18 ) ) ;
nand ( 
    .Z ( config0_decoder2.n7 ) ,
    .I0 ( config0_decoder2.n34 ) ,
    .I1 ( config0_decoder2.n18 ) ) ;
nand ( 
    .Z ( config0_decoder2.n21 ) ,
    .I0 ( config0_decoder2.n23 ) ,
    .I1 ( config0_decoder2.n18 ) ) ;
or ( 
    .Z ( config0_decoder2.U42.AB ) ,
    .I0 ( config0_decoder2.n15 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U42.ZN ) ,
    .I0 ( config0_decoder2.U42.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_33 ) ,
    .IN ( config0_decoder2.U42.ZN ) ) ;
not ( 
    .O1 ( config0_decoder2.n28 ) ,
    .IN ( masks_hold_reg_1_6 ) ) ;
nand ( 
    .Z ( config0_decoder2.n19 ) ,
    .I0 ( config0_decoder2.n29 ) ,
    .I1 ( masks_hold_reg_1_8 ) ) ;
or ( 
    .Z ( config0_decoder2.U18.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n16 ) ) ;
and ( 
    .Z ( config0_decoder2.U18.ZN ) ,
    .I0 ( config0_decoder2.U18.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_0 ) ,
    .IN ( config0_decoder2.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U15.AB ) ,
    .I0 ( config0_decoder2.n10 ) ,
    .I1 ( config0_decoder2.n13 ) ) ;
and ( 
    .Z ( config0_decoder2.U15.ZN ) ,
    .I0 ( config0_decoder2.U15.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_4 ) ,
    .IN ( config0_decoder2.U15.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U6.AB ) ,
    .I0 ( config0_decoder2.n13 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U6.ZN ) ,
    .I0 ( config0_decoder2.U6.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_19 ) ,
    .IN ( config0_decoder2.U6.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U85.AB ) ,
    .I0 ( config0_decoder2.n21 ) ,
    .I1 ( config0_decoder2.n22 ) ) ;
and ( 
    .Z ( config0_decoder2.U85.ZN ) ,
    .I0 ( config0_decoder2.U85.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_43 ) ,
    .IN ( config0_decoder2.U85.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n13 ) ,
    .I0 ( config0_decoder2.n28 ) ,
    .I1 ( config0_decoder2.n30 ) ,
    .I2 ( masks_hold_reg_1_7 ) ) ;
or ( 
    .Z ( config0_decoder2.U45.AB ) ,
    .I0 ( config0_decoder2.n16 ) ,
    .I1 ( config0_decoder2.n26 ) ) ;
and ( 
    .Z ( config0_decoder2.U45.ZN ) ,
    .I0 ( config0_decoder2.U45.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_15 ) ,
    .IN ( config0_decoder2.U45.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U71.AB ) ,
    .I0 ( config0_decoder2.n20 ) ,
    .I1 ( config0_decoder2.n22 ) ) ;
and ( 
    .Z ( config0_decoder2.U71.ZN ) ,
    .I0 ( config0_decoder2.U71.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_44 ) ,
    .IN ( config0_decoder2.U71.ZN ) ) ;
nand ( 
    .Z ( config0_decoder2.n6 ) ,
    .I0 ( masks_hold_reg_1_6 ) ,
    .I1 ( config0_decoder2.n27 ) ) ;
or ( 
    .Z ( config0_decoder2.U19.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n13 ) ) ;
and ( 
    .Z ( config0_decoder2.U19.ZN ) ,
    .I0 ( config0_decoder2.U19.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_3 ) ,
    .IN ( config0_decoder2.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U16.AB ) ,
    .I0 ( config0_decoder2.n7 ) ,
    .I1 ( config0_decoder2.n9 ) ) ;
and ( 
    .Z ( config0_decoder2.U16.ZN ) ,
    .I0 ( config0_decoder2.U16.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_7 ) ,
    .IN ( config0_decoder2.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U36.AB ) ,
    .I0 ( config0_decoder2.n11 ) ,
    .I1 ( config0_decoder2.n20 ) ) ;
and ( 
    .Z ( config0_decoder2.U36.ZN ) ,
    .I0 ( config0_decoder2.U36.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_38 ) ,
    .IN ( config0_decoder2.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U1.AB ) ,
    .I0 ( config0_decoder2.n22 ) ,
    .I1 ( config0_decoder2.n25 ) ) ;
and ( 
    .Z ( config0_decoder2.U1.ZN ) ,
    .I0 ( config0_decoder2.U1.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_28 ) ,
    .IN ( config0_decoder2.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder2.U84.AB ) ,
    .I0 ( config0_decoder2.n6 ) ,
    .I1 ( config0_decoder2.n21 ) ) ;
and ( 
    .Z ( config0_decoder2.U84.ZN ) ,
    .I0 ( config0_decoder2.U84.AB ) ,
    .I1 ( config0_decoder2.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_1_41 ) ,
    .IN ( config0_decoder2.U84.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n1 ) ,
    .I0 ( config0_decoder1.n16 ) ,
    .I1 ( config0_decoder1.n40 ) ) ;
nand ( 
    .Z ( config0_decoder1.n14 ) ,
    .I0 ( config0_decoder1.n15 ) ,
    .I1 ( config0_decoder1.n16 ) ) ;
or ( 
    .Z ( config0_decoder1.U84.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n34 ) ) ;
and ( 
    .Z ( config0_decoder1.U84.ZN ) ,
    .I0 ( config0_decoder1.U84.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_17 ) ,
    .IN ( config0_decoder1.U84.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n10 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( config0_decoder1.n39 ) ) ;
or ( 
    .Z ( config0_decoder1.U44.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n29 ) ) ;
and ( 
    .Z ( config0_decoder1.U44.ZN ) ,
    .I0 ( config0_decoder1.U44.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_2 ) ,
    .IN ( config0_decoder1.U44.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U76.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n28 ) ) ;
and ( 
    .Z ( config0_decoder1.U76.ZN ) ,
    .I0 ( config0_decoder1.U76.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_27 ) ,
    .IN ( config0_decoder1.U76.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n39 ) ,
    .IN ( masks_hold_reg_0_5 ) ) ;
or ( 
    .Z ( config0_decoder1.U17.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n26 ) ) ;
and ( 
    .Z ( config0_decoder1.U17.ZN ) ,
    .I0 ( config0_decoder1.U17.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_33 ) ,
    .IN ( config0_decoder1.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U37.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n17 ) ) ;
and ( 
    .Z ( config0_decoder1.U37.ZN ) ,
    .I0 ( config0_decoder1.U37.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_49 ) ,
    .IN ( config0_decoder1.U37.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n26 ) ,
    .I0 ( config0_decoder1.n20 ) ,
    .I1 ( config0_decoder1.n18 ) ) ;
or ( 
    .Z ( config0_decoder1.U87.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n17 ) ) ;
and ( 
    .Z ( config0_decoder1.U87.ZN ) ,
    .I0 ( config0_decoder1.U87.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_50 ) ,
    .IN ( config0_decoder1.U87.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n37 ) ,
    .IN ( masks_hold_reg_0_4 ) ) ;
or ( 
    .Z ( config0_decoder1.U47.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n36 ) ) ;
and ( 
    .Z ( config0_decoder1.U47.ZN ) ,
    .I0 ( config0_decoder1.U47.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_14 ) ,
    .IN ( config0_decoder1.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U77.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n31 ) ) ;
and ( 
    .Z ( config0_decoder1.U77.ZN ) ,
    .I0 ( config0_decoder1.U77.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_24 ) ,
    .IN ( config0_decoder1.U77.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n38 ) ,
    .IN ( masks_hold_reg_0_7 ) ) ;
or ( 
    .Z ( config0_decoder1.U10.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n19 ) ) ;
and ( 
    .Z ( config0_decoder1.U10.ZN ) ,
    .I0 ( config0_decoder1.U10.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_43 ) ,
    .IN ( config0_decoder1.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n31 ) ,
    .I0 ( config0_decoder1.n30 ) ,
    .I1 ( config0_decoder1.n24 ) ) ;
nand ( 
    .Z ( config0_decoder1.n25 ) ,
    .I0 ( config0_decoder1.n20 ) ,
    .I1 ( config0_decoder1.n15 ) ) ;
or ( 
    .Z ( config0_decoder1.U90.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n36 ) ) ;
and ( 
    .Z ( config0_decoder1.U90.ZN ) ,
    .I0 ( config0_decoder1.U90.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_11 ) ,
    .IN ( config0_decoder1.U90.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U86.AB ) ,
    .I0 ( config0_decoder1.n7 ) ,
    .I1 ( config0_decoder1.n8 ) ) ;
and ( 
    .Z ( config0_decoder1.U86.ZN ) ,
    .I0 ( config0_decoder1.U86.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_9 ) ,
    .IN ( config0_decoder1.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n8 ) ,
    .I0 ( masks_hold_reg_0_5 ) ,
    .I1 ( config0_decoder1.n37 ) ) ;
or ( 
    .Z ( config0_decoder1.U46.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n34 ) ) ;
and ( 
    .Z ( config0_decoder1.U46.ZN ) ,
    .I0 ( config0_decoder1.U46.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_15 ) ,
    .IN ( config0_decoder1.U46.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U74.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n26 ) ) ;
and ( 
    .Z ( config0_decoder1.U74.ZN ) ,
    .I0 ( config0_decoder1.U74.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_31 ) ,
    .IN ( config0_decoder1.U74.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n35 ) ,
    .IN ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config0_decoder1.U11.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n19 ) ) ;
and ( 
    .Z ( config0_decoder1.U11.ZN ) ,
    .I0 ( config0_decoder1.U11.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_44 ) ,
    .IN ( config0_decoder1.U11.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U38.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n17 ) ) ;
and ( 
    .Z ( config0_decoder1.U38.ZN ) ,
    .I0 ( config0_decoder1.U38.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_48 ) ,
    .IN ( config0_decoder1.U38.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n29 ) ,
    .I0 ( config0_decoder1.n18 ) ,
    .I1 ( config0_decoder1.n23 ) ) ;
nand ( 
    .Z ( config0_decoder1.n22 ) ,
    .I0 ( config0_decoder1.n20 ) ,
    .I1 ( config0_decoder1.n24 ) ) ;
or ( 
    .Z ( config0_decoder1.U91.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n29 ) ) ;
and ( 
    .Z ( config0_decoder1.U91.ZN ) ,
    .I0 ( config0_decoder1.U91.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_1 ) ,
    .IN ( config0_decoder1.U91.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U81.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n31 ) ) ;
and ( 
    .Z ( config0_decoder1.U81.ZN ) ,
    .I0 ( config0_decoder1.U81.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_26 ) ,
    .IN ( config0_decoder1.U81.ZN ) ) ;
nor ( 
    .Z ( config0_decoder1.n23 ) ,
    .I0 ( masks_hold_reg_0_8 ) ,
    .I1 ( masks_hold_reg_0_9 ) ) ;
or ( 
    .Z ( config0_decoder1.U49.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n13 ) ) ;
and ( 
    .Z ( config0_decoder1.U49.ZN ) ,
    .I0 ( config0_decoder1.U49.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_4 ) ,
    .IN ( config0_decoder1.U49.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U75.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n28 ) ) ;
and ( 
    .Z ( config0_decoder1.U75.ZN ) ,
    .I0 ( config0_decoder1.U75.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_29 ) ,
    .IN ( config0_decoder1.U75.ZN ) ) ;
nor ( 
    .Z ( config0_decoder1.n24 ) ,
    .I0 ( config0_decoder1.n38 ) ,
    .I1 ( masks_hold_reg_0_6 ) ) ;
or ( 
    .Z ( config0_decoder1.U12.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n19 ) ) ;
and ( 
    .Z ( config0_decoder1.U12.ZN ) ,
    .I0 ( config0_decoder1.U12.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_46 ) ,
    .IN ( config0_decoder1.U12.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U39.AB ) ,
    .I0 ( config0_decoder1.n7 ) ,
    .I1 ( config0_decoder1.n12 ) ) ;
and ( 
    .Z ( config0_decoder1.U39.ZN ) ,
    .I0 ( config0_decoder1.U39.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_10 ) ,
    .IN ( config0_decoder1.U39.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n34 ) ,
    .I0 ( config0_decoder1.n30 ) ,
    .I1 ( config0_decoder1.n18 ) ) ;
nand ( 
    .Z ( config0_decoder1.n13 ) ,
    .I0 ( config0_decoder1.n15 ) ,
    .I1 ( config0_decoder1.n23 ) ) ;
nand ( 
    .Z ( config0_decoder1.n19 ) ,
    .I0 ( config0_decoder1.n20 ) ,
    .I1 ( config0_decoder1.n21 ) ) ;
or ( 
    .Z ( config0_decoder1.U92.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n14 ) ) ;
and ( 
    .Z ( config0_decoder1.U92.ZN ) ,
    .I0 ( config0_decoder1.U92.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_53 ) ,
    .IN ( config0_decoder1.U92.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U80.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n28 ) ) ;
and ( 
    .Z ( config0_decoder1.U80.ZN ) ,
    .I0 ( config0_decoder1.U80.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_30 ) ,
    .IN ( config0_decoder1.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U48.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n13 ) ) ;
and ( 
    .Z ( config0_decoder1.U48.ZN ) ,
    .I0 ( config0_decoder1.U48.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_5 ) ,
    .IN ( config0_decoder1.U48.ZN ) ) ;
nor ( 
    .Z ( config0_decoder1.n30 ) ,
    .I0 ( config0_decoder1.n35 ) ,
    .I1 ( masks_hold_reg_0_9 ) ) ;
or ( 
    .Z ( config0_decoder1.U13.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n17 ) ) ;
and ( 
    .Z ( config0_decoder1.U13.ZN ) ,
    .I0 ( config0_decoder1.U13.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_47 ) ,
    .IN ( config0_decoder1.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n28 ) ,
    .I0 ( config0_decoder1.n30 ) ,
    .I1 ( config0_decoder1.n21 ) ) ;
nand ( 
    .Z ( config0_decoder1.n17 ) ,
    .I0 ( config0_decoder1.n18 ) ,
    .I1 ( config0_decoder1.n16 ) ) ;
nor ( 
    .Z ( config0_decoder1.n16 ) ,
    .I0 ( config0_decoder1.n27 ) ,
    .I1 ( config0_decoder1.n35 ) ) ;
or ( 
    .Z ( config0_decoder1.U93.AB ) ,
    .I0 ( config0_decoder1.n7 ) ,
    .I1 ( config0_decoder1.n11 ) ) ;
and ( 
    .Z ( config0_decoder1.U93.ZN ) ,
    .I0 ( config0_decoder1.U93.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_7 ) ,
    .IN ( config0_decoder1.U93.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U83.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n28 ) ) ;
and ( 
    .Z ( config0_decoder1.U83.ZN ) ,
    .I0 ( config0_decoder1.U83.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_28 ) ,
    .IN ( config0_decoder1.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U50.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n13 ) ) ;
and ( 
    .Z ( config0_decoder1.U50.ZN ) ,
    .I0 ( config0_decoder1.U50.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_6 ) ,
    .IN ( config0_decoder1.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n36 ) ,
    .I0 ( config0_decoder1.n21 ) ,
    .I1 ( config0_decoder1.n23 ) ) ;
nor ( 
    .Z ( config0_decoder1.n21 ) ,
    .I0 ( config0_decoder1.n33 ) ,
    .I1 ( config0_decoder1.n38 ) ) ;
or ( 
    .Z ( config0_decoder1.U82.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n32 ) ) ;
and ( 
    .Z ( config0_decoder1.U82.ZN ) ,
    .I0 ( config0_decoder1.U82.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_20 ) ,
    .IN ( config0_decoder1.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U89.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n14 ) ) ;
and ( 
    .Z ( config0_decoder1.U89.ZN ) ,
    .I0 ( config0_decoder1.U89.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_51 ) ,
    .IN ( config0_decoder1.U89.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n12 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( masks_hold_reg_0_5 ) ) ;
or ( 
    .Z ( config0_decoder1.U41.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n36 ) ) ;
and ( 
    .Z ( config0_decoder1.U41.ZN ) ,
    .I0 ( config0_decoder1.U41.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_13 ) ,
    .IN ( config0_decoder1.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U78.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n32 ) ) ;
and ( 
    .Z ( config0_decoder1.U78.ZN ) ,
    .I0 ( config0_decoder1.U78.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_22 ) ,
    .IN ( config0_decoder1.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder1.n32 ) ,
    .I0 ( config0_decoder1.n30 ) ,
    .I1 ( config0_decoder1.n15 ) ) ;
nand ( 
    .Z ( config0_decoder1.n7 ) ,
    .I0 ( config0_decoder1.n23 ) ,
    .I1 ( config0_decoder1.n24 ) ) ;
or ( 
    .Z ( config0_decoder1.U88.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n14 ) ) ;
and ( 
    .Z ( config0_decoder1.U88.ZN ) ,
    .I0 ( config0_decoder1.U88.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_52 ) ,
    .IN ( config0_decoder1.U88.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U52.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n22 ) ) ;
and ( 
    .Z ( config0_decoder1.U52.ZN ) ,
    .I0 ( config0_decoder1.U52.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_41 ) ,
    .IN ( config0_decoder1.U52.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U40.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n36 ) ) ;
and ( 
    .Z ( config0_decoder1.U40.ZN ) ,
    .I0 ( config0_decoder1.U40.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_12 ) ,
    .IN ( config0_decoder1.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U79.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n34 ) ) ;
and ( 
    .Z ( config0_decoder1.U79.ZN ) ,
    .I0 ( config0_decoder1.U79.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_18 ) ,
    .IN ( config0_decoder1.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U72.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n32 ) ) ;
and ( 
    .Z ( config0_decoder1.U72.ZN ) ,
    .I0 ( config0_decoder1.U72.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_19 ) ,
    .IN ( config0_decoder1.U72.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n27 ) ,
    .IN ( masks_hold_reg_0_9 ) ) ;
nand ( 
    .Z ( config0_decoder1.n11 ) ,
    .I0 ( config0_decoder1.n37 ) ,
    .I1 ( config0_decoder1.n39 ) ) ;
or ( 
    .Z ( config0_decoder1.U9.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n22 ) ) ;
and ( 
    .Z ( config0_decoder1.U9.ZN ) ,
    .I0 ( config0_decoder1.U9.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_42 ) ,
    .IN ( config0_decoder1.U9.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U53.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n19 ) ) ;
and ( 
    .Z ( config0_decoder1.U53.ZN ) ,
    .I0 ( config0_decoder1.U53.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_45 ) ,
    .IN ( config0_decoder1.U53.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U43.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n29 ) ) ;
and ( 
    .Z ( config0_decoder1.U43.ZN ) ,
    .I0 ( config0_decoder1.U43.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_0 ) ,
    .IN ( config0_decoder1.U43.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U73.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n34 ) ) ;
and ( 
    .Z ( config0_decoder1.U73.ZN ) ,
    .I0 ( config0_decoder1.U73.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_16 ) ,
    .IN ( config0_decoder1.U73.ZN ) ) ;
not ( 
    .O1 ( config0_decoder1.n33 ) ,
    .IN ( masks_hold_reg_0_6 ) ) ;
nor ( 
    .Z ( config0_decoder1.n15 ) ,
    .I0 ( config0_decoder1.n33 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
or ( 
    .Z ( config0_decoder1.U14.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n22 ) ) ;
and ( 
    .Z ( config0_decoder1.U14.ZN ) ,
    .I0 ( config0_decoder1.U14.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_39 ) ,
    .IN ( config0_decoder1.U14.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U8.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n22 ) ) ;
and ( 
    .Z ( config0_decoder1.U8.ZN ) ,
    .I0 ( config0_decoder1.U8.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_40 ) ,
    .IN ( config0_decoder1.U8.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U7.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n33 ) ) ;
and ( 
    .Z ( config0_decoder1.U7.ZN ) ,
    .I0 ( config0_decoder1.U7.AB ) ,
    .I1 ( config0_decoder1.n38 ) ) ;
not ( 
    .O1 ( config0_decoder1.n40 ) ,
    .IN ( config0_decoder1.U7.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U54.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n25 ) ) ;
and ( 
    .Z ( config0_decoder1.U54.ZN ) ,
    .I0 ( config0_decoder1.U54.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_37 ) ,
    .IN ( config0_decoder1.U54.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U42.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n13 ) ) ;
and ( 
    .Z ( config0_decoder1.U42.ZN ) ,
    .I0 ( config0_decoder1.U42.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_3 ) ,
    .IN ( config0_decoder1.U42.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U70.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n31 ) ) ;
and ( 
    .Z ( config0_decoder1.U70.ZN ) ,
    .I0 ( config0_decoder1.U70.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_23 ) ,
    .IN ( config0_decoder1.U70.ZN ) ) ;
nor ( 
    .Z ( config0_decoder1.n18 ) ,
    .I0 ( masks_hold_reg_0_6 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
or ( 
    .Z ( config0_decoder1.U18.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n26 ) ) ;
and ( 
    .Z ( config0_decoder1.U18.ZN ) ,
    .I0 ( config0_decoder1.U18.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_32 ) ,
    .IN ( config0_decoder1.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U15.AB ) ,
    .I0 ( config0_decoder1.n10 ) ,
    .I1 ( config0_decoder1.n25 ) ) ;
and ( 
    .Z ( config0_decoder1.U15.ZN ) ,
    .I0 ( config0_decoder1.U15.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_36 ) ,
    .IN ( config0_decoder1.U15.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U85.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n31 ) ) ;
and ( 
    .Z ( config0_decoder1.U85.ZN ) ,
    .I0 ( config0_decoder1.U85.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_25 ) ,
    .IN ( config0_decoder1.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U55.AB ) ,
    .I0 ( config0_decoder1.n11 ) ,
    .I1 ( config0_decoder1.n25 ) ) ;
and ( 
    .Z ( config0_decoder1.U55.ZN ) ,
    .I0 ( config0_decoder1.U55.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_35 ) ,
    .IN ( config0_decoder1.U55.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U45.AB ) ,
    .I0 ( config0_decoder1.n7 ) ,
    .I1 ( config0_decoder1.n10 ) ) ;
and ( 
    .Z ( config0_decoder1.U45.ZN ) ,
    .I0 ( config0_decoder1.U45.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_8 ) ,
    .IN ( config0_decoder1.U45.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U71.AB ) ,
    .I0 ( config0_decoder1.n8 ) ,
    .I1 ( config0_decoder1.n32 ) ) ;
and ( 
    .Z ( config0_decoder1.U71.ZN ) ,
    .I0 ( config0_decoder1.U71.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_21 ) ,
    .IN ( config0_decoder1.U71.ZN ) ) ;
nor ( 
    .Z ( config0_decoder1.n20 ) ,
    .I0 ( config0_decoder1.n27 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config0_decoder1.U19.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n26 ) ) ;
and ( 
    .Z ( config0_decoder1.U19.ZN ) ,
    .I0 ( config0_decoder1.U19.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_34 ) ,
    .IN ( config0_decoder1.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder1.U16.AB ) ,
    .I0 ( config0_decoder1.n12 ) ,
    .I1 ( config0_decoder1.n25 ) ) ;
and ( 
    .Z ( config0_decoder1.U16.ZN ) ,
    .I0 ( config0_decoder1.U16.AB ) ,
    .I1 ( config0_decoder1.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_0_38 ) ,
    .IN ( config0_decoder1.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U54.AB ) ,
    .I0 ( config0_decoder7.n40 ) ,
    .I1 ( masks_hold_reg_5_2 ) ) ;
and ( 
    .Z ( config0_decoder7.U54.ZN ) ,
    .I0 ( config0_decoder7.U54.AB ) ,
    .I1 ( config0_decoder7.n52 ) ) ;
not ( 
    .O1 ( config0_decoder7.n1 ) ,
    .IN ( config0_decoder7.U54.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n59 ) ,
    .I0 ( masks_hold_reg_6_10 ) ,
    .I1 ( config0_decoder7.n35 ) ) ;
or ( 
    .Z ( config0_decoder7.U44.AB ) ,
    .I0 ( config0_decoder7.n58 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U44.ZN ) ,
    .I0 ( config0_decoder7.U44.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_21 ) ,
    .IN ( config0_decoder7.U44.ZN ) ) ;
not ( 
    .O1 ( config0_decoder7.n45 ) ,
    .IN ( masks_hold_reg_5_4 ) ) ;
nand ( 
    .Z ( config0_decoder7.n54 ) ,
    .I0 ( config0_decoder7.n38 ) ,
    .I1 ( masks_hold_reg_5_0 ) ) ;
or ( 
    .Z ( config0_decoder7.U17.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n53 ) ) ;
and ( 
    .Z ( config0_decoder7.U17.ZN ) ,
    .I0 ( config0_decoder7.U17.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_0 ) ,
    .IN ( config0_decoder7.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U37.AB ) ,
    .I0 ( config0_decoder7.n60 ) ,
    .I1 ( config0_decoder7.n59 ) ) ;
and ( 
    .Z ( config0_decoder7.U37.ZN ) ,
    .I0 ( config0_decoder7.U37.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_8 ) ,
    .IN ( config0_decoder7.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U87.AB ) ,
    .I0 ( config0_decoder7.n57 ) ,
    .I1 ( config0_decoder7.n54 ) ) ;
and ( 
    .Z ( config0_decoder7.U87.ZN ) ,
    .I0 ( config0_decoder7.U87.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_50 ) ,
    .IN ( config0_decoder7.U87.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n47 ) ,
    .I0 ( masks_hold_reg_5_2 ) ,
    .I1 ( config0_decoder7.n41 ) ,
    .I2 ( masks_hold_reg_5_1 ) ) ;
or ( 
    .Z ( config0_decoder7.U47.AB ) ,
    .I0 ( config0_decoder7.n54 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U47.ZN ) ,
    .I0 ( config0_decoder7.U47.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_17 ) ,
    .IN ( config0_decoder7.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U77.AB ) ,
    .I0 ( config0_decoder7.n50 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U77.ZN ) ,
    .I0 ( config0_decoder7.U77.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_46 ) ,
    .IN ( config0_decoder7.U77.ZN ) ) ;
nor ( 
    .Z ( config0_decoder7.n42 ) ,
    .I0 ( config0_decoder7.n39 ) ,
    .I1 ( masks_hold_reg_5_1 ) ) ;
nand ( 
    .Z ( config0_decoder7.n60 ) ,
    .I0 ( config0_decoder7.n42 ) ,
    .I1 ( config0_decoder7.n41 ) ) ;
or ( 
    .Z ( config0_decoder7.U34.AB ) ,
    .I0 ( config0_decoder7.n54 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U34.ZN ) ,
    .I0 ( config0_decoder7.U34.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_34 ) ,
    .IN ( config0_decoder7.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U3.AB ) ,
    .I0 ( config0_decoder7.n50 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U3.ZN ) ,
    .I0 ( config0_decoder7.U3.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_30 ) ,
    .IN ( config0_decoder7.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U86.AB ) ,
    .I0 ( config0_decoder7.n57 ) ,
    .I1 ( config0_decoder7.n56 ) ) ;
and ( 
    .Z ( config0_decoder7.U86.ZN ) ,
    .I0 ( config0_decoder7.U86.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_52 ) ,
    .IN ( config0_decoder7.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n49 ) ,
    .I0 ( config0_decoder7.n46 ) ,
    .I1 ( masks_hold_reg_6_10 ) ) ;
or ( 
    .Z ( config0_decoder7.U46.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n47 ) ) ;
and ( 
    .Z ( config0_decoder7.U46.ZN ) ,
    .I0 ( config0_decoder7.U46.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_11 ) ,
    .IN ( config0_decoder7.U46.ZN ) ) ;
and ( 
    .Z ( config0_decoder7.n40 ) ,
    .I0 ( masks_hold_reg_5_1 ) ,
    .I1 ( masks_hold_reg_5_0 ) ) ;
nor ( 
    .Z ( config0_decoder7.n35 ) ,
    .I0 ( masks_hold_reg_5_3 ) ,
    .I1 ( masks_hold_reg_5_4 ) ) ;
nand ( 
    .Z ( config0_decoder7.n58 ) ,
    .I0 ( config0_decoder7.n40 ) ,
    .I1 ( config0_decoder7.n39 ) ) ;
or ( 
    .Z ( config0_decoder7.U38.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n47 ) ) ;
and ( 
    .Z ( config0_decoder7.U38.ZN ) ,
    .I0 ( config0_decoder7.U38.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_12 ) ,
    .IN ( config0_decoder7.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U35.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U35.ZN ) ,
    .I0 ( config0_decoder7.U35.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_26 ) ,
    .IN ( config0_decoder7.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U2.AB ) ,
    .I0 ( config0_decoder7.n53 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U2.ZN ) ,
    .I0 ( config0_decoder7.U2.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_31 ) ,
    .IN ( config0_decoder7.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U81.AB ) ,
    .I0 ( config0_decoder7.n55 ) ,
    .I1 ( config0_decoder7.n53 ) ) ;
and ( 
    .Z ( config0_decoder7.U81.ZN ) ,
    .I0 ( config0_decoder7.U81.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_47 ) ,
    .IN ( config0_decoder7.U81.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n44 ) ,
    .I0 ( config0_decoder7.n37 ) ,
    .I1 ( masks_hold_reg_6_10 ) ) ;
or ( 
    .Z ( config0_decoder7.U49.AB ) ,
    .I0 ( config0_decoder7.n47 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U49.ZN ) ,
    .I0 ( config0_decoder7.U49.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_27 ) ,
    .IN ( config0_decoder7.U49.ZN ) ) ;
not ( 
    .O1 ( config0_decoder7.n36 ) ,
    .IN ( masks_hold_reg_5_3 ) ) ;
nor ( 
    .Z ( config0_decoder7.n38 ) ,
    .I0 ( masks_hold_reg_5_1 ) ,
    .I1 ( masks_hold_reg_5_2 ) ) ;
nor ( 
    .Z ( config0_decoder7.n52 ) ,
    .I0 ( config0_decoder7.n45 ) ,
    .I1 ( config0_decoder7.n36 ) ) ;
or ( 
    .Z ( config0_decoder7.U39.AB ) ,
    .I0 ( config0_decoder7.n54 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U39.ZN ) ,
    .I0 ( config0_decoder7.U39.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_18 ) ,
    .IN ( config0_decoder7.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U32.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n59 ) ) ;
and ( 
    .Z ( config0_decoder7.U32.ZN ) ,
    .I0 ( config0_decoder7.U32.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_10 ) ,
    .IN ( config0_decoder7.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U29.AB ) ,
    .I0 ( config0_decoder7.n60 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U29.ZN ) ,
    .I0 ( config0_decoder7.U29.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_24 ) ,
    .IN ( config0_decoder7.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U80.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n54 ) ) ;
and ( 
    .Z ( config0_decoder7.U80.ZN ) ,
    .I0 ( config0_decoder7.U80.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_1 ) ,
    .IN ( config0_decoder7.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U48.AB ) ,
    .I0 ( config0_decoder7.n56 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U48.ZN ) ,
    .I0 ( config0_decoder7.U48.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_35 ) ,
    .IN ( config0_decoder7.U48.ZN ) ) ;
not ( 
    .O1 ( config0_decoder7.n51 ) ,
    .IN ( masks_hold_reg_6_10 ) ) ;
nand ( 
    .Z ( config0_decoder7.n55 ) ,
    .I0 ( config0_decoder7.n52 ) ,
    .I1 ( config0_decoder7.n51 ) ) ;
or ( 
    .Z ( config0_decoder7.U33.AB ) ,
    .I0 ( config0_decoder7.n53 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U33.ZN ) ,
    .I0 ( config0_decoder7.U33.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_16 ) ,
    .IN ( config0_decoder7.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U28.AB ) ,
    .I0 ( config0_decoder7.n53 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U28.ZN ) ,
    .I0 ( config0_decoder7.U28.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_32 ) ,
    .IN ( config0_decoder7.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U83.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U83.ZN ) ,
    .I0 ( config0_decoder7.U83.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_42 ) ,
    .IN ( config0_decoder7.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U50.AB ) ,
    .I0 ( config0_decoder7.n60 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U50.ZN ) ,
    .I0 ( config0_decoder7.U50.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_39 ) ,
    .IN ( config0_decoder7.U50.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U30.AB ) ,
    .I0 ( config0_decoder7.n56 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U30.ZN ) ,
    .I0 ( config0_decoder7.U30.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_36 ) ,
    .IN ( config0_decoder7.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U22.AB ) ,
    .I0 ( config0_decoder7.n56 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U22.ZN ) ,
    .I0 ( config0_decoder7.U22.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_20 ) ,
    .IN ( config0_decoder7.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U82.AB ) ,
    .I0 ( config0_decoder7.n60 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U82.ZN ) ,
    .I0 ( config0_decoder7.U82.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_40 ) ,
    .IN ( config0_decoder7.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U51.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n62 ) ) ;
and ( 
    .Z ( config0_decoder7.U51.ZN ) ,
    .I0 ( config0_decoder7.U51.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_9 ) ,
    .IN ( config0_decoder7.U51.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U41.AB ) ,
    .I0 ( config0_decoder7.n54 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U41.ZN ) ,
    .I0 ( config0_decoder7.U41.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_33 ) ,
    .IN ( config0_decoder7.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U78.AB ) ,
    .I0 ( config0_decoder7.n49 ) ,
    .I1 ( config0_decoder7.n47 ) ) ;
and ( 
    .Z ( config0_decoder7.U78.ZN ) ,
    .I0 ( config0_decoder7.U78.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_44 ) ,
    .IN ( config0_decoder7.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U31.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n50 ) ) ;
and ( 
    .Z ( config0_decoder7.U31.ZN ) ,
    .I0 ( config0_decoder7.U31.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_14 ) ,
    .IN ( config0_decoder7.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U21.AB ) ,
    .I0 ( config0_decoder7.n55 ) ,
    .I1 ( config0_decoder7.n54 ) ) ;
and ( 
    .Z ( config0_decoder7.U21.ZN ) ,
    .I0 ( config0_decoder7.U21.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_49 ) ,
    .IN ( config0_decoder7.U21.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U5.AB ) ,
    .I0 ( config0_decoder7.n60 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U5.ZN ) ,
    .I0 ( config0_decoder7.U5.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_23 ) ,
    .IN ( config0_decoder7.U5.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U52.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n50 ) ) ;
and ( 
    .Z ( config0_decoder7.U52.ZN ) ,
    .I0 ( config0_decoder7.U52.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_13 ) ,
    .IN ( config0_decoder7.U52.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U40.AB ) ,
    .I0 ( config0_decoder7.n50 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U40.ZN ) ,
    .I0 ( config0_decoder7.U40.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_29 ) ,
    .IN ( config0_decoder7.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U79.AB ) ,
    .I0 ( config0_decoder7.n50 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U79.ZN ) ,
    .I0 ( config0_decoder7.U79.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_45 ) ,
    .IN ( config0_decoder7.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U72.AB ) ,
    .I0 ( config0_decoder7.n56 ) ,
    .I1 ( config0_decoder7.n55 ) ) ;
and ( 
    .Z ( config0_decoder7.U72.ZN ) ,
    .I0 ( config0_decoder7.U72.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_51 ) ,
    .IN ( config0_decoder7.U72.ZN ) ) ;
nor ( 
    .Z ( config0_decoder7.n37 ) ,
    .I0 ( config0_decoder7.n36 ) ,
    .I1 ( masks_hold_reg_5_4 ) ) ;
or ( 
    .Z ( config0_decoder7.U20.AB ) ,
    .I0 ( config0_decoder7.n57 ) ,
    .I1 ( config0_decoder7.n53 ) ) ;
and ( 
    .Z ( config0_decoder7.U20.ZN ) ,
    .I0 ( config0_decoder7.U20.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_48 ) ,
    .IN ( config0_decoder7.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n53 ) ,
    .I0 ( config0_decoder7.n38 ) ,
    .I1 ( config0_decoder7.n41 ) ) ;
or ( 
    .Z ( config0_decoder7.U4.AB ) ,
    .I0 ( config0_decoder7.n58 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U4.ZN ) ,
    .I0 ( config0_decoder7.U4.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_22 ) ,
    .IN ( config0_decoder7.U4.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U53.AB ) ,
    .I0 ( config0_decoder7.n56 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U53.ZN ) ,
    .I0 ( config0_decoder7.U53.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_19 ) ,
    .IN ( config0_decoder7.U53.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U43.AB ) ,
    .I0 ( config0_decoder7.n58 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U43.ZN ) ,
    .I0 ( config0_decoder7.U43.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_37 ) ,
    .IN ( config0_decoder7.U43.ZN ) ) ;
not ( 
    .O1 ( config0_decoder7.n39 ) ,
    .IN ( masks_hold_reg_5_2 ) ) ;
not ( 
    .O1 ( config0_decoder7.n41 ) ,
    .IN ( masks_hold_reg_5_0 ) ) ;
nand ( 
    .Z ( config0_decoder7.n50 ) ,
    .I0 ( config0_decoder7.n40 ) ,
    .I1 ( masks_hold_reg_5_2 ) ) ;
or ( 
    .Z ( config0_decoder7.U14.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n58 ) ) ;
and ( 
    .Z ( config0_decoder7.U14.ZN ) ,
    .I0 ( config0_decoder7.U14.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_5 ) ,
    .IN ( config0_decoder7.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n62 ) ,
    .I0 ( config0_decoder7.n35 ) ,
    .I1 ( config0_decoder7.n51 ) ) ;
nand ( 
    .Z ( config0_decoder7.n43 ) ,
    .I0 ( config0_decoder7.n37 ) ,
    .I1 ( config0_decoder7.n51 ) ) ;
or ( 
    .Z ( config0_decoder7.U42.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U42.ZN ) ,
    .I0 ( config0_decoder7.U42.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_25 ) ,
    .IN ( config0_decoder7.U42.ZN ) ) ;
nor ( 
    .Z ( config0_decoder7.n46 ) ,
    .I0 ( config0_decoder7.n45 ) ,
    .I1 ( masks_hold_reg_5_3 ) ) ;
nand ( 
    .Z ( config0_decoder7.n63 ) ,
    .I0 ( masks_hold_reg_5_0 ) ,
    .I1 ( config0_decoder7.n42 ) ) ;
or ( 
    .Z ( config0_decoder7.U18.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n56 ) ) ;
and ( 
    .Z ( config0_decoder7.U18.ZN ) ,
    .I0 ( config0_decoder7.U18.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_3 ) ,
    .IN ( config0_decoder7.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U15.AB ) ,
    .I0 ( config0_decoder7.n62 ) ,
    .I1 ( config0_decoder7.n60 ) ) ;
and ( 
    .Z ( config0_decoder7.U15.ZN ) ,
    .I0 ( config0_decoder7.U15.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_7 ) ,
    .IN ( config0_decoder7.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n48 ) ,
    .I0 ( config0_decoder7.n46 ) ,
    .I1 ( config0_decoder7.n51 ) ) ;
or ( 
    .Z ( config0_decoder7.U85.AB ) ,
    .I0 ( config0_decoder7.n48 ) ,
    .I1 ( config0_decoder7.n47 ) ) ;
and ( 
    .Z ( config0_decoder7.U85.ZN ) ,
    .I0 ( config0_decoder7.U85.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_43 ) ,
    .IN ( config0_decoder7.U85.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n56 ) ,
    .I0 ( config0_decoder7.n41 ) ,
    .I1 ( config0_decoder7.n39 ) ,
    .I2 ( masks_hold_reg_5_1 ) ) ;
or ( 
    .Z ( config0_decoder7.U45.AB ) ,
    .I0 ( config0_decoder7.n53 ) ,
    .I1 ( config0_decoder7.n43 ) ) ;
and ( 
    .Z ( config0_decoder7.U45.ZN ) ,
    .I0 ( config0_decoder7.U45.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_15 ) ,
    .IN ( config0_decoder7.U45.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U71.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n56 ) ) ;
and ( 
    .Z ( config0_decoder7.U71.ZN ) ,
    .I0 ( config0_decoder7.U71.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_4 ) ,
    .IN ( config0_decoder7.U71.ZN ) ) ;
nand ( 
    .Z ( config0_decoder7.n57 ) ,
    .I0 ( masks_hold_reg_6_10 ) ,
    .I1 ( config0_decoder7.n52 ) ) ;
or ( 
    .Z ( config0_decoder7.U19.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n54 ) ) ;
and ( 
    .Z ( config0_decoder7.U19.ZN ) ,
    .I0 ( config0_decoder7.U19.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_2 ) ,
    .IN ( config0_decoder7.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U16.AB ) ,
    .I0 ( config0_decoder7.n59 ) ,
    .I1 ( config0_decoder7.n58 ) ) ;
and ( 
    .Z ( config0_decoder7.U16.ZN ) ,
    .I0 ( config0_decoder7.U16.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_6 ) ,
    .IN ( config0_decoder7.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U36.AB ) ,
    .I0 ( config0_decoder7.n58 ) ,
    .I1 ( config0_decoder7.n49 ) ) ;
and ( 
    .Z ( config0_decoder7.U36.ZN ) ,
    .I0 ( config0_decoder7.U36.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_38 ) ,
    .IN ( config0_decoder7.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U1.AB ) ,
    .I0 ( config0_decoder7.n47 ) ,
    .I1 ( config0_decoder7.n44 ) ) ;
and ( 
    .Z ( config0_decoder7.U1.ZN ) ,
    .I0 ( config0_decoder7.U1.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_28 ) ,
    .IN ( config0_decoder7.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder7.U84.AB ) ,
    .I0 ( config0_decoder7.n63 ) ,
    .I1 ( config0_decoder7.n48 ) ) ;
and ( 
    .Z ( config0_decoder7.U84.ZN ) ,
    .I0 ( config0_decoder7.U84.AB ) ,
    .I1 ( config0_decoder7.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_6_41 ) ,
    .IN ( config0_decoder7.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U28.AB ) ,
    .I0 ( config0_decoder6.n40 ) ,
    .I1 ( masks_hold_reg_4_1 ) ) ;
and ( 
    .Z ( config0_decoder6.U28.ZN ) ,
    .I0 ( config0_decoder6.U28.AB ) ,
    .I1 ( config0_decoder6.n52 ) ) ;
not ( 
    .O1 ( config0_decoder6.n1 ) ,
    .IN ( config0_decoder6.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U56.AB ) ,
    .I0 ( config0_decoder6.n53 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U56.ZN ) ,
    .I0 ( config0_decoder6.U56.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_32 ) ,
    .IN ( config0_decoder6.U56.ZN ) ) ;
not ( 
    .O1 ( config0_decoder6.n41 ) ,
    .IN ( masks_hold_reg_5_10 ) ) ;
or ( 
    .Z ( config0_decoder6.U76.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n47 ) ) ;
and ( 
    .Z ( config0_decoder6.U76.ZN ) ,
    .I0 ( config0_decoder6.U76.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_11 ) ,
    .IN ( config0_decoder6.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U60.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n59 ) ) ;
and ( 
    .Z ( config0_decoder6.U60.ZN ) ,
    .I0 ( config0_decoder6.U60.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_10 ) ,
    .IN ( config0_decoder6.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U17.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n56 ) ) ;
and ( 
    .Z ( config0_decoder6.U17.ZN ) ,
    .I0 ( config0_decoder6.U17.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_3 ) ,
    .IN ( config0_decoder6.U17.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n57 ) ,
    .I0 ( masks_hold_reg_5_9 ) ,
    .I1 ( config0_decoder6.n52 ) ) ;
or ( 
    .Z ( config0_decoder6.U87.AB ) ,
    .I0 ( config0_decoder6.n57 ) ,
    .I1 ( config0_decoder6.n54 ) ) ;
and ( 
    .Z ( config0_decoder6.U87.ZN ) ,
    .I0 ( config0_decoder6.U87.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_50 ) ,
    .IN ( config0_decoder6.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U57.AB ) ,
    .I0 ( config0_decoder6.n56 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U57.ZN ) ,
    .I0 ( config0_decoder6.U57.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_36 ) ,
    .IN ( config0_decoder6.U57.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U47.AB ) ,
    .I0 ( config0_decoder6.n55 ) ,
    .I1 ( config0_decoder6.n53 ) ) ;
and ( 
    .Z ( config0_decoder6.U47.ZN ) ,
    .I0 ( config0_decoder6.U47.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_47 ) ,
    .IN ( config0_decoder6.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U77.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U77.ZN ) ,
    .I0 ( config0_decoder6.U77.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_41 ) ,
    .IN ( config0_decoder6.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U67.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n47 ) ) ;
and ( 
    .Z ( config0_decoder6.U67.ZN ) ,
    .I0 ( config0_decoder6.U67.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_12 ) ,
    .IN ( config0_decoder6.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U10.AB ) ,
    .I0 ( config0_decoder6.n50 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U10.ZN ) ,
    .I0 ( config0_decoder6.U10.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_30 ) ,
    .IN ( config0_decoder6.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n44 ) ,
    .I0 ( config0_decoder6.n37 ) ,
    .I1 ( masks_hold_reg_5_9 ) ) ;
or ( 
    .Z ( config0_decoder6.U26.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n56 ) ) ;
and ( 
    .Z ( config0_decoder6.U26.ZN ) ,
    .I0 ( config0_decoder6.U26.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_4 ) ,
    .IN ( config0_decoder6.U26.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n62 ) ,
    .I0 ( config0_decoder6.n35 ) ,
    .I1 ( config0_decoder6.n51 ) ) ;
or ( 
    .Z ( config0_decoder6.U86.AB ) ,
    .I0 ( config0_decoder6.n57 ) ,
    .I1 ( config0_decoder6.n56 ) ) ;
and ( 
    .Z ( config0_decoder6.U86.ZN ) ,
    .I0 ( config0_decoder6.U86.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_52 ) ,
    .IN ( config0_decoder6.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U58.AB ) ,
    .I0 ( config0_decoder6.n56 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U58.ZN ) ,
    .I0 ( config0_decoder6.U58.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_20 ) ,
    .IN ( config0_decoder6.U58.ZN ) ) ;
not ( 
    .O1 ( config0_decoder6.n45 ) ,
    .IN ( masks_hold_reg_4_3 ) ) ;
or ( 
    .Z ( config0_decoder6.U74.AB ) ,
    .I0 ( config0_decoder6.n58 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U74.ZN ) ,
    .I0 ( config0_decoder6.U74.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_21 ) ,
    .IN ( config0_decoder6.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U66.AB ) ,
    .I0 ( config0_decoder6.n60 ) ,
    .I1 ( config0_decoder6.n59 ) ) ;
and ( 
    .Z ( config0_decoder6.U66.ZN ) ,
    .I0 ( config0_decoder6.U66.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_8 ) ,
    .IN ( config0_decoder6.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U11.AB ) ,
    .I0 ( config0_decoder6.n53 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U11.ZN ) ,
    .I0 ( config0_decoder6.U11.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_31 ) ,
    .IN ( config0_decoder6.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder6.n38 ) ,
    .I0 ( masks_hold_reg_4_0 ) ,
    .I1 ( masks_hold_reg_4_1 ) ) ;
nand ( 
    .Z ( config0_decoder6.n63 ) ,
    .I0 ( masks_hold_reg_5_10 ) ,
    .I1 ( config0_decoder6.n42 ) ) ;
nand ( 
    .Z ( config0_decoder6.n43 ) ,
    .I0 ( config0_decoder6.n37 ) ,
    .I1 ( config0_decoder6.n51 ) ) ;
or ( 
    .Z ( config0_decoder6.U81.AB ) ,
    .I0 ( config0_decoder6.n60 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U81.ZN ) ,
    .I0 ( config0_decoder6.U81.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_23 ) ,
    .IN ( config0_decoder6.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U59.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n50 ) ) ;
and ( 
    .Z ( config0_decoder6.U59.ZN ) ,
    .I0 ( config0_decoder6.U59.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_14 ) ,
    .IN ( config0_decoder6.U59.ZN ) ) ;
and ( 
    .Z ( config0_decoder6.n40 ) ,
    .I0 ( masks_hold_reg_4_0 ) ,
    .I1 ( masks_hold_reg_5_10 ) ) ;
or ( 
    .Z ( config0_decoder6.U75.AB ) ,
    .I0 ( config0_decoder6.n53 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U75.ZN ) ,
    .I0 ( config0_decoder6.U75.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_15 ) ,
    .IN ( config0_decoder6.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U65.AB ) ,
    .I0 ( config0_decoder6.n58 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U65.ZN ) ,
    .I0 ( config0_decoder6.U65.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_22 ) ,
    .IN ( config0_decoder6.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U12.AB ) ,
    .I0 ( config0_decoder6.n53 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U12.ZN ) ,
    .I0 ( config0_decoder6.U12.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_16 ) ,
    .IN ( config0_decoder6.U12.ZN ) ) ;
not ( 
    .O1 ( config0_decoder6.n51 ) ,
    .IN ( masks_hold_reg_5_9 ) ) ;
nand ( 
    .Z ( config0_decoder6.n49 ) ,
    .I0 ( config0_decoder6.n46 ) ,
    .I1 ( masks_hold_reg_5_9 ) ) ;
nand ( 
    .Z ( config0_decoder6.n56 ) ,
    .I0 ( config0_decoder6.n41 ) ,
    .I1 ( config0_decoder6.n39 ) ,
    .I2 ( masks_hold_reg_4_0 ) ) ;
or ( 
    .Z ( config0_decoder6.U80.AB ) ,
    .I0 ( config0_decoder6.n60 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U80.ZN ) ,
    .I0 ( config0_decoder6.U80.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_39 ) ,
    .IN ( config0_decoder6.U80.ZN ) ) ;
not ( 
    .O1 ( config0_decoder6.n36 ) ,
    .IN ( masks_hold_reg_4_2 ) ) ;
or ( 
    .Z ( config0_decoder6.U64.AB ) ,
    .I0 ( config0_decoder6.n58 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U64.ZN ) ,
    .I0 ( config0_decoder6.U64.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_38 ) ,
    .IN ( config0_decoder6.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U13.AB ) ,
    .I0 ( config0_decoder6.n54 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U13.ZN ) ,
    .I0 ( config0_decoder6.U13.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_18 ) ,
    .IN ( config0_decoder6.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n54 ) ,
    .I0 ( config0_decoder6.n38 ) ,
    .I1 ( masks_hold_reg_5_10 ) ) ;
or ( 
    .Z ( config0_decoder6.U83.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n50 ) ) ;
and ( 
    .Z ( config0_decoder6.U83.ZN ) ,
    .I0 ( config0_decoder6.U83.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_13 ) ,
    .IN ( config0_decoder6.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U50.AB ) ,
    .I0 ( config0_decoder6.n50 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U50.ZN ) ,
    .I0 ( config0_decoder6.U50.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_46 ) ,
    .IN ( config0_decoder6.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n47 ) ,
    .I0 ( masks_hold_reg_4_1 ) ,
    .I1 ( config0_decoder6.n41 ) ,
    .I2 ( masks_hold_reg_4_0 ) ) ;
or ( 
    .Z ( config0_decoder6.U82.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n62 ) ) ;
and ( 
    .Z ( config0_decoder6.U82.ZN ) ,
    .I0 ( config0_decoder6.U82.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_9 ) ,
    .IN ( config0_decoder6.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U51.AB ) ,
    .I0 ( config0_decoder6.n49 ) ,
    .I1 ( config0_decoder6.n47 ) ) ;
and ( 
    .Z ( config0_decoder6.U51.ZN ) ,
    .I0 ( config0_decoder6.U51.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_44 ) ,
    .IN ( config0_decoder6.U51.ZN ) ) ;
nor ( 
    .Z ( config0_decoder6.n37 ) ,
    .I0 ( config0_decoder6.n36 ) ,
    .I1 ( masks_hold_reg_4_3 ) ) ;
or ( 
    .Z ( config0_decoder6.U78.AB ) ,
    .I0 ( config0_decoder6.n47 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U78.ZN ) ,
    .I0 ( config0_decoder6.U78.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_27 ) ,
    .IN ( config0_decoder6.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n59 ) ,
    .I0 ( masks_hold_reg_5_9 ) ,
    .I1 ( config0_decoder6.n35 ) ) ;
or ( 
    .Z ( config0_decoder6.U21.AB ) ,
    .I0 ( config0_decoder6.n56 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U21.ZN ) ,
    .I0 ( config0_decoder6.U21.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_19 ) ,
    .IN ( config0_decoder6.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n60 ) ,
    .I0 ( config0_decoder6.n42 ) ,
    .I1 ( config0_decoder6.n41 ) ) ;
or ( 
    .Z ( config0_decoder6.U52.AB ) ,
    .I0 ( config0_decoder6.n50 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U52.ZN ) ,
    .I0 ( config0_decoder6.U52.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_45 ) ,
    .IN ( config0_decoder6.U52.ZN ) ) ;
nor ( 
    .Z ( config0_decoder6.n35 ) ,
    .I0 ( masks_hold_reg_4_2 ) ,
    .I1 ( masks_hold_reg_4_3 ) ) ;
or ( 
    .Z ( config0_decoder6.U79.AB ) ,
    .I0 ( config0_decoder6.n56 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U79.ZN ) ,
    .I0 ( config0_decoder6.U79.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_35 ) ,
    .IN ( config0_decoder6.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U72.AB ) ,
    .I0 ( config0_decoder6.n58 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U72.ZN ) ,
    .I0 ( config0_decoder6.U72.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_37 ) ,
    .IN ( config0_decoder6.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U69.AB ) ,
    .I0 ( config0_decoder6.n50 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U69.ZN ) ,
    .I0 ( config0_decoder6.U69.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_29 ) ,
    .IN ( config0_decoder6.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U20.AB ) ,
    .I0 ( config0_decoder6.n55 ) ,
    .I1 ( config0_decoder6.n54 ) ) ;
and ( 
    .Z ( config0_decoder6.U20.ZN ) ,
    .I0 ( config0_decoder6.U20.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_49 ) ,
    .IN ( config0_decoder6.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U9.AB ) ,
    .I0 ( config0_decoder6.n47 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U9.ZN ) ,
    .I0 ( config0_decoder6.U9.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_28 ) ,
    .IN ( config0_decoder6.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n53 ) ,
    .I0 ( config0_decoder6.n38 ) ,
    .I1 ( config0_decoder6.n41 ) ) ;
or ( 
    .Z ( config0_decoder6.U53.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n58 ) ) ;
and ( 
    .Z ( config0_decoder6.U53.ZN ) ,
    .I0 ( config0_decoder6.U53.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_5 ) ,
    .IN ( config0_decoder6.U53.ZN ) ) ;
not ( 
    .O1 ( config0_decoder6.n39 ) ,
    .IN ( masks_hold_reg_4_1 ) ) ;
or ( 
    .Z ( config0_decoder6.U73.AB ) ,
    .I0 ( config0_decoder6.n54 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U73.ZN ) ,
    .I0 ( config0_decoder6.U73.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_17 ) ,
    .IN ( config0_decoder6.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U68.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U68.ZN ) ,
    .I0 ( config0_decoder6.U68.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_42 ) ,
    .IN ( config0_decoder6.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U63.AB ) ,
    .I0 ( config0_decoder6.n54 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U63.ZN ) ,
    .I0 ( config0_decoder6.U63.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_34 ) ,
    .IN ( config0_decoder6.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U14.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n60 ) ) ;
and ( 
    .Z ( config0_decoder6.U14.ZN ) ,
    .I0 ( config0_decoder6.U14.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_7 ) ,
    .IN ( config0_decoder6.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n55 ) ,
    .I0 ( config0_decoder6.n52 ) ,
    .I1 ( config0_decoder6.n51 ) ) ;
nor ( 
    .Z ( config0_decoder6.n52 ) ,
    .I0 ( config0_decoder6.n45 ) ,
    .I1 ( config0_decoder6.n36 ) ) ;
or ( 
    .Z ( config0_decoder6.U54.AB ) ,
    .I0 ( config0_decoder6.n62 ) ,
    .I1 ( config0_decoder6.n54 ) ) ;
and ( 
    .Z ( config0_decoder6.U54.ZN ) ,
    .I0 ( config0_decoder6.U54.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_1 ) ,
    .IN ( config0_decoder6.U54.ZN ) ) ;
nor ( 
    .Z ( config0_decoder6.n42 ) ,
    .I0 ( config0_decoder6.n39 ) ,
    .I1 ( masks_hold_reg_4_0 ) ) ;
or ( 
    .Z ( config0_decoder6.U70.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n43 ) ) ;
and ( 
    .Z ( config0_decoder6.U70.ZN ) ,
    .I0 ( config0_decoder6.U70.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_25 ) ,
    .IN ( config0_decoder6.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U62.AB ) ,
    .I0 ( config0_decoder6.n63 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U62.ZN ) ,
    .I0 ( config0_decoder6.U62.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_26 ) ,
    .IN ( config0_decoder6.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U18.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n54 ) ) ;
and ( 
    .Z ( config0_decoder6.U18.ZN ) ,
    .I0 ( config0_decoder6.U18.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_2 ) ,
    .IN ( config0_decoder6.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U15.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n58 ) ) ;
and ( 
    .Z ( config0_decoder6.U15.ZN ) ,
    .I0 ( config0_decoder6.U15.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_6 ) ,
    .IN ( config0_decoder6.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n58 ) ,
    .I0 ( config0_decoder6.n40 ) ,
    .I1 ( config0_decoder6.n39 ) ) ;
or ( 
    .Z ( config0_decoder6.U85.AB ) ,
    .I0 ( config0_decoder6.n56 ) ,
    .I1 ( config0_decoder6.n55 ) ) ;
and ( 
    .Z ( config0_decoder6.U85.ZN ) ,
    .I0 ( config0_decoder6.U85.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_51 ) ,
    .IN ( config0_decoder6.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U55.AB ) ,
    .I0 ( config0_decoder6.n60 ) ,
    .I1 ( config0_decoder6.n44 ) ) ;
and ( 
    .Z ( config0_decoder6.U55.ZN ) ,
    .I0 ( config0_decoder6.U55.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_24 ) ,
    .IN ( config0_decoder6.U55.ZN ) ) ;
nor ( 
    .Z ( config0_decoder6.n46 ) ,
    .I0 ( config0_decoder6.n45 ) ,
    .I1 ( masks_hold_reg_4_2 ) ) ;
or ( 
    .Z ( config0_decoder6.U71.AB ) ,
    .I0 ( config0_decoder6.n54 ) ,
    .I1 ( config0_decoder6.n48 ) ) ;
and ( 
    .Z ( config0_decoder6.U71.ZN ) ,
    .I0 ( config0_decoder6.U71.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_33 ) ,
    .IN ( config0_decoder6.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U61.AB ) ,
    .I0 ( config0_decoder6.n60 ) ,
    .I1 ( config0_decoder6.n49 ) ) ;
and ( 
    .Z ( config0_decoder6.U61.ZN ) ,
    .I0 ( config0_decoder6.U61.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_40 ) ,
    .IN ( config0_decoder6.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U19.AB ) ,
    .I0 ( config0_decoder6.n57 ) ,
    .I1 ( config0_decoder6.n53 ) ) ;
and ( 
    .Z ( config0_decoder6.U19.ZN ) ,
    .I0 ( config0_decoder6.U19.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_48 ) ,
    .IN ( config0_decoder6.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder6.U16.AB ) ,
    .I0 ( config0_decoder6.n59 ) ,
    .I1 ( config0_decoder6.n53 ) ) ;
and ( 
    .Z ( config0_decoder6.U16.ZN ) ,
    .I0 ( config0_decoder6.U16.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_0 ) ,
    .IN ( config0_decoder6.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder6.n50 ) ,
    .I0 ( config0_decoder6.n40 ) ,
    .I1 ( masks_hold_reg_4_1 ) ) ;
nand ( 
    .Z ( config0_decoder6.n48 ) ,
    .I0 ( config0_decoder6.n46 ) ,
    .I1 ( config0_decoder6.n51 ) ) ;
or ( 
    .Z ( config0_decoder6.U84.AB ) ,
    .I0 ( config0_decoder6.n48 ) ,
    .I1 ( config0_decoder6.n47 ) ) ;
and ( 
    .Z ( config0_decoder6.U84.ZN ) ,
    .I0 ( config0_decoder6.U84.AB ) ,
    .I1 ( config0_decoder6.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_5_43 ) ,
    .IN ( config0_decoder6.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U49.AB ) ,
    .I0 ( config0_decoder5.n40 ) ,
    .I1 ( masks_hold_reg_3_0 ) ) ;
and ( 
    .Z ( config0_decoder5.U49.ZN ) ,
    .I0 ( config0_decoder5.U49.AB ) ,
    .I1 ( config0_decoder5.n52 ) ) ;
not ( 
    .O1 ( config0_decoder5.n1 ) ,
    .IN ( config0_decoder5.U49.ZN ) ) ;
not ( 
    .O1 ( config0_decoder5.n36 ) ,
    .IN ( masks_hold_reg_3_1 ) ) ;
nor ( 
    .Z ( config0_decoder5.n38 ) ,
    .I0 ( masks_hold_reg_4_10 ) ,
    .I1 ( masks_hold_reg_3_0 ) ) ;
or ( 
    .Z ( config0_decoder5.U19.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n54 ) ) ;
and ( 
    .Z ( config0_decoder5.U19.ZN ) ,
    .I0 ( config0_decoder5.U19.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_2 ) ,
    .IN ( config0_decoder5.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U16.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n58 ) ) ;
and ( 
    .Z ( config0_decoder5.U16.ZN ) ,
    .I0 ( config0_decoder5.U16.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_6 ) ,
    .IN ( config0_decoder5.U16.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U36.AB ) ,
    .I0 ( config0_decoder5.n50 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U36.ZN ) ,
    .I0 ( config0_decoder5.U36.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_29 ) ,
    .IN ( config0_decoder5.U36.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U1.AB ) ,
    .I0 ( config0_decoder5.n47 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U1.ZN ) ,
    .I0 ( config0_decoder5.U1.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_28 ) ,
    .IN ( config0_decoder5.U1.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U84.AB ) ,
    .I0 ( config0_decoder5.n48 ) ,
    .I1 ( config0_decoder5.n47 ) ) ;
and ( 
    .Z ( config0_decoder5.U84.ZN ) ,
    .I0 ( config0_decoder5.U84.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_43 ) ,
    .IN ( config0_decoder5.U84.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n63 ) ,
    .I0 ( n92 ) ,
    .I1 ( config0_decoder5.n42 ) ) ;
or ( 
    .Z ( config0_decoder5.U44.AB ) ,
    .I0 ( config0_decoder5.n56 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U44.ZN ) ,
    .I0 ( config0_decoder5.U44.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_35 ) ,
    .IN ( config0_decoder5.U44.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U76.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n59 ) ) ;
and ( 
    .Z ( config0_decoder5.U76.ZN ) ,
    .I0 ( config0_decoder5.U76.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_10 ) ,
    .IN ( config0_decoder5.U76.ZN ) ) ;
not ( 
    .O1 ( config0_decoder5.n41 ) ,
    .IN ( n92 ) ) ;
or ( 
    .Z ( config0_decoder5.U17.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n53 ) ) ;
and ( 
    .Z ( config0_decoder5.U17.ZN ) ,
    .I0 ( config0_decoder5.U17.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_0 ) ,
    .IN ( config0_decoder5.U17.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U37.AB ) ,
    .I0 ( config0_decoder5.n54 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U37.ZN ) ,
    .I0 ( config0_decoder5.U37.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_33 ) ,
    .IN ( config0_decoder5.U37.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U87.AB ) ,
    .I0 ( config0_decoder5.n57 ) ,
    .I1 ( config0_decoder5.n54 ) ) ;
and ( 
    .Z ( config0_decoder5.U87.ZN ) ,
    .I0 ( config0_decoder5.U87.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_50 ) ,
    .IN ( config0_decoder5.U87.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n57 ) ,
    .I0 ( masks_hold_reg_4_8 ) ,
    .I1 ( config0_decoder5.n52 ) ) ;
or ( 
    .Z ( config0_decoder5.U47.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n62 ) ) ;
and ( 
    .Z ( config0_decoder5.U47.ZN ) ,
    .I0 ( config0_decoder5.U47.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_9 ) ,
    .IN ( config0_decoder5.U47.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U77.AB ) ,
    .I0 ( config0_decoder5.n53 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U77.ZN ) ,
    .I0 ( config0_decoder5.U77.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_16 ) ,
    .IN ( config0_decoder5.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U67.AB ) ,
    .I0 ( config0_decoder5.n49 ) ,
    .I1 ( config0_decoder5.n47 ) ) ;
and ( 
    .Z ( config0_decoder5.U67.ZN ) ,
    .I0 ( config0_decoder5.U67.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_44 ) ,
    .IN ( config0_decoder5.U67.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n58 ) ,
    .I0 ( config0_decoder5.n40 ) ,
    .I1 ( config0_decoder5.n39 ) ) ;
or ( 
    .Z ( config0_decoder5.U34.AB ) ,
    .I0 ( config0_decoder5.n58 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U34.ZN ) ,
    .I0 ( config0_decoder5.U34.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_38 ) ,
    .IN ( config0_decoder5.U34.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U3.AB ) ,
    .I0 ( config0_decoder5.n50 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U3.ZN ) ,
    .I0 ( config0_decoder5.U3.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_30 ) ,
    .IN ( config0_decoder5.U3.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U86.AB ) ,
    .I0 ( config0_decoder5.n57 ) ,
    .I1 ( config0_decoder5.n56 ) ) ;
and ( 
    .Z ( config0_decoder5.U86.ZN ) ,
    .I0 ( config0_decoder5.U86.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_52 ) ,
    .IN ( config0_decoder5.U86.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n50 ) ,
    .I0 ( config0_decoder5.n40 ) ,
    .I1 ( masks_hold_reg_3_0 ) ) ;
or ( 
    .Z ( config0_decoder5.U46.AB ) ,
    .I0 ( config0_decoder5.n60 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U46.ZN ) ,
    .I0 ( config0_decoder5.U46.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_39 ) ,
    .IN ( config0_decoder5.U46.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U74.AB ) ,
    .I0 ( config0_decoder5.n50 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U74.ZN ) ,
    .I0 ( config0_decoder5.U74.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_45 ) ,
    .IN ( config0_decoder5.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U66.AB ) ,
    .I0 ( config0_decoder5.n55 ) ,
    .I1 ( config0_decoder5.n53 ) ) ;
and ( 
    .Z ( config0_decoder5.U66.ZN ) ,
    .I0 ( config0_decoder5.U66.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_47 ) ,
    .IN ( config0_decoder5.U66.ZN ) ) ;
nor ( 
    .Z ( config0_decoder5.n52 ) ,
    .I0 ( config0_decoder5.n45 ) ,
    .I1 ( config0_decoder5.n36 ) ) ;
or ( 
    .Z ( config0_decoder5.U38.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U38.ZN ) ,
    .I0 ( config0_decoder5.U38.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_25 ) ,
    .IN ( config0_decoder5.U38.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U35.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n47 ) ) ;
and ( 
    .Z ( config0_decoder5.U35.ZN ) ,
    .I0 ( config0_decoder5.U35.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_12 ) ,
    .IN ( config0_decoder5.U35.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U2.AB ) ,
    .I0 ( config0_decoder5.n53 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U2.ZN ) ,
    .I0 ( config0_decoder5.U2.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_31 ) ,
    .IN ( config0_decoder5.U2.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U81.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U81.ZN ) ,
    .I0 ( config0_decoder5.U81.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_42 ) ,
    .IN ( config0_decoder5.U81.ZN ) ) ;
not ( 
    .O1 ( config0_decoder5.n51 ) ,
    .IN ( masks_hold_reg_4_8 ) ) ;
or ( 
    .Z ( config0_decoder5.U75.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n54 ) ) ;
and ( 
    .Z ( config0_decoder5.U75.ZN ) ,
    .I0 ( config0_decoder5.U75.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_1 ) ,
    .IN ( config0_decoder5.U75.ZN ) ) ;
nor ( 
    .Z ( config0_decoder5.n46 ) ,
    .I0 ( config0_decoder5.n45 ) ,
    .I1 ( masks_hold_reg_3_1 ) ) ;
nand ( 
    .Z ( config0_decoder5.n55 ) ,
    .I0 ( config0_decoder5.n52 ) ,
    .I1 ( config0_decoder5.n51 ) ) ;
or ( 
    .Z ( config0_decoder5.U39.AB ) ,
    .I0 ( config0_decoder5.n58 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U39.ZN ) ,
    .I0 ( config0_decoder5.U39.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_37 ) ,
    .IN ( config0_decoder5.U39.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U32.AB ) ,
    .I0 ( config0_decoder5.n54 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U32.ZN ) ,
    .I0 ( config0_decoder5.U32.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_34 ) ,
    .IN ( config0_decoder5.U32.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U29.AB ) ,
    .I0 ( config0_decoder5.n60 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U29.ZN ) ,
    .I0 ( config0_decoder5.U29.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_24 ) ,
    .IN ( config0_decoder5.U29.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U80.AB ) ,
    .I0 ( config0_decoder5.n54 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U80.ZN ) ,
    .I0 ( config0_decoder5.U80.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_18 ) ,
    .IN ( config0_decoder5.U80.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U48.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n50 ) ) ;
and ( 
    .Z ( config0_decoder5.U48.ZN ) ,
    .I0 ( config0_decoder5.U48.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_13 ) ,
    .IN ( config0_decoder5.U48.ZN ) ) ;
nor ( 
    .Z ( config0_decoder5.n37 ) ,
    .I0 ( config0_decoder5.n36 ) ,
    .I1 ( n91 ) ) ;
or ( 
    .Z ( config0_decoder5.U13.AB ) ,
    .I0 ( config0_decoder5.n60 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U13.ZN ) ,
    .I0 ( config0_decoder5.U13.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_23 ) ,
    .IN ( config0_decoder5.U13.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U33.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U33.ZN ) ,
    .I0 ( config0_decoder5.U33.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_26 ) ,
    .IN ( config0_decoder5.U33.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U28.AB ) ,
    .I0 ( config0_decoder5.n53 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U28.ZN ) ,
    .I0 ( config0_decoder5.U28.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_32 ) ,
    .IN ( config0_decoder5.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U83.AB ) ,
    .I0 ( config0_decoder5.n56 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U83.ZN ) ,
    .I0 ( config0_decoder5.U83.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_19 ) ,
    .IN ( config0_decoder5.U83.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n56 ) ,
    .I0 ( config0_decoder5.n41 ) ,
    .I1 ( config0_decoder5.n39 ) ,
    .I2 ( masks_hold_reg_4_10 ) ) ;
or ( 
    .Z ( config0_decoder5.U30.AB ) ,
    .I0 ( config0_decoder5.n56 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U30.ZN ) ,
    .I0 ( config0_decoder5.U30.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_36 ) ,
    .IN ( config0_decoder5.U30.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U22.AB ) ,
    .I0 ( config0_decoder5.n56 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U22.ZN ) ,
    .I0 ( config0_decoder5.U22.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_20 ) ,
    .IN ( config0_decoder5.U22.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U82.AB ) ,
    .I0 ( config0_decoder5.n63 ) ,
    .I1 ( config0_decoder5.n48 ) ) ;
and ( 
    .Z ( config0_decoder5.U82.ZN ) ,
    .I0 ( config0_decoder5.U82.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_41 ) ,
    .IN ( config0_decoder5.U82.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n59 ) ,
    .I0 ( masks_hold_reg_4_8 ) ,
    .I1 ( config0_decoder5.n35 ) ) ;
or ( 
    .Z ( config0_decoder5.U41.AB ) ,
    .I0 ( config0_decoder5.n53 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U41.ZN ) ,
    .I0 ( config0_decoder5.U41.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_15 ) ,
    .IN ( config0_decoder5.U41.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U78.AB ) ,
    .I0 ( config0_decoder5.n60 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U78.ZN ) ,
    .I0 ( config0_decoder5.U78.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_40 ) ,
    .IN ( config0_decoder5.U78.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U31.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n50 ) ) ;
and ( 
    .Z ( config0_decoder5.U31.ZN ) ,
    .I0 ( config0_decoder5.U31.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_14 ) ,
    .IN ( config0_decoder5.U31.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U21.AB ) ,
    .I0 ( config0_decoder5.n55 ) ,
    .I1 ( config0_decoder5.n54 ) ) ;
and ( 
    .Z ( config0_decoder5.U21.ZN ) ,
    .I0 ( config0_decoder5.U21.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_49 ) ,
    .IN ( config0_decoder5.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n48 ) ,
    .I0 ( config0_decoder5.n46 ) ,
    .I1 ( config0_decoder5.n51 ) ) ;
nand ( 
    .Z ( config0_decoder5.n47 ) ,
    .I0 ( masks_hold_reg_3_0 ) ,
    .I1 ( config0_decoder5.n41 ) ,
    .I2 ( masks_hold_reg_4_10 ) ) ;
or ( 
    .Z ( config0_decoder5.U40.AB ) ,
    .I0 ( config0_decoder5.n58 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U40.ZN ) ,
    .I0 ( config0_decoder5.U40.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_21 ) ,
    .IN ( config0_decoder5.U40.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U79.AB ) ,
    .I0 ( config0_decoder5.n60 ) ,
    .I1 ( config0_decoder5.n59 ) ) ;
and ( 
    .Z ( config0_decoder5.U79.ZN ) ,
    .I0 ( config0_decoder5.U79.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_8 ) ,
    .IN ( config0_decoder5.U79.ZN ) ) ;
not ( 
    .O1 ( config0_decoder5.n45 ) ,
    .IN ( n91 ) ) ;
not ( 
    .O1 ( config0_decoder5.n39 ) ,
    .IN ( masks_hold_reg_3_0 ) ) ;
or ( 
    .Z ( config0_decoder5.U20.AB ) ,
    .I0 ( config0_decoder5.n57 ) ,
    .I1 ( config0_decoder5.n53 ) ) ;
and ( 
    .Z ( config0_decoder5.U20.ZN ) ,
    .I0 ( config0_decoder5.U20.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_48 ) ,
    .IN ( config0_decoder5.U20.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n60 ) ,
    .I0 ( config0_decoder5.n42 ) ,
    .I1 ( config0_decoder5.n41 ) ) ;
or ( 
    .Z ( config0_decoder5.U4.AB ) ,
    .I0 ( config0_decoder5.n58 ) ,
    .I1 ( config0_decoder5.n44 ) ) ;
and ( 
    .Z ( config0_decoder5.U4.ZN ) ,
    .I0 ( config0_decoder5.U4.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_22 ) ,
    .IN ( config0_decoder5.U4.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n54 ) ,
    .I0 ( config0_decoder5.n38 ) ,
    .I1 ( n92 ) ) ;
or ( 
    .Z ( config0_decoder5.U43.AB ) ,
    .I0 ( config0_decoder5.n54 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U43.ZN ) ,
    .I0 ( config0_decoder5.U43.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_17 ) ,
    .IN ( config0_decoder5.U43.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U73.AB ) ,
    .I0 ( config0_decoder5.n50 ) ,
    .I1 ( config0_decoder5.n49 ) ) ;
and ( 
    .Z ( config0_decoder5.U73.ZN ) ,
    .I0 ( config0_decoder5.U73.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_46 ) ,
    .IN ( config0_decoder5.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U68.AB ) ,
    .I0 ( config0_decoder5.n59 ) ,
    .I1 ( config0_decoder5.n56 ) ) ;
and ( 
    .Z ( config0_decoder5.U68.ZN ) ,
    .I0 ( config0_decoder5.U68.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_4 ) ,
    .IN ( config0_decoder5.U68.ZN ) ) ;
nor ( 
    .Z ( config0_decoder5.n35 ) ,
    .I0 ( masks_hold_reg_3_1 ) ,
    .I1 ( n91 ) ) ;
or ( 
    .Z ( config0_decoder5.U14.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n58 ) ) ;
and ( 
    .Z ( config0_decoder5.U14.ZN ) ,
    .I0 ( config0_decoder5.U14.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_5 ) ,
    .IN ( config0_decoder5.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n53 ) ,
    .I0 ( config0_decoder5.n38 ) ,
    .I1 ( config0_decoder5.n41 ) ) ;
nand ( 
    .Z ( config0_decoder5.n62 ) ,
    .I0 ( config0_decoder5.n35 ) ,
    .I1 ( config0_decoder5.n51 ) ) ;
nand ( 
    .Z ( config0_decoder5.n49 ) ,
    .I0 ( config0_decoder5.n46 ) ,
    .I1 ( masks_hold_reg_4_8 ) ) ;
or ( 
    .Z ( config0_decoder5.U42.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n47 ) ) ;
and ( 
    .Z ( config0_decoder5.U42.ZN ) ,
    .I0 ( config0_decoder5.U42.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_11 ) ,
    .IN ( config0_decoder5.U42.ZN ) ) ;
and ( 
    .Z ( config0_decoder5.n40 ) ,
    .I0 ( masks_hold_reg_4_10 ) ,
    .I1 ( n92 ) ) ;
nor ( 
    .Z ( config0_decoder5.n42 ) ,
    .I0 ( config0_decoder5.n39 ) ,
    .I1 ( masks_hold_reg_4_10 ) ) ;
or ( 
    .Z ( config0_decoder5.U18.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n56 ) ) ;
and ( 
    .Z ( config0_decoder5.U18.ZN ) ,
    .I0 ( config0_decoder5.U18.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_3 ) ,
    .IN ( config0_decoder5.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder5.U15.AB ) ,
    .I0 ( config0_decoder5.n62 ) ,
    .I1 ( config0_decoder5.n60 ) ) ;
and ( 
    .Z ( config0_decoder5.U15.ZN ) ,
    .I0 ( config0_decoder5.U15.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_7 ) ,
    .IN ( config0_decoder5.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n43 ) ,
    .I0 ( config0_decoder5.n37 ) ,
    .I1 ( config0_decoder5.n51 ) ) ;
or ( 
    .Z ( config0_decoder5.U85.AB ) ,
    .I0 ( config0_decoder5.n56 ) ,
    .I1 ( config0_decoder5.n55 ) ) ;
and ( 
    .Z ( config0_decoder5.U85.ZN ) ,
    .I0 ( config0_decoder5.U85.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_51 ) ,
    .IN ( config0_decoder5.U85.ZN ) ) ;
nand ( 
    .Z ( config0_decoder5.n44 ) ,
    .I0 ( config0_decoder5.n37 ) ,
    .I1 ( masks_hold_reg_4_8 ) ) ;
or ( 
    .Z ( config0_decoder5.U45.AB ) ,
    .I0 ( config0_decoder5.n47 ) ,
    .I1 ( config0_decoder5.n43 ) ) ;
and ( 
    .Z ( config0_decoder5.U45.ZN ) ,
    .I0 ( config0_decoder5.U45.AB ) ,
    .I1 ( config0_decoder5.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_4_27 ) ,
    .IN ( config0_decoder5.U45.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U28.AB ) ,
    .I0 ( config0_decoder4.n40 ) ,
    .I1 ( masks_hold_reg_3_10 ) ) ;
and ( 
    .Z ( config0_decoder4.U28.ZN ) ,
    .I0 ( config0_decoder4.U28.AB ) ,
    .I1 ( config0_decoder4.n52 ) ) ;
not ( 
    .O1 ( config0_decoder4.n1 ) ,
    .IN ( config0_decoder4.U28.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U46.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n54 ) ) ;
and ( 
    .Z ( config0_decoder4.U46.ZN ) ,
    .I0 ( config0_decoder4.U46.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_1 ) ,
    .IN ( config0_decoder4.U46.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U74.AB ) ,
    .I0 ( config0_decoder4.n53 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U74.ZN ) ,
    .I0 ( config0_decoder4.U74.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_15 ) ,
    .IN ( config0_decoder4.U74.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U66.AB ) ,
    .I0 ( config0_decoder4.n60 ) ,
    .I1 ( config0_decoder4.n59 ) ) ;
and ( 
    .Z ( config0_decoder4.U66.ZN ) ,
    .I0 ( config0_decoder4.U66.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_8 ) ,
    .IN ( config0_decoder4.U66.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U11.AB ) ,
    .I0 ( config0_decoder4.n56 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U11.ZN ) ,
    .I0 ( config0_decoder4.U11.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_35 ) ,
    .IN ( config0_decoder4.U11.ZN ) ) ;
nor ( 
    .Z ( config0_decoder4.n38 ) ,
    .I0 ( masks_hold_reg_3_9 ) ,
    .I1 ( masks_hold_reg_3_10 ) ) ;
nand ( 
    .Z ( config0_decoder4.n50 ) ,
    .I0 ( config0_decoder4.n40 ) ,
    .I1 ( masks_hold_reg_3_10 ) ) ;
nand ( 
    .Z ( config0_decoder4.n62 ) ,
    .I0 ( config0_decoder4.n35 ) ,
    .I1 ( config0_decoder4.n51 ) ) ;
or ( 
    .Z ( config0_decoder4.U81.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n62 ) ) ;
and ( 
    .Z ( config0_decoder4.U81.ZN ) ,
    .I0 ( config0_decoder4.U81.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_9 ) ,
    .IN ( config0_decoder4.U81.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U59.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n50 ) ) ;
and ( 
    .Z ( config0_decoder4.U59.ZN ) ,
    .I0 ( config0_decoder4.U59.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_14 ) ,
    .IN ( config0_decoder4.U59.ZN ) ) ;
and ( 
    .Z ( config0_decoder4.n40 ) ,
    .I0 ( masks_hold_reg_3_9 ) ,
    .I1 ( masks_hold_reg_3_8 ) ) ;
or ( 
    .Z ( config0_decoder4.U75.AB ) ,
    .I0 ( config0_decoder4.n54 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U75.ZN ) ,
    .I0 ( config0_decoder4.U75.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_17 ) ,
    .IN ( config0_decoder4.U75.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U65.AB ) ,
    .I0 ( config0_decoder4.n58 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U65.ZN ) ,
    .I0 ( config0_decoder4.U65.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_38 ) ,
    .IN ( config0_decoder4.U65.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U12.AB ) ,
    .I0 ( config0_decoder4.n58 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U12.ZN ) ,
    .I0 ( config0_decoder4.U12.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_22 ) ,
    .IN ( config0_decoder4.U12.ZN ) ) ;
nor ( 
    .Z ( config0_decoder4.n35 ) ,
    .I0 ( masks_hold_reg_2_0 ) ,
    .I1 ( masks_hold_reg_2_1 ) ) ;
nand ( 
    .Z ( config0_decoder4.n54 ) ,
    .I0 ( config0_decoder4.n38 ) ,
    .I1 ( masks_hold_reg_3_8 ) ) ;
nand ( 
    .Z ( config0_decoder4.n56 ) ,
    .I0 ( config0_decoder4.n41 ) ,
    .I1 ( config0_decoder4.n39 ) ,
    .I2 ( masks_hold_reg_3_9 ) ) ;
or ( 
    .Z ( config0_decoder4.U80.AB ) ,
    .I0 ( config0_decoder4.n60 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U80.ZN ) ,
    .I0 ( config0_decoder4.U80.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_39 ) ,
    .IN ( config0_decoder4.U80.ZN ) ) ;
not ( 
    .O1 ( config0_decoder4.n45 ) ,
    .IN ( masks_hold_reg_2_1 ) ) ;
or ( 
    .Z ( config0_decoder4.U64.AB ) ,
    .I0 ( config0_decoder4.n50 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U64.ZN ) ,
    .I0 ( config0_decoder4.U64.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_30 ) ,
    .IN ( config0_decoder4.U64.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U13.AB ) ,
    .I0 ( config0_decoder4.n60 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U13.ZN ) ,
    .I0 ( config0_decoder4.U13.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_23 ) ,
    .IN ( config0_decoder4.U13.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n49 ) ,
    .I0 ( config0_decoder4.n46 ) ,
    .I1 ( masks_hold_reg_3_7 ) ) ;
or ( 
    .Z ( config0_decoder4.U83.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n50 ) ) ;
and ( 
    .Z ( config0_decoder4.U83.ZN ) ,
    .I0 ( config0_decoder4.U83.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_13 ) ,
    .IN ( config0_decoder4.U83.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U50.AB ) ,
    .I0 ( config0_decoder4.n50 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U50.ZN ) ,
    .I0 ( config0_decoder4.U50.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_46 ) ,
    .IN ( config0_decoder4.U50.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n47 ) ,
    .I0 ( masks_hold_reg_3_10 ) ,
    .I1 ( config0_decoder4.n41 ) ,
    .I2 ( masks_hold_reg_3_9 ) ) ;
or ( 
    .Z ( config0_decoder4.U82.AB ) ,
    .I0 ( config0_decoder4.n56 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U82.ZN ) ,
    .I0 ( config0_decoder4.U82.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_19 ) ,
    .IN ( config0_decoder4.U82.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U51.AB ) ,
    .I0 ( config0_decoder4.n49 ) ,
    .I1 ( config0_decoder4.n47 ) ) ;
and ( 
    .Z ( config0_decoder4.U51.ZN ) ,
    .I0 ( config0_decoder4.U51.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_44 ) ,
    .IN ( config0_decoder4.U51.ZN ) ) ;
not ( 
    .O1 ( config0_decoder4.n39 ) ,
    .IN ( masks_hold_reg_3_10 ) ) ;
or ( 
    .Z ( config0_decoder4.U78.AB ) ,
    .I0 ( config0_decoder4.n47 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U78.ZN ) ,
    .I0 ( config0_decoder4.U78.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_27 ) ,
    .IN ( config0_decoder4.U78.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n59 ) ,
    .I0 ( masks_hold_reg_3_7 ) ,
    .I1 ( config0_decoder4.n35 ) ) ;
or ( 
    .Z ( config0_decoder4.U21.AB ) ,
    .I0 ( config0_decoder4.n56 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U21.ZN ) ,
    .I0 ( config0_decoder4.U21.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_20 ) ,
    .IN ( config0_decoder4.U21.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n60 ) ,
    .I0 ( config0_decoder4.n42 ) ,
    .I1 ( config0_decoder4.n41 ) ) ;
or ( 
    .Z ( config0_decoder4.U52.AB ) ,
    .I0 ( config0_decoder4.n50 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U52.ZN ) ,
    .I0 ( config0_decoder4.U52.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_45 ) ,
    .IN ( config0_decoder4.U52.ZN ) ) ;
nor ( 
    .Z ( config0_decoder4.n42 ) ,
    .I0 ( config0_decoder4.n39 ) ,
    .I1 ( masks_hold_reg_3_9 ) ) ;
or ( 
    .Z ( config0_decoder4.U79.AB ) ,
    .I0 ( config0_decoder4.n53 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U79.ZN ) ,
    .I0 ( config0_decoder4.U79.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_31 ) ,
    .IN ( config0_decoder4.U79.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U72.AB ) ,
    .I0 ( config0_decoder4.n58 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U72.ZN ) ,
    .I0 ( config0_decoder4.U72.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_37 ) ,
    .IN ( config0_decoder4.U72.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U69.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U69.ZN ) ,
    .I0 ( config0_decoder4.U69.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_42 ) ,
    .IN ( config0_decoder4.U69.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U20.AB ) ,
    .I0 ( config0_decoder4.n57 ) ,
    .I1 ( config0_decoder4.n53 ) ) ;
and ( 
    .Z ( config0_decoder4.U20.ZN ) ,
    .I0 ( config0_decoder4.U20.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_48 ) ,
    .IN ( config0_decoder4.U20.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U9.AB ) ,
    .I0 ( config0_decoder4.n54 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U9.ZN ) ,
    .I0 ( config0_decoder4.U9.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_34 ) ,
    .IN ( config0_decoder4.U9.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n53 ) ,
    .I0 ( config0_decoder4.n38 ) ,
    .I1 ( config0_decoder4.n41 ) ) ;
or ( 
    .Z ( config0_decoder4.U53.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n58 ) ) ;
and ( 
    .Z ( config0_decoder4.U53.ZN ) ,
    .I0 ( config0_decoder4.U53.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_5 ) ,
    .IN ( config0_decoder4.U53.ZN ) ) ;
nor ( 
    .Z ( config0_decoder4.n37 ) ,
    .I0 ( config0_decoder4.n36 ) ,
    .I1 ( masks_hold_reg_2_1 ) ) ;
or ( 
    .Z ( config0_decoder4.U73.AB ) ,
    .I0 ( config0_decoder4.n58 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U73.ZN ) ,
    .I0 ( config0_decoder4.U73.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_21 ) ,
    .IN ( config0_decoder4.U73.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U68.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n47 ) ) ;
and ( 
    .Z ( config0_decoder4.U68.ZN ) ,
    .I0 ( config0_decoder4.U68.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_12 ) ,
    .IN ( config0_decoder4.U68.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U63.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U63.ZN ) ,
    .I0 ( config0_decoder4.U63.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_26 ) ,
    .IN ( config0_decoder4.U63.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U14.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n56 ) ) ;
and ( 
    .Z ( config0_decoder4.U14.ZN ) ,
    .I0 ( config0_decoder4.U14.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_4 ) ,
    .IN ( config0_decoder4.U14.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n55 ) ,
    .I0 ( config0_decoder4.n52 ) ,
    .I1 ( config0_decoder4.n51 ) ) ;
nor ( 
    .Z ( config0_decoder4.n52 ) ,
    .I0 ( config0_decoder4.n45 ) ,
    .I1 ( config0_decoder4.n36 ) ) ;
or ( 
    .Z ( config0_decoder4.U54.AB ) ,
    .I0 ( config0_decoder4.n55 ) ,
    .I1 ( config0_decoder4.n53 ) ) ;
and ( 
    .Z ( config0_decoder4.U54.ZN ) ,
    .I0 ( config0_decoder4.U54.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_47 ) ,
    .IN ( config0_decoder4.U54.ZN ) ) ;
not ( 
    .O1 ( config0_decoder4.n51 ) ,
    .IN ( masks_hold_reg_3_7 ) ) ;
or ( 
    .Z ( config0_decoder4.U70.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U70.ZN ) ,
    .I0 ( config0_decoder4.U70.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_25 ) ,
    .IN ( config0_decoder4.U70.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U62.AB ) ,
    .I0 ( config0_decoder4.n60 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U62.ZN ) ,
    .I0 ( config0_decoder4.U62.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_40 ) ,
    .IN ( config0_decoder4.U62.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U18.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n56 ) ) ;
and ( 
    .Z ( config0_decoder4.U18.ZN ) ,
    .I0 ( config0_decoder4.U18.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_3 ) ,
    .IN ( config0_decoder4.U18.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U15.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n60 ) ) ;
and ( 
    .Z ( config0_decoder4.U15.ZN ) ,
    .I0 ( config0_decoder4.U15.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_7 ) ,
    .IN ( config0_decoder4.U15.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n58 ) ,
    .I0 ( config0_decoder4.n40 ) ,
    .I1 ( config0_decoder4.n39 ) ) ;
or ( 
    .Z ( config0_decoder4.U85.AB ) ,
    .I0 ( config0_decoder4.n56 ) ,
    .I1 ( config0_decoder4.n55 ) ) ;
and ( 
    .Z ( config0_decoder4.U85.ZN ) ,
    .I0 ( config0_decoder4.U85.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_51 ) ,
    .IN ( config0_decoder4.U85.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U55.AB ) ,
    .I0 ( config0_decoder4.n53 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U55.ZN ) ,
    .I0 ( config0_decoder4.U55.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_32 ) ,
    .IN ( config0_decoder4.U55.ZN ) ) ;
not ( 
    .O1 ( config0_decoder4.n41 ) ,
    .IN ( masks_hold_reg_3_8 ) ) ;
or ( 
    .Z ( config0_decoder4.U71.AB ) ,
    .I0 ( config0_decoder4.n50 ) ,
    .I1 ( config0_decoder4.n43 ) ) ;
and ( 
    .Z ( config0_decoder4.U71.ZN ) ,
    .I0 ( config0_decoder4.U71.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_29 ) ,
    .IN ( config0_decoder4.U71.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U61.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n59 ) ) ;
and ( 
    .Z ( config0_decoder4.U61.ZN ) ,
    .I0 ( config0_decoder4.U61.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_10 ) ,
    .IN ( config0_decoder4.U61.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U19.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n54 ) ) ;
and ( 
    .Z ( config0_decoder4.U19.ZN ) ,
    .I0 ( config0_decoder4.U19.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_2 ) ,
    .IN ( config0_decoder4.U19.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U16.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n58 ) ) ;
and ( 
    .Z ( config0_decoder4.U16.ZN ) ,
    .I0 ( config0_decoder4.U16.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_6 ) ,
    .IN ( config0_decoder4.U16.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n63 ) ,
    .I0 ( masks_hold_reg_3_8 ) ,
    .I1 ( config0_decoder4.n42 ) ) ;
nand ( 
    .Z ( config0_decoder4.n48 ) ,
    .I0 ( config0_decoder4.n46 ) ,
    .I1 ( config0_decoder4.n51 ) ) ;
or ( 
    .Z ( config0_decoder4.U84.AB ) ,
    .I0 ( config0_decoder4.n48 ) ,
    .I1 ( config0_decoder4.n47 ) ) ;
and ( 
    .Z ( config0_decoder4.U84.ZN ) ,
    .I0 ( config0_decoder4.U84.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_43 ) ,
    .IN ( config0_decoder4.U84.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U56.AB ) ,
    .I0 ( config0_decoder4.n60 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U56.ZN ) ,
    .I0 ( config0_decoder4.U56.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_24 ) ,
    .IN ( config0_decoder4.U56.ZN ) ) ;
nor ( 
    .Z ( config0_decoder4.n46 ) ,
    .I0 ( config0_decoder4.n45 ) ,
    .I1 ( masks_hold_reg_2_0 ) ) ;
or ( 
    .Z ( config0_decoder4.U76.AB ) ,
    .I0 ( config0_decoder4.n62 ) ,
    .I1 ( config0_decoder4.n47 ) ) ;
and ( 
    .Z ( config0_decoder4.U76.ZN ) ,
    .I0 ( config0_decoder4.U76.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_11 ) ,
    .IN ( config0_decoder4.U76.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U60.AB ) ,
    .I0 ( config0_decoder4.n53 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U60.ZN ) ,
    .I0 ( config0_decoder4.U60.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_16 ) ,
    .IN ( config0_decoder4.U60.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U17.AB ) ,
    .I0 ( config0_decoder4.n59 ) ,
    .I1 ( config0_decoder4.n53 ) ) ;
and ( 
    .Z ( config0_decoder4.U17.ZN ) ,
    .I0 ( config0_decoder4.U17.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_0 ) ,
    .IN ( config0_decoder4.U17.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n57 ) ,
    .I0 ( masks_hold_reg_3_7 ) ,
    .I1 ( config0_decoder4.n52 ) ) ;
or ( 
    .Z ( config0_decoder4.U87.AB ) ,
    .I0 ( config0_decoder4.n57 ) ,
    .I1 ( config0_decoder4.n54 ) ) ;
and ( 
    .Z ( config0_decoder4.U87.ZN ) ,
    .I0 ( config0_decoder4.U87.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_50 ) ,
    .IN ( config0_decoder4.U87.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U57.AB ) ,
    .I0 ( config0_decoder4.n47 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U57.ZN ) ,
    .I0 ( config0_decoder4.U57.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_28 ) ,
    .IN ( config0_decoder4.U57.ZN ) ) ;
not ( 
    .O1 ( config0_decoder4.n36 ) ,
    .IN ( masks_hold_reg_2_0 ) ) ;
or ( 
    .Z ( config0_decoder4.U77.AB ) ,
    .I0 ( config0_decoder4.n63 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U77.ZN ) ,
    .I0 ( config0_decoder4.U77.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_41 ) ,
    .IN ( config0_decoder4.U77.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U67.AB ) ,
    .I0 ( config0_decoder4.n54 ) ,
    .I1 ( config0_decoder4.n44 ) ) ;
and ( 
    .Z ( config0_decoder4.U67.ZN ) ,
    .I0 ( config0_decoder4.U67.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_18 ) ,
    .IN ( config0_decoder4.U67.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U10.AB ) ,
    .I0 ( config0_decoder4.n54 ) ,
    .I1 ( config0_decoder4.n48 ) ) ;
and ( 
    .Z ( config0_decoder4.U10.ZN ) ,
    .I0 ( config0_decoder4.U10.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_33 ) ,
    .IN ( config0_decoder4.U10.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n44 ) ,
    .I0 ( config0_decoder4.n37 ) ,
    .I1 ( masks_hold_reg_3_7 ) ) ;
or ( 
    .Z ( config0_decoder4.U26.AB ) ,
    .I0 ( config0_decoder4.n55 ) ,
    .I1 ( config0_decoder4.n54 ) ) ;
and ( 
    .Z ( config0_decoder4.U26.ZN ) ,
    .I0 ( config0_decoder4.U26.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_49 ) ,
    .IN ( config0_decoder4.U26.ZN ) ) ;
nand ( 
    .Z ( config0_decoder4.n43 ) ,
    .I0 ( config0_decoder4.n37 ) ,
    .I1 ( config0_decoder4.n51 ) ) ;
or ( 
    .Z ( config0_decoder4.U86.AB ) ,
    .I0 ( config0_decoder4.n57 ) ,
    .I1 ( config0_decoder4.n56 ) ) ;
and ( 
    .Z ( config0_decoder4.U86.ZN ) ,
    .I0 ( config0_decoder4.U86.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_52 ) ,
    .IN ( config0_decoder4.U86.ZN ) ) ;
or ( 
    .Z ( config0_decoder4.U58.AB ) ,
    .I0 ( config0_decoder4.n56 ) ,
    .I1 ( config0_decoder4.n49 ) ) ;
and ( 
    .Z ( config0_decoder4.U58.ZN ) ,
    .I0 ( config0_decoder4.U58.AB ) ,
    .I1 ( config0_decoder4.n1 ) ) ;
not ( 
    .O1 ( config0_onehot_decoded_masks_3_36 ) ,
    .IN ( config0_decoder4.U58.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder2.n2 ) ,
    .IN ( config1_decoder2.n1 ) ) ;
or ( 
    .Z ( config1_decoder2.U56.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U56.ZN ) ,
    .I0 ( config1_decoder2.U56.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_52 ) ,
    .IN ( config1_decoder2.U56.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.U44.BN ) ,
    .IN ( config1_decoder2.n32 ) ) ;
nand ( 
    .Z ( config1_decoder2.n13 ) ,
    .I0 ( config1_decoder2.U44.BN ) ,
    .I1 ( config1_decoder2.n20 ) ) ;
or ( 
    .Z ( config1_decoder2.U76.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U76.ZN ) ,
    .I0 ( config1_decoder2.U76.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_55 ) ,
    .IN ( config1_decoder2.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U60.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U60.ZN ) ,
    .I0 ( config1_decoder2.U60.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_33 ) ,
    .IN ( config1_decoder2.U60.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n43 ) ,
    .I0 ( config1_decoder2.n44 ) ,
    .I1 ( config1_decoder2.n38 ) ) ;
or ( 
    .Z ( config1_decoder2.U27.AB ) ,
    .I0 ( config1_decoder2.n25 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U27.ZN ) ,
    .I0 ( config1_decoder2.U27.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_75 ) ,
    .IN ( config1_decoder2.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U110.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n21 ) ) ;
and ( 
    .Z ( config1_decoder2.U110.ZN ) ,
    .I0 ( config1_decoder2.U110.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_70 ) ,
    .IN ( config1_decoder2.U110.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U100.AB ) ,
    .I0 ( config1_decoder2.n25 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U100.ZN ) ,
    .I0 ( config1_decoder2.U100.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_79 ) ,
    .IN ( config1_decoder2.U100.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U139.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U139.ZN ) ,
    .I0 ( config1_decoder2.U139.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_57 ) ,
    .IN ( config1_decoder2.U139.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n15 ) ,
    .I0 ( masks_hold_reg_2_2 ) ,
    .I1 ( masks_hold_reg_2_3 ) ) ;
nand ( 
    .Z ( config1_decoder2.n1 ) ,
    .I0 ( config1_decoder2.n20 ) ,
    .I1 ( config1_decoder2.n54 ) ) ;
or ( 
    .Z ( config1_decoder2.U13.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n19 ) ) ;
and ( 
    .Z ( config1_decoder2.U13.ZN ) ,
    .I0 ( config1_decoder2.U13.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_1 ) ,
    .IN ( config1_decoder2.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n27 ) ,
    .I0 ( config1_decoder2.n37 ) ,
    .I1 ( config1_decoder2.n50 ) ) ;
nand ( 
    .Z ( config1_decoder2.n10 ) ,
    .I0 ( config1_decoder2.n50 ) ,
    .I1 ( config1_decoder2.n36 ) ) ;
nor ( 
    .Z ( config1_decoder2.n34 ) ,
    .I0 ( config1_decoder2.n39 ) ,
    .I1 ( masks_hold_reg_2_7 ) ) ;
not ( 
    .O1 ( config1_decoder2.n47 ) ,
    .IN ( masks_hold_reg_2_4 ) ) ;
or ( 
    .Z ( config1_decoder2.U154.AB ) ,
    .I0 ( config1_decoder2.n14 ) ,
    .I1 ( config1_decoder2.n16 ) ) ;
and ( 
    .Z ( config1_decoder2.U154.ZN ) ,
    .I0 ( config1_decoder2.U154.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_95 ) ,
    .IN ( config1_decoder2.U154.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U144.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U144.ZN ) ,
    .I0 ( config1_decoder2.U144.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_47 ) ,
    .IN ( config1_decoder2.U144.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U160.AB ) ,
    .I0 ( config1_decoder2.n31 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U160.ZN ) ,
    .I0 ( config1_decoder2.U160.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_43 ) ,
    .IN ( config1_decoder2.U160.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U98.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n25 ) ) ;
and ( 
    .Z ( config1_decoder2.U98.ZN ) ,
    .I0 ( config1_decoder2.U98.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_67 ) ,
    .IN ( config1_decoder2.U98.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U83.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U83.ZN ) ,
    .I0 ( config1_decoder2.U83.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_19 ) ,
    .IN ( config1_decoder2.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U2.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U2.ZN ) ,
    .I0 ( config1_decoder2.U2.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_17 ) ,
    .IN ( config1_decoder2.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U81.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n23 ) ) ;
and ( 
    .Z ( config1_decoder2.U81.ZN ) ,
    .I0 ( config1_decoder2.U81.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_73 ) ,
    .IN ( config1_decoder2.U81.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U59.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U59.ZN ) ,
    .I0 ( config1_decoder2.U59.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_34 ) ,
    .IN ( config1_decoder2.U59.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U49.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n27 ) ) ;
and ( 
    .Z ( config1_decoder2.U49.ZN ) ,
    .I0 ( config1_decoder2.U49.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_28 ) ,
    .IN ( config1_decoder2.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U75.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U75.ZN ) ,
    .I0 ( config1_decoder2.U75.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_56 ) ,
    .IN ( config1_decoder2.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U65.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n27 ) ) ;
and ( 
    .Z ( config1_decoder2.U65.ZN ) ,
    .I0 ( config1_decoder2.U65.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_4 ) ,
    .IN ( config1_decoder2.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U12.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U12.ZN ) ,
    .I0 ( config1_decoder2.U12.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_13 ) ,
    .IN ( config1_decoder2.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n33 ) ,
    .I0 ( config1_decoder2.n35 ) ,
    .I1 ( config1_decoder2.n50 ) ) ;
nand ( 
    .Z ( config1_decoder2.n23 ) ,
    .I0 ( config1_decoder2.n34 ) ,
    .I1 ( config1_decoder2.n36 ) ) ;
nand ( 
    .Z ( config1_decoder2.n21 ) ,
    .I0 ( config1_decoder2.n34 ) ,
    .I1 ( config1_decoder2.n35 ) ) ;
or ( 
    .Z ( config1_decoder2.U24.AB ) ,
    .I0 ( config1_decoder2.n23 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U24.ZN ) ,
    .I0 ( config1_decoder2.U24.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_81 ) ,
    .IN ( config1_decoder2.U24.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U103.AB ) ,
    .I0 ( config1_decoder2.n21 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U103.ZN ) ,
    .I0 ( config1_decoder2.U103.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_82 ) ,
    .IN ( config1_decoder2.U103.ZN ) ) ;
nor ( 
    .Z ( config1_decoder2.n37 ) ,
    .I0 ( config1_decoder2.n52 ) ,
    .I1 ( masks_hold_reg_2_3 ) ) ;
nand ( 
    .Z ( config1_decoder2.n28 ) ,
    .I0 ( config1_decoder2.n48 ) ,
    .I1 ( masks_hold_reg_2_4 ) ) ;
or ( 
    .Z ( config1_decoder2.U155.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n26 ) ) ;
and ( 
    .Z ( config1_decoder2.U155.ZN ) ,
    .I0 ( config1_decoder2.U155.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_25 ) ,
    .IN ( config1_decoder2.U155.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U143.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U143.ZN ) ,
    .I0 ( config1_decoder2.U143.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_54 ) ,
    .IN ( config1_decoder2.U143.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U163.AB ) ,
    .I0 ( config1_decoder2.n18 ) ,
    .I1 ( config1_decoder2.n51 ) ) ;
and ( 
    .Z ( config1_decoder2.U163.ZN ) ,
    .I0 ( config1_decoder2.U163.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_104 ) ,
    .IN ( config1_decoder2.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U80.AB ) ,
    .I0 ( config1_decoder2.n27 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U80.ZN ) ,
    .I0 ( config1_decoder2.U80.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_20 ) ,
    .IN ( config1_decoder2.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U48.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n27 ) ) ;
and ( 
    .Z ( config1_decoder2.U48.ZN ) ,
    .I0 ( config1_decoder2.U48.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_24 ) ,
    .IN ( config1_decoder2.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U64.AB ) ,
    .I0 ( config1_decoder2.n24 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U64.ZN ) ,
    .I0 ( config1_decoder2.U64.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_76 ) ,
    .IN ( config1_decoder2.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U50.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U50.ZN ) ,
    .I0 ( config1_decoder2.U50.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_39 ) ,
    .IN ( config1_decoder2.U50.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n25 ) ,
    .I0 ( config1_decoder2.n34 ) ,
    .I1 ( config1_decoder2.n38 ) ) ;
nand ( 
    .Z ( config1_decoder2.n11 ) ,
    .I0 ( config1_decoder2.n47 ) ,
    .I1 ( config1_decoder2.n49 ) ,
    .I2 ( masks_hold_reg_2_5 ) ) ;
or ( 
    .Z ( config1_decoder2.U157.AB ) ,
    .I0 ( config1_decoder2.n21 ) ,
    .I1 ( config1_decoder2.n22 ) ) ;
and ( 
    .Z ( config1_decoder2.U157.ZN ) ,
    .I0 ( config1_decoder2.U157.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_94 ) ,
    .IN ( config1_decoder2.U157.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U145.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U145.ZN ) ,
    .I0 ( config1_decoder2.U145.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_32 ) ,
    .IN ( config1_decoder2.U145.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U161.AB ) ,
    .I0 ( config1_decoder2.n16 ) ,
    .I1 ( config1_decoder2.n18 ) ) ;
and ( 
    .Z ( config1_decoder2.U161.ZN ) ,
    .I0 ( config1_decoder2.U161.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_96 ) ,
    .IN ( config1_decoder2.U161.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U99.AB ) ,
    .I0 ( config1_decoder2.n25 ) ,
    .I1 ( config1_decoder2.n26 ) ) ;
and ( 
    .Z ( config1_decoder2.U99.ZN ) ,
    .I0 ( config1_decoder2.U99.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_87 ) ,
    .IN ( config1_decoder2.U99.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U82.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U82.ZN ) ,
    .I0 ( config1_decoder2.U82.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_27 ) ,
    .IN ( config1_decoder2.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U51.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U51.ZN ) ,
    .I0 ( config1_decoder2.U51.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_37 ) ,
    .IN ( config1_decoder2.U51.ZN ) ) ;
nor ( 
    .Z ( config1_decoder2.n20 ) ,
    .I0 ( config1_decoder2.n39 ) ,
    .I1 ( config1_decoder2.n45 ) ) ;
or ( 
    .Z ( config1_decoder2.U78.AB ) ,
    .I0 ( config1_decoder2.n17 ) ,
    .I1 ( config1_decoder2.n13 ) ) ;
and ( 
    .Z ( config1_decoder2.U78.ZN ) ,
    .I0 ( config1_decoder2.U78.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_101 ) ,
    .IN ( config1_decoder2.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n24 ) ,
    .I0 ( config1_decoder2.n34 ) ,
    .I1 ( config1_decoder2.n37 ) ) ;
or ( 
    .Z ( config1_decoder2.U115.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n21 ) ) ;
and ( 
    .Z ( config1_decoder2.U115.ZN ) ,
    .I0 ( config1_decoder2.U115.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_66 ) ,
    .IN ( config1_decoder2.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U156.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U156.ZN ) ,
    .I0 ( config1_decoder2.U156.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_21 ) ,
    .IN ( config1_decoder2.U156.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U146.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n25 ) ) ;
and ( 
    .Z ( config1_decoder2.U146.ZN ) ,
    .I0 ( config1_decoder2.U146.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_63 ) ,
    .IN ( config1_decoder2.U146.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U5.AB ) ,
    .I0 ( config1_decoder2.n31 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U5.ZN ) ,
    .I0 ( config1_decoder2.U5.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_46 ) ,
    .IN ( config1_decoder2.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U88.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U88.ZN ) ,
    .I0 ( config1_decoder2.U88.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_49 ) ,
    .IN ( config1_decoder2.U88.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U52.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U52.ZN ) ,
    .I0 ( config1_decoder2.U52.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_36 ) ,
    .IN ( config1_decoder2.U52.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n30 ) ,
    .I0 ( config1_decoder2.n38 ) ,
    .I1 ( config1_decoder2.n50 ) ) ;
or ( 
    .Z ( config1_decoder2.U79.AB ) ,
    .I0 ( config1_decoder2.n15 ) ,
    .I1 ( config1_decoder2.n13 ) ) ;
and ( 
    .Z ( config1_decoder2.U79.ZN ) ,
    .I0 ( config1_decoder2.U79.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_102 ) ,
    .IN ( config1_decoder2.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U72.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U72.ZN ) ,
    .I0 ( config1_decoder2.U72.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_60 ) ,
    .IN ( config1_decoder2.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U69.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U69.ZN ) ,
    .I0 ( config1_decoder2.U69.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_3 ) ,
    .IN ( config1_decoder2.U69.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n22 ) ,
    .I0 ( n79 ) ,
    .I1 ( config1_decoder2.n46 ) ) ;
or ( 
    .Z ( config1_decoder2.U114.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U114.ZN ) ,
    .I0 ( config1_decoder2.U114.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_62 ) ,
    .IN ( config1_decoder2.U114.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U104.AB ) ,
    .I0 ( config1_decoder2.n21 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U104.ZN ) ,
    .I0 ( config1_decoder2.U104.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_86 ) ,
    .IN ( config1_decoder2.U104.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U159.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n24 ) ) ;
and ( 
    .Z ( config1_decoder2.U159.ZN ) ,
    .I0 ( config1_decoder2.U159.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_72 ) ,
    .IN ( config1_decoder2.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U147.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n23 ) ) ;
and ( 
    .Z ( config1_decoder2.U147.ZN ) ,
    .I0 ( config1_decoder2.U147.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_69 ) ,
    .IN ( config1_decoder2.U147.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U9.AB ) ,
    .I0 ( config1_decoder2.n31 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U9.ZN ) ,
    .I0 ( config1_decoder2.U9.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_14 ) ,
    .IN ( config1_decoder2.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U4.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U4.ZN ) ,
    .I0 ( config1_decoder2.U4.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_31 ) ,
    .IN ( config1_decoder2.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U53.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U53.ZN ) ,
    .I0 ( config1_decoder2.U53.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_38 ) ,
    .IN ( config1_decoder2.U53.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n31 ) ,
    .I0 ( config1_decoder2.n46 ) ,
    .I1 ( config1_decoder2.n49 ) ) ;
or ( 
    .Z ( config1_decoder2.U73.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U73.ZN ) ,
    .I0 ( config1_decoder2.U73.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_59 ) ,
    .IN ( config1_decoder2.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U68.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n27 ) ) ;
and ( 
    .Z ( config1_decoder2.U68.ZN ) ,
    .I0 ( config1_decoder2.U68.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_0 ) ,
    .IN ( config1_decoder2.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U63.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U63.ZN ) ,
    .I0 ( config1_decoder2.U63.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_23 ) ,
    .IN ( config1_decoder2.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U14.AB ) ,
    .I0 ( config1_decoder2.n27 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U14.ZN ) ,
    .I0 ( config1_decoder2.U14.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_12 ) ,
    .IN ( config1_decoder2.U14.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n49 ) ,
    .IN ( n79 ) ) ;
nor ( 
    .Z ( config1_decoder2.n53 ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( n79 ) ) ;
or ( 
    .Z ( config1_decoder2.U108.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n24 ) ) ;
and ( 
    .Z ( config1_decoder2.U108.ZN ) ,
    .I0 ( config1_decoder2.U108.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_68 ) ,
    .IN ( config1_decoder2.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U105.AB ) ,
    .I0 ( config1_decoder2.n21 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U105.ZN ) ,
    .I0 ( config1_decoder2.U105.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_78 ) ,
    .IN ( config1_decoder2.U105.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U137.AB ) ,
    .I0 ( config1_decoder2.n13 ) ,
    .I1 ( config1_decoder2.n18 ) ) ;
and ( 
    .Z ( config1_decoder2.U137.ZN ) ,
    .I0 ( config1_decoder2.U137.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_100 ) ,
    .IN ( config1_decoder2.U137.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U158.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n11 ) ) ;
and ( 
    .Z ( config1_decoder2.U158.ZN ) ,
    .I0 ( config1_decoder2.U158.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_9 ) ,
    .IN ( config1_decoder2.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U148.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n23 ) ) ;
and ( 
    .Z ( config1_decoder2.U148.ZN ) ,
    .I0 ( config1_decoder2.U148.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_93 ) ,
    .IN ( config1_decoder2.U148.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U164.AB ) ,
    .I0 ( config1_decoder2.n17 ) ,
    .I1 ( config1_decoder2.n51 ) ) ;
and ( 
    .Z ( config1_decoder2.U164.ZN ) ,
    .I0 ( config1_decoder2.U164.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_105 ) ,
    .IN ( config1_decoder2.U164.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U8.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U8.ZN ) ,
    .I0 ( config1_decoder2.U8.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_50 ) ,
    .IN ( config1_decoder2.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U7.AB ) ,
    .I0 ( config1_decoder2.n31 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U7.ZN ) ,
    .I0 ( config1_decoder2.U7.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_44 ) ,
    .IN ( config1_decoder2.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U54.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U54.ZN ) ,
    .I0 ( config1_decoder2.U54.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_41 ) ,
    .IN ( config1_decoder2.U54.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n19 ) ,
    .I0 ( config1_decoder2.n53 ) ,
    .I1 ( config1_decoder2.n47 ) ) ;
or ( 
    .Z ( config1_decoder2.U70.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U70.ZN ) ,
    .I0 ( config1_decoder2.U70.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_2 ) ,
    .IN ( config1_decoder2.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U62.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U62.ZN ) ,
    .I0 ( config1_decoder2.U62.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_22 ) ,
    .IN ( config1_decoder2.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U15.AB ) ,
    .I0 ( config1_decoder2.n30 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U15.ZN ) ,
    .I0 ( config1_decoder2.U15.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_11 ) ,
    .IN ( config1_decoder2.U15.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n26 ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( config1_decoder2.n47 ) ,
    .I2 ( n79 ) ) ;
or ( 
    .Z ( config1_decoder2.U109.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n24 ) ) ;
and ( 
    .Z ( config1_decoder2.U109.ZN ) ,
    .I0 ( config1_decoder2.U109.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_64 ) ,
    .IN ( config1_decoder2.U109.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U106.AB ) ,
    .I0 ( config1_decoder2.n21 ) ,
    .I1 ( config1_decoder2.n26 ) ) ;
and ( 
    .Z ( config1_decoder2.U106.ZN ) ,
    .I0 ( config1_decoder2.U106.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_90 ) ,
    .IN ( config1_decoder2.U106.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n45 ) ,
    .IN ( masks_hold_reg_2_7 ) ) ;
nor ( 
    .Z ( config1_decoder2.n50 ) ,
    .I0 ( masks_hold_reg_2_7 ) ,
    .I1 ( masks_hold_reg_2_8 ) ) ;
or ( 
    .Z ( config1_decoder2.U149.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U149.ZN ) ,
    .I0 ( config1_decoder2.U149.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_30 ) ,
    .IN ( config1_decoder2.U149.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U165.AB ) ,
    .I0 ( config1_decoder2.n14 ) ,
    .I1 ( config1_decoder2.n51 ) ) ;
and ( 
    .Z ( config1_decoder2.U165.ZN ) ,
    .I0 ( config1_decoder2.U165.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_103 ) ,
    .IN ( config1_decoder2.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U95.AB ) ,
    .I0 ( config1_decoder2.n23 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U95.ZN ) ,
    .I0 ( config1_decoder2.U95.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_85 ) ,
    .IN ( config1_decoder2.U95.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U6.AB ) ,
    .I0 ( config1_decoder2.n31 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U6.ZN ) ,
    .I0 ( config1_decoder2.U6.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_45 ) ,
    .IN ( config1_decoder2.U6.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n35 ) ,
    .IN ( config1_decoder2.n15 ) ) ;
or ( 
    .Z ( config1_decoder2.U55.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U55.ZN ) ,
    .I0 ( config1_decoder2.U55.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_40 ) ,
    .IN ( config1_decoder2.U55.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U45.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n22 ) ) ;
and ( 
    .Z ( config1_decoder2.U45.ZN ) ,
    .I0 ( config1_decoder2.U45.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_29 ) ,
    .IN ( config1_decoder2.U45.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U71.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U71.ZN ) ,
    .I0 ( config1_decoder2.U71.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_58 ) ,
    .IN ( config1_decoder2.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U61.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U61.ZN ) ,
    .I0 ( config1_decoder2.U61.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_35 ) ,
    .IN ( config1_decoder2.U61.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n42 ) ,
    .I0 ( config1_decoder2.n44 ) ,
    .I1 ( config1_decoder2.n37 ) ) ;
or ( 
    .Z ( config1_decoder2.U111.AB ) ,
    .I0 ( config1_decoder2.n24 ) ,
    .I1 ( config1_decoder2.n26 ) ) ;
and ( 
    .Z ( config1_decoder2.U111.ZN ) ,
    .I0 ( config1_decoder2.U111.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_88 ) ,
    .IN ( config1_decoder2.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U107.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n21 ) ) ;
and ( 
    .Z ( config1_decoder2.U107.ZN ) ,
    .I0 ( config1_decoder2.U107.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_74 ) ,
    .IN ( config1_decoder2.U107.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n39 ) ,
    .IN ( masks_hold_reg_2_8 ) ) ;
nor ( 
    .Z ( config1_decoder2.n48 ) ,
    .I0 ( config1_decoder2.n49 ) ,
    .I1 ( masks_hold_reg_2_5 ) ) ;
or ( 
    .Z ( config1_decoder2.U151.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U151.ZN ) ,
    .I0 ( config1_decoder2.U151.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_61 ) ,
    .IN ( config1_decoder2.U151.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U96.AB ) ,
    .I0 ( config1_decoder2.n23 ) ,
    .I1 ( config1_decoder2.n31 ) ) ;
and ( 
    .Z ( config1_decoder2.U96.ZN ) ,
    .I0 ( config1_decoder2.U96.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_77 ) ,
    .IN ( config1_decoder2.U96.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.U1.BN ) ,
    .IN ( config1_decoder2.n19 ) ) ;
nand ( 
    .Z ( config1_decoder2.n16 ) ,
    .I0 ( config1_decoder2.U1.BN ) ,
    .I1 ( config1_decoder2.n20 ) ) ;
not ( 
    .O1 ( config1_decoder2.n36 ) ,
    .IN ( config1_decoder2.n17 ) ) ;
or ( 
    .Z ( config1_decoder2.U150.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n27 ) ) ;
and ( 
    .Z ( config1_decoder2.U150.ZN ) ,
    .I0 ( config1_decoder2.U150.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_8 ) ,
    .IN ( config1_decoder2.U150.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n52 ) ,
    .IN ( masks_hold_reg_2_2 ) ) ;
or ( 
    .Z ( config1_decoder2.U97.AB ) ,
    .I0 ( config1_decoder2.n23 ) ,
    .I1 ( config1_decoder2.n26 ) ) ;
and ( 
    .Z ( config1_decoder2.U97.ZN ) ,
    .I0 ( config1_decoder2.U97.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_89 ) ,
    .IN ( config1_decoder2.U97.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n18 ) ,
    .IN ( config1_decoder2.n37 ) ) ;
or ( 
    .Z ( config1_decoder2.U57.AB ) ,
    .I0 ( config1_decoder2.n26 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U57.ZN ) ,
    .I0 ( config1_decoder2.U57.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_26 ) ,
    .IN ( config1_decoder2.U57.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.U47.BN ) ,
    .IN ( config1_decoder2.n11 ) ) ;
nand ( 
    .Z ( config1_decoder2.n51 ) ,
    .I0 ( config1_decoder2.U47.BN ) ,
    .I1 ( config1_decoder2.n20 ) ) ;
or ( 
    .Z ( config1_decoder2.U77.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n42 ) ) ;
and ( 
    .Z ( config1_decoder2.U77.ZN ) ,
    .I0 ( config1_decoder2.U77.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_48 ) ,
    .IN ( config1_decoder2.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U67.AB ) ,
    .I0 ( config1_decoder2.n32 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U67.ZN ) ,
    .I0 ( config1_decoder2.U67.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_6 ) ,
    .IN ( config1_decoder2.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U10.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U10.ZN ) ,
    .I0 ( config1_decoder2.U10.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_18 ) ,
    .IN ( config1_decoder2.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n29 ) ,
    .I0 ( config1_decoder2.n48 ) ,
    .I1 ( config1_decoder2.n47 ) ) ;
or ( 
    .Z ( config1_decoder2.U26.AB ) ,
    .I0 ( config1_decoder2.n25 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U26.ZN ) ,
    .I0 ( config1_decoder2.U26.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_83 ) ,
    .IN ( config1_decoder2.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U113.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n24 ) ) ;
and ( 
    .Z ( config1_decoder2.U113.ZN ) ,
    .I0 ( config1_decoder2.U113.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_92 ) ,
    .IN ( config1_decoder2.U113.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U101.AB ) ,
    .I0 ( config1_decoder2.n22 ) ,
    .I1 ( config1_decoder2.n25 ) ) ;
and ( 
    .Z ( config1_decoder2.U101.ZN ) ,
    .I0 ( config1_decoder2.U101.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_91 ) ,
    .IN ( config1_decoder2.U101.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U138.AB ) ,
    .I0 ( config1_decoder2.n17 ) ,
    .I1 ( config1_decoder2.n16 ) ) ;
and ( 
    .Z ( config1_decoder2.U138.ZN ) ,
    .I0 ( config1_decoder2.U138.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_97 ) ,
    .IN ( config1_decoder2.U138.ZN ) ) ;
and ( 
    .Z ( config1_decoder2.n46 ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( masks_hold_reg_2_4 ) ) ;
nor ( 
    .Z ( config1_decoder2.n44 ) ,
    .I0 ( config1_decoder2.n45 ) ,
    .I1 ( masks_hold_reg_2_8 ) ) ;
and ( 
    .Z ( config1_decoder2.U125.AB ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( config1_decoder2.n35 ) ) ;
or ( 
    .Z ( config1_decoder2.n54 ) ,
    .I0 ( config1_decoder2.U125.AB ) ,
    .I1 ( config1_decoder2.n46 ) ,
    .I2 ( n79 ) ) ;
or ( 
    .Z ( config1_decoder2.U153.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n40 ) ) ;
and ( 
    .Z ( config1_decoder2.U153.ZN ) ,
    .I0 ( config1_decoder2.U153.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_42 ) ,
    .IN ( config1_decoder2.U153.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U141.AB ) ,
    .I0 ( config1_decoder2.n13 ) ,
    .I1 ( config1_decoder2.n14 ) ) ;
and ( 
    .Z ( config1_decoder2.U141.ZN ) ,
    .I0 ( config1_decoder2.U141.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_99 ) ,
    .IN ( config1_decoder2.U141.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U3.AB ) ,
    .I0 ( config1_decoder2.n27 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U3.ZN ) ,
    .I0 ( config1_decoder2.U3.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_16 ) ,
    .IN ( config1_decoder2.U3.ZN ) ) ;
not ( 
    .O1 ( config1_decoder2.n14 ) ,
    .IN ( config1_decoder2.n38 ) ) ;
or ( 
    .Z ( config1_decoder2.U58.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n33 ) ) ;
and ( 
    .Z ( config1_decoder2.U58.ZN ) ,
    .I0 ( config1_decoder2.U58.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_10 ) ,
    .IN ( config1_decoder2.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U46.AB ) ,
    .I0 ( config1_decoder2.n10 ) ,
    .I1 ( config1_decoder2.n32 ) ) ;
and ( 
    .Z ( config1_decoder2.U46.ZN ) ,
    .I0 ( config1_decoder2.U46.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_5 ) ,
    .IN ( config1_decoder2.U46.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U74.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n41 ) ) ;
and ( 
    .Z ( config1_decoder2.U74.ZN ) ,
    .I0 ( config1_decoder2.U74.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_53 ) ,
    .IN ( config1_decoder2.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U66.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U66.ZN ) ,
    .I0 ( config1_decoder2.U66.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_7 ) ,
    .IN ( config1_decoder2.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U11.AB ) ,
    .I0 ( config1_decoder2.n29 ) ,
    .I1 ( config1_decoder2.n30 ) ) ;
and ( 
    .Z ( config1_decoder2.U11.ZN ) ,
    .I0 ( config1_decoder2.U11.AB ) ,
    .I1 ( config1_decoder2.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_15 ) ,
    .IN ( config1_decoder2.U11.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n41 ) ,
    .I0 ( config1_decoder2.n44 ) ,
    .I1 ( config1_decoder2.n36 ) ) ;
nand ( 
    .Z ( config1_decoder2.n40 ) ,
    .I0 ( config1_decoder2.n44 ) ,
    .I1 ( config1_decoder2.n35 ) ) ;
or ( 
    .Z ( config1_decoder2.U25.AB ) ,
    .I0 ( config1_decoder2.n24 ) ,
    .I1 ( config1_decoder2.n28 ) ) ;
and ( 
    .Z ( config1_decoder2.U25.ZN ) ,
    .I0 ( config1_decoder2.U25.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_84 ) ,
    .IN ( config1_decoder2.U25.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U112.AB ) ,
    .I0 ( config1_decoder2.n24 ) ,
    .I1 ( config1_decoder2.n29 ) ) ;
and ( 
    .Z ( config1_decoder2.U112.ZN ) ,
    .I0 ( config1_decoder2.U112.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_80 ) ,
    .IN ( config1_decoder2.U112.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U102.AB ) ,
    .I0 ( config1_decoder2.n19 ) ,
    .I1 ( config1_decoder2.n23 ) ) ;
and ( 
    .Z ( config1_decoder2.U102.ZN ) ,
    .I0 ( config1_decoder2.U102.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_65 ) ,
    .IN ( config1_decoder2.U102.ZN ) ) ;
nand ( 
    .Z ( config1_decoder2.n17 ) ,
    .I0 ( masks_hold_reg_2_3 ) ,
    .I1 ( config1_decoder2.n52 ) ) ;
nor ( 
    .Z ( config1_decoder2.n38 ) ,
    .I0 ( masks_hold_reg_2_2 ) ,
    .I1 ( masks_hold_reg_2_3 ) ) ;
nand ( 
    .Z ( config1_decoder2.n32 ) ,
    .I0 ( config1_decoder2.n53 ) ,
    .I1 ( masks_hold_reg_2_4 ) ) ;
or ( 
    .Z ( config1_decoder2.U152.AB ) ,
    .I0 ( config1_decoder2.n11 ) ,
    .I1 ( config1_decoder2.n25 ) ) ;
and ( 
    .Z ( config1_decoder2.U152.ZN ) ,
    .I0 ( config1_decoder2.U152.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_71 ) ,
    .IN ( config1_decoder2.U152.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U142.AB ) ,
    .I0 ( config1_decoder2.n15 ) ,
    .I1 ( config1_decoder2.n16 ) ) ;
and ( 
    .Z ( config1_decoder2.U142.ZN ) ,
    .I0 ( config1_decoder2.U142.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_98 ) ,
    .IN ( config1_decoder2.U142.ZN ) ) ;
or ( 
    .Z ( config1_decoder2.U162.AB ) ,
    .I0 ( config1_decoder2.n28 ) ,
    .I1 ( config1_decoder2.n43 ) ) ;
and ( 
    .Z ( config1_decoder2.U162.ZN ) ,
    .I0 ( config1_decoder2.U162.AB ) ,
    .I1 ( config1_decoder2.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_1_51 ) ,
    .IN ( config1_decoder2.U162.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n99 ) ,
    .I0 ( masks_hold_reg_4_3 ) ,
    .I1 ( masks_hold_reg_4_4 ) ) ;
nand ( 
    .Z ( config1_decoder3.n97 ) ,
    .I0 ( masks_hold_reg_4_4 ) ,
    .I1 ( config1_decoder3.n62 ) ) ;
nor ( 
    .Z ( config1_decoder3.n94 ) ,
    .I0 ( config1_decoder3.n75 ) ,
    .I1 ( config1_decoder3.n69 ) ) ;
nor ( 
    .Z ( config1_decoder3.n80 ) ,
    .I0 ( config1_decoder3.n75 ) ,
    .I1 ( masks_hold_reg_4_8 ) ) ;
nor ( 
    .Z ( config1_decoder3.n76 ) ,
    .I0 ( masks_hold_reg_4_3 ) ,
    .I1 ( masks_hold_reg_4_4 ) ) ;
nand ( 
    .Z ( config1_decoder3.n1 ) ,
    .I0 ( config1_decoder3.n94 ) ,
    .I1 ( config1_decoder3.n60 ) ) ;
nand ( 
    .Z ( config1_decoder3.n85 ) ,
    .I0 ( config1_decoder3.n66 ) ,
    .I1 ( config1_decoder3.n67 ) ) ;
nand ( 
    .Z ( config1_decoder3.n95 ) ,
    .I0 ( config1_decoder3.n61 ) ,
    .I1 ( config1_decoder3.n67 ) ) ;
nand ( 
    .Z ( config1_decoder3.n71 ) ,
    .I0 ( config1_decoder3.n70 ) ,
    .I1 ( config1_decoder3.n76 ) ) ;
nand ( 
    .Z ( config1_decoder3.n86 ) ,
    .I0 ( config1_decoder3.n66 ) ,
    .I1 ( masks_hold_reg_4_5 ) ) ;
nand ( 
    .Z ( config1_decoder3.n72 ) ,
    .I0 ( config1_decoder3.n70 ) ,
    .I1 ( config1_decoder3.n77 ) ) ;
nand ( 
    .Z ( config1_decoder3.n74 ) ,
    .I0 ( config1_decoder3.n70 ) ,
    .I1 ( config1_decoder3.n79 ) ) ;
nand ( 
    .Z ( config1_decoder3.n73 ) ,
    .I0 ( config1_decoder3.n70 ) ,
    .I1 ( config1_decoder3.n78 ) ) ;
nand ( 
    .Z ( config1_decoder3.n82 ) ,
    .I0 ( config1_decoder3.n61 ) ,
    .I1 ( masks_hold_reg_4_5 ) ) ;
nand ( 
    .Z ( config1_decoder3.n83 ) ,
    .I0 ( config1_decoder3.n68 ) ,
    .I1 ( config1_decoder3.n65 ) ) ;
nand ( 
    .Z ( config1_decoder3.n103 ) ,
    .I0 ( config1_decoder3.n67 ) ,
    .I1 ( config1_decoder3.n65 ) ,
    .I2 ( masks_hold_reg_4_6 ) ) ;
nand ( 
    .Z ( config1_decoder3.n88 ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( config1_decoder3.n67 ) ,
    .I2 ( masks_hold_reg_4_7 ) ) ;
buf ( 
    .O1 ( config1_decoder3.n3 ) ,
    .IN ( config1_decoder3.n1 ) ) ;
not ( 
    .O1 ( config1_decoder3.n79 ) ,
    .IN ( config1_decoder3.n99 ) ) ;
not ( 
    .O1 ( config1_decoder3.n78 ) ,
    .IN ( config1_decoder3.n97 ) ) ;
buf ( 
    .O1 ( config1_decoder3.n2 ) ,
    .IN ( config1_decoder3.n1 ) ) ;
nor ( 
    .Z ( config1_decoder3.n77 ) ,
    .I0 ( config1_decoder3.n62 ) ,
    .I1 ( masks_hold_reg_4_4 ) ) ;
nand ( 
    .Z ( config1_decoder3.n92 ) ,
    .I0 ( masks_hold_reg_4_7 ) ,
    .I1 ( config1_decoder3.n68 ) ) ;
or ( 
    .Z ( config1_decoder3.U67.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U67.ZN ) ,
    .I0 ( config1_decoder3.U67.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_26 ) ,
    .IN ( config1_decoder3.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U10.AB ) ,
    .I0 ( config1_decoder3.n83 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U10.ZN ) ,
    .I0 ( config1_decoder3.U10.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_43 ) ,
    .IN ( config1_decoder3.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n90 ) ,
    .I0 ( config1_decoder3.n80 ) ,
    .I1 ( config1_decoder3.n77 ) ) ;
or ( 
    .Z ( config1_decoder3.U26.AB ) ,
    .I0 ( config1_decoder3.n91 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U26.ZN ) ,
    .I0 ( config1_decoder3.U26.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_81 ) ,
    .IN ( config1_decoder3.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U113.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n89 ) ) ;
and ( 
    .Z ( config1_decoder3.U113.ZN ) ,
    .I0 ( config1_decoder3.U113.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_91 ) ,
    .IN ( config1_decoder3.U113.ZN ) ) ;
nor ( 
    .Z ( config1_decoder3.n64 ) ,
    .I0 ( masks_hold_reg_4_8 ) ,
    .I1 ( n92 ) ) ;
nor ( 
    .Z ( config1_decoder3.n61 ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( masks_hold_reg_4_7 ) ) ;
or ( 
    .Z ( config1_decoder3.U128.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U128.ZN ) ,
    .I0 ( config1_decoder3.U128.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_62 ) ,
    .IN ( config1_decoder3.U128.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U125.AB ) ,
    .I0 ( config1_decoder3.n90 ) ,
    .I1 ( config1_decoder3.n88 ) ) ;
and ( 
    .Z ( config1_decoder3.U125.ZN ) ,
    .I0 ( config1_decoder3.U125.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_88 ) ,
    .IN ( config1_decoder3.U125.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U153.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U153.ZN ) ,
    .I0 ( config1_decoder3.U153.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_57 ) ,
    .IN ( config1_decoder3.U153.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.n65 ) ,
    .IN ( masks_hold_reg_4_7 ) ) ;
or ( 
    .Z ( config1_decoder3.U90.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n91 ) ) ;
and ( 
    .Z ( config1_decoder3.U90.ZN ) ,
    .I0 ( config1_decoder3.U90.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_73 ) ,
    .IN ( config1_decoder3.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U3.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U3.ZN ) ,
    .I0 ( config1_decoder3.U3.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_33 ) ,
    .IN ( config1_decoder3.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U13.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U13.ZN ) ,
    .I0 ( config1_decoder3.U13.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_15 ) ,
    .IN ( config1_decoder3.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n89 ) ,
    .I0 ( config1_decoder3.n80 ) ,
    .I1 ( config1_decoder3.n76 ) ) ;
or ( 
    .Z ( config1_decoder3.U28.AB ) ,
    .I0 ( config1_decoder3.n89 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U28.ZN ) ,
    .I0 ( config1_decoder3.U28.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_83 ) ,
    .IN ( config1_decoder3.U28.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U130.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n90 ) ) ;
and ( 
    .Z ( config1_decoder3.U130.ZN ) ,
    .I0 ( config1_decoder3.U130.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_72 ) ,
    .IN ( config1_decoder3.U130.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U120.AB ) ,
    .I0 ( config1_decoder3.n93 ) ,
    .I1 ( config1_decoder3.n88 ) ) ;
and ( 
    .Z ( config1_decoder3.U120.ZN ) ,
    .I0 ( config1_decoder3.U120.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_90 ) ,
    .IN ( config1_decoder3.U120.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U154.AB ) ,
    .I0 ( config1_decoder3.n96 ) ,
    .I1 ( config1_decoder3.n63 ) ) ;
and ( 
    .Z ( config1_decoder3.U154.ZN ) ,
    .I0 ( config1_decoder3.U154.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_104 ) ,
    .IN ( config1_decoder3.U154.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U160.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n91 ) ) ;
and ( 
    .Z ( config1_decoder3.U160.ZN ) ,
    .I0 ( config1_decoder3.U160.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_93 ) ,
    .IN ( config1_decoder3.U160.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U93.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U93.ZN ) ,
    .I0 ( config1_decoder3.U93.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_27 ) ,
    .IN ( config1_decoder3.U93.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U98.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n87 ) ) ;
and ( 
    .Z ( config1_decoder3.U98.ZN ) ,
    .I0 ( config1_decoder3.U98.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_4 ) ,
    .IN ( config1_decoder3.U98.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U83.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U83.ZN ) ,
    .I0 ( config1_decoder3.U83.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_53 ) ,
    .IN ( config1_decoder3.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U50.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n103 ) ) ;
and ( 
    .Z ( config1_decoder3.U50.ZN ) ,
    .I0 ( config1_decoder3.U50.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_9 ) ,
    .IN ( config1_decoder3.U50.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U30.AB ) ,
    .I0 ( config1_decoder3.n90 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U30.ZN ) ,
    .I0 ( config1_decoder3.U30.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_76 ) ,
    .IN ( config1_decoder3.U30.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U121.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n93 ) ) ;
and ( 
    .Z ( config1_decoder3.U121.ZN ) ,
    .I0 ( config1_decoder3.U121.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_74 ) ,
    .IN ( config1_decoder3.U121.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U157.AB ) ,
    .I0 ( config1_decoder3.n99 ) ,
    .I1 ( config1_decoder3.n98 ) ) ;
and ( 
    .Z ( config1_decoder3.U157.ZN ) ,
    .I0 ( config1_decoder3.U157.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_98 ) ,
    .IN ( config1_decoder3.U157.ZN ) ) ;
nor ( 
    .Z ( config1_decoder3.n70 ) ,
    .I0 ( config1_decoder3.n69 ) ,
    .I1 ( n92 ) ) ;
or ( 
    .Z ( config1_decoder3.U161.AB ) ,
    .I0 ( config1_decoder3.n100 ) ,
    .I1 ( config1_decoder3.n98 ) ) ;
and ( 
    .Z ( config1_decoder3.U161.ZN ) ,
    .I0 ( config1_decoder3.U161.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_95 ) ,
    .IN ( config1_decoder3.U161.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U82.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U82.ZN ) ,
    .I0 ( config1_decoder3.U82.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_59 ) ,
    .IN ( config1_decoder3.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U89.AB ) ,
    .I0 ( config1_decoder3.n99 ) ,
    .I1 ( config1_decoder3.n101 ) ) ;
and ( 
    .Z ( config1_decoder3.U89.ZN ) ,
    .I0 ( config1_decoder3.U89.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_102 ) ,
    .IN ( config1_decoder3.U89.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U51.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n82 ) ) ;
and ( 
    .Z ( config1_decoder3.U51.ZN ) ,
    .I0 ( config1_decoder3.U51.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_5 ) ,
    .IN ( config1_decoder3.U51.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U78.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U78.ZN ) ,
    .I0 ( config1_decoder3.U78.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_3 ) ,
    .IN ( config1_decoder3.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n104 ) ,
    .I0 ( config1_decoder3.n64 ) ,
    .I1 ( config1_decoder3.n78 ) ) ;
or ( 
    .Z ( config1_decoder3.U115.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n91 ) ) ;
and ( 
    .Z ( config1_decoder3.U115.ZN ) ,
    .I0 ( config1_decoder3.U115.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_65 ) ,
    .IN ( config1_decoder3.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U156.AB ) ,
    .I0 ( config1_decoder3.n97 ) ,
    .I1 ( config1_decoder3.n98 ) ) ;
and ( 
    .Z ( config1_decoder3.U156.ZN ) ,
    .I0 ( config1_decoder3.U156.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_97 ) ,
    .IN ( config1_decoder3.U156.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U5.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U5.ZN ) ,
    .I0 ( config1_decoder3.U5.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_34 ) ,
    .IN ( config1_decoder3.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U88.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U88.ZN ) ,
    .I0 ( config1_decoder3.U88.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_49 ) ,
    .IN ( config1_decoder3.U88.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.U52.BN ) ,
    .IN ( config1_decoder3.n103 ) ) ;
nand ( 
    .Z ( config1_decoder3.n63 ) ,
    .I0 ( config1_decoder3.U52.BN ) ,
    .I1 ( config1_decoder3.n94 ) ) ;
or ( 
    .Z ( config1_decoder3.U2.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U2.ZN ) ,
    .I0 ( config1_decoder3.U2.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_17 ) ,
    .IN ( config1_decoder3.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U81.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U81.ZN ) ,
    .I0 ( config1_decoder3.U81.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_60 ) ,
    .IN ( config1_decoder3.U81.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U59.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U59.ZN ) ,
    .I0 ( config1_decoder3.U59.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_37 ) ,
    .IN ( config1_decoder3.U59.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U49.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n92 ) ) ;
and ( 
    .Z ( config1_decoder3.U49.ZN ) ,
    .I0 ( config1_decoder3.U49.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_29 ) ,
    .IN ( config1_decoder3.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U75.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U75.ZN ) ,
    .I0 ( config1_decoder3.U75.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_7 ) ,
    .IN ( config1_decoder3.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U65.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U65.ZN ) ,
    .I0 ( config1_decoder3.U65.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_52 ) ,
    .IN ( config1_decoder3.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U12.AB ) ,
    .I0 ( config1_decoder3.n83 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U12.ZN ) ,
    .I0 ( config1_decoder3.U12.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_14 ) ,
    .IN ( config1_decoder3.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n93 ) ,
    .I0 ( config1_decoder3.n80 ) ,
    .I1 ( config1_decoder3.n79 ) ) ;
or ( 
    .Z ( config1_decoder3.U29.AB ) ,
    .I0 ( config1_decoder3.n89 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U29.ZN ) ,
    .I0 ( config1_decoder3.U29.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_75 ) ,
    .IN ( config1_decoder3.U29.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U123.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n90 ) ) ;
and ( 
    .Z ( config1_decoder3.U123.ZN ) ,
    .I0 ( config1_decoder3.U123.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_64 ) ,
    .IN ( config1_decoder3.U123.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U155.AB ) ,
    .I0 ( config1_decoder3.n101 ) ,
    .I1 ( config1_decoder3.n100 ) ) ;
and ( 
    .Z ( config1_decoder3.U155.ZN ) ,
    .I0 ( config1_decoder3.U155.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_99 ) ,
    .IN ( config1_decoder3.U155.ZN ) ) ;
nor ( 
    .Z ( config1_decoder3.n66 ) ,
    .I0 ( config1_decoder3.n65 ) ,
    .I1 ( masks_hold_reg_4_6 ) ) ;
or ( 
    .Z ( config1_decoder3.U163.AB ) ,
    .I0 ( config1_decoder3.n98 ) ,
    .I1 ( config1_decoder3.n96 ) ) ;
and ( 
    .Z ( config1_decoder3.U163.ZN ) ,
    .I0 ( config1_decoder3.U163.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_96 ) ,
    .IN ( config1_decoder3.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U80.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U80.ZN ) ,
    .I0 ( config1_decoder3.U80.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_58 ) ,
    .IN ( config1_decoder3.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U48.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n88 ) ) ;
and ( 
    .Z ( config1_decoder3.U48.ZN ) ,
    .I0 ( config1_decoder3.U48.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_25 ) ,
    .IN ( config1_decoder3.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U64.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U64.ZN ) ,
    .I0 ( config1_decoder3.U64.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_42 ) ,
    .IN ( config1_decoder3.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U79.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U79.ZN ) ,
    .I0 ( config1_decoder3.U79.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_2 ) ,
    .IN ( config1_decoder3.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U72.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U72.ZN ) ,
    .I0 ( config1_decoder3.U72.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_31 ) ,
    .IN ( config1_decoder3.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U69.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U69.ZN ) ,
    .I0 ( config1_decoder3.U69.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_10 ) ,
    .IN ( config1_decoder3.U69.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U119.AB ) ,
    .I0 ( config1_decoder3.n93 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U119.ZN ) ,
    .I0 ( config1_decoder3.U119.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_78 ) ,
    .IN ( config1_decoder3.U119.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U114.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U114.ZN ) ,
    .I0 ( config1_decoder3.U114.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_61 ) ,
    .IN ( config1_decoder3.U114.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U159.AB ) ,
    .I0 ( config1_decoder3.n101 ) ,
    .I1 ( config1_decoder3.n96 ) ) ;
and ( 
    .Z ( config1_decoder3.U159.ZN ) ,
    .I0 ( config1_decoder3.U159.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_100 ) ,
    .IN ( config1_decoder3.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U9.AB ) ,
    .I0 ( config1_decoder3.n83 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U9.ZN ) ,
    .I0 ( config1_decoder3.U9.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_44 ) ,
    .IN ( config1_decoder3.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U4.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U4.ZN ) ,
    .I0 ( config1_decoder3.U4.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_32 ) ,
    .IN ( config1_decoder3.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U53.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U53.ZN ) ,
    .I0 ( config1_decoder3.U53.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_21 ) ,
    .IN ( config1_decoder3.U53.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n84 ) ,
    .I0 ( config1_decoder3.n76 ) ,
    .I1 ( config1_decoder3.n64 ) ) ;
or ( 
    .Z ( config1_decoder3.U73.AB ) ,
    .I0 ( config1_decoder3.n87 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U73.ZN ) ,
    .I0 ( config1_decoder3.U73.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_16 ) ,
    .IN ( config1_decoder3.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U68.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U68.ZN ) ,
    .I0 ( config1_decoder3.U68.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_22 ) ,
    .IN ( config1_decoder3.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U63.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U63.ZN ) ,
    .I0 ( config1_decoder3.U63.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_40 ) ,
    .IN ( config1_decoder3.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U14.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U14.ZN ) ,
    .I0 ( config1_decoder3.U14.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_13 ) ,
    .IN ( config1_decoder3.U14.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U118.AB ) ,
    .I0 ( config1_decoder3.n93 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U118.ZN ) ,
    .I0 ( config1_decoder3.U118.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_86 ) ,
    .IN ( config1_decoder3.U118.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U117.AB ) ,
    .I0 ( config1_decoder3.n93 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U117.ZN ) ,
    .I0 ( config1_decoder3.U117.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_82 ) ,
    .IN ( config1_decoder3.U117.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U108.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n89 ) ) ;
and ( 
    .Z ( config1_decoder3.U108.ZN ) ,
    .I0 ( config1_decoder3.U108.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_67 ) ,
    .IN ( config1_decoder3.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U105.AB ) ,
    .I0 ( config1_decoder3.n91 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U105.ZN ) ,
    .I0 ( config1_decoder3.U105.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_85 ) ,
    .IN ( config1_decoder3.U105.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U158.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U158.ZN ) ,
    .I0 ( config1_decoder3.U158.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_54 ) ,
    .IN ( config1_decoder3.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U164.AB ) ,
    .I0 ( config1_decoder3.n97 ) ,
    .I1 ( config1_decoder3.n63 ) ) ;
and ( 
    .Z ( config1_decoder3.U164.ZN ) ,
    .I0 ( config1_decoder3.U164.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_105 ) ,
    .IN ( config1_decoder3.U164.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U94.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U94.ZN ) ,
    .I0 ( config1_decoder3.U94.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_19 ) ,
    .IN ( config1_decoder3.U94.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U8.AB ) ,
    .I0 ( config1_decoder3.n83 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U8.ZN ) ,
    .I0 ( config1_decoder3.U8.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_45 ) ,
    .IN ( config1_decoder3.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U7.AB ) ,
    .I0 ( config1_decoder3.n83 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U7.ZN ) ,
    .I0 ( config1_decoder3.U7.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_46 ) ,
    .IN ( config1_decoder3.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U54.AB ) ,
    .I0 ( config1_decoder3.n87 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U54.ZN ) ,
    .I0 ( config1_decoder3.U54.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_20 ) ,
    .IN ( config1_decoder3.U54.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n81 ) ,
    .I0 ( config1_decoder3.n79 ) ,
    .I1 ( config1_decoder3.n64 ) ) ;
or ( 
    .Z ( config1_decoder3.U70.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n87 ) ) ;
and ( 
    .Z ( config1_decoder3.U70.ZN ) ,
    .I0 ( config1_decoder3.U70.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_28 ) ,
    .IN ( config1_decoder3.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U62.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n73 ) ) ;
and ( 
    .Z ( config1_decoder3.U62.ZN ) ,
    .I0 ( config1_decoder3.U62.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_41 ) ,
    .IN ( config1_decoder3.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U15.AB ) ,
    .I0 ( config1_decoder3.n104 ) ,
    .I1 ( config1_decoder3.n95 ) ) ;
and ( 
    .Z ( config1_decoder3.U15.ZN ) ,
    .I0 ( config1_decoder3.U15.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_1 ) ,
    .IN ( config1_decoder3.U15.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U116.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n89 ) ) ;
and ( 
    .Z ( config1_decoder3.U116.ZN ) ,
    .I0 ( config1_decoder3.U116.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_71 ) ,
    .IN ( config1_decoder3.U116.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U109.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n89 ) ) ;
and ( 
    .Z ( config1_decoder3.U109.ZN ) ,
    .I0 ( config1_decoder3.U109.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_63 ) ,
    .IN ( config1_decoder3.U109.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U106.AB ) ,
    .I0 ( config1_decoder3.n91 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U106.ZN ) ,
    .I0 ( config1_decoder3.U106.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_77 ) ,
    .IN ( config1_decoder3.U106.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U126.AB ) ,
    .I0 ( config1_decoder3.n90 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U126.ZN ) ,
    .I0 ( config1_decoder3.U126.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_80 ) ,
    .IN ( config1_decoder3.U126.ZN ) ) ;
and ( 
    .Z ( config1_decoder3.n68 ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( masks_hold_reg_4_5 ) ) ;
or ( 
    .Z ( config1_decoder3.U165.AB ) ,
    .I0 ( config1_decoder3.n100 ) ,
    .I1 ( config1_decoder3.n63 ) ) ;
and ( 
    .Z ( config1_decoder3.U165.ZN ) ,
    .I0 ( config1_decoder3.U165.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_103 ) ,
    .IN ( config1_decoder3.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U6.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U6.ZN ) ,
    .I0 ( config1_decoder3.U6.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_47 ) ,
    .IN ( config1_decoder3.U6.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U85.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U85.ZN ) ,
    .I0 ( config1_decoder3.U85.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_55 ) ,
    .IN ( config1_decoder3.U85.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U55.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n87 ) ) ;
and ( 
    .Z ( config1_decoder3.U55.ZN ) ,
    .I0 ( config1_decoder3.U55.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_24 ) ,
    .IN ( config1_decoder3.U55.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U71.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U71.ZN ) ,
    .I0 ( config1_decoder3.U71.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_30 ) ,
    .IN ( config1_decoder3.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U61.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U61.ZN ) ,
    .I0 ( config1_decoder3.U61.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_38 ) ,
    .IN ( config1_decoder3.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U16.AB ) ,
    .I0 ( config1_decoder3.n87 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U16.ZN ) ,
    .I0 ( config1_decoder3.U16.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_12 ) ,
    .IN ( config1_decoder3.U16.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n87 ) ,
    .I0 ( config1_decoder3.n77 ) ,
    .I1 ( config1_decoder3.n64 ) ) ;
or ( 
    .Z ( config1_decoder3.U111.AB ) ,
    .I0 ( config1_decoder3.n89 ) ,
    .I1 ( config1_decoder3.n88 ) ) ;
and ( 
    .Z ( config1_decoder3.U111.ZN ) ,
    .I0 ( config1_decoder3.U111.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_87 ) ,
    .IN ( config1_decoder3.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U107.AB ) ,
    .I0 ( config1_decoder3.n91 ) ,
    .I1 ( config1_decoder3.n88 ) ) ;
and ( 
    .Z ( config1_decoder3.U107.ZN ) ,
    .I0 ( config1_decoder3.U107.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_89 ) ,
    .IN ( config1_decoder3.U107.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U127.AB ) ,
    .I0 ( config1_decoder3.n92 ) ,
    .I1 ( config1_decoder3.n90 ) ) ;
and ( 
    .Z ( config1_decoder3.U127.ZN ) ,
    .I0 ( config1_decoder3.U127.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_92 ) ,
    .IN ( config1_decoder3.U127.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.n75 ) ,
    .IN ( n92 ) ) ;
not ( 
    .O1 ( config1_decoder3.n100 ) ,
    .IN ( config1_decoder3.n76 ) ) ;
not ( 
    .O1 ( config1_decoder3.U1.BN ) ,
    .IN ( config1_decoder3.n95 ) ) ;
nand ( 
    .Z ( config1_decoder3.n98 ) ,
    .I0 ( config1_decoder3.U1.BN ) ,
    .I1 ( config1_decoder3.n94 ) ) ;
or ( 
    .Z ( config1_decoder3.U84.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U84.ZN ) ,
    .I0 ( config1_decoder3.U84.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_56 ) ,
    .IN ( config1_decoder3.U84.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U56.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n87 ) ) ;
and ( 
    .Z ( config1_decoder3.U56.ZN ) ,
    .I0 ( config1_decoder3.U56.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_8 ) ,
    .IN ( config1_decoder3.U56.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U76.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U76.ZN ) ,
    .I0 ( config1_decoder3.U76.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_6 ) ,
    .IN ( config1_decoder3.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U60.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U60.ZN ) ,
    .I0 ( config1_decoder3.U60.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_36 ) ,
    .IN ( config1_decoder3.U60.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U17.AB ) ,
    .I0 ( config1_decoder3.n84 ) ,
    .I1 ( config1_decoder3.n83 ) ) ;
and ( 
    .Z ( config1_decoder3.U17.ZN ) ,
    .I0 ( config1_decoder3.U17.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_11 ) ,
    .IN ( config1_decoder3.U17.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U27.AB ) ,
    .I0 ( config1_decoder3.n90 ) ,
    .I1 ( config1_decoder3.n86 ) ) ;
and ( 
    .Z ( config1_decoder3.U27.ZN ) ,
    .I0 ( config1_decoder3.U27.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_84 ) ,
    .IN ( config1_decoder3.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U110.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n91 ) ) ;
and ( 
    .Z ( config1_decoder3.U110.ZN ) ,
    .I0 ( config1_decoder3.U110.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_69 ) ,
    .IN ( config1_decoder3.U110.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.n67 ) ,
    .IN ( masks_hold_reg_4_5 ) ) ;
or ( 
    .Z ( config1_decoder3.U124.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n93 ) ) ;
and ( 
    .Z ( config1_decoder3.U124.ZN ) ,
    .I0 ( config1_decoder3.U124.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_70 ) ,
    .IN ( config1_decoder3.U124.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.n69 ) ,
    .IN ( masks_hold_reg_4_8 ) ) ;
and ( 
    .Z ( config1_decoder3.U140.AB ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( config1_decoder3.n79 ) ) ;
or ( 
    .Z ( config1_decoder3.n60 ) ,
    .I0 ( config1_decoder3.U140.AB ) ,
    .I1 ( config1_decoder3.n68 ) ,
    .I2 ( masks_hold_reg_4_7 ) ) ;
not ( 
    .O1 ( config1_decoder3.n96 ) ,
    .IN ( config1_decoder3.n77 ) ) ;
or ( 
    .Z ( config1_decoder3.U87.AB ) ,
    .I0 ( config1_decoder3.n97 ) ,
    .I1 ( config1_decoder3.n101 ) ) ;
and ( 
    .Z ( config1_decoder3.U87.ZN ) ,
    .I0 ( config1_decoder3.U87.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_101 ) ,
    .IN ( config1_decoder3.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U57.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U57.ZN ) ,
    .I0 ( config1_decoder3.U57.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_35 ) ,
    .IN ( config1_decoder3.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U77.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n87 ) ) ;
and ( 
    .Z ( config1_decoder3.U77.ZN ) ,
    .I0 ( config1_decoder3.U77.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_0 ) ,
    .IN ( config1_decoder3.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U86.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n72 ) ) ;
and ( 
    .Z ( config1_decoder3.U86.ZN ) ,
    .I0 ( config1_decoder3.U86.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_48 ) ,
    .IN ( config1_decoder3.U86.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U58.AB ) ,
    .I0 ( config1_decoder3.n103 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U58.ZN ) ,
    .I0 ( config1_decoder3.U58.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_39 ) ,
    .IN ( config1_decoder3.U58.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.U46.BN ) ,
    .IN ( config1_decoder3.n82 ) ) ;
nand ( 
    .Z ( config1_decoder3.n101 ) ,
    .I0 ( config1_decoder3.U46.BN ) ,
    .I1 ( config1_decoder3.n94 ) ) ;
or ( 
    .Z ( config1_decoder3.U74.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n81 ) ) ;
and ( 
    .Z ( config1_decoder3.U74.ZN ) ,
    .I0 ( config1_decoder3.U74.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_18 ) ,
    .IN ( config1_decoder3.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U66.AB ) ,
    .I0 ( config1_decoder3.n86 ) ,
    .I1 ( config1_decoder3.n71 ) ) ;
and ( 
    .Z ( config1_decoder3.U66.ZN ) ,
    .I0 ( config1_decoder3.U66.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_51 ) ,
    .IN ( config1_decoder3.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U11.AB ) ,
    .I0 ( config1_decoder3.n85 ) ,
    .I1 ( config1_decoder3.n74 ) ) ;
and ( 
    .Z ( config1_decoder3.U11.ZN ) ,
    .I0 ( config1_decoder3.U11.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_50 ) ,
    .IN ( config1_decoder3.U11.ZN ) ) ;
nand ( 
    .Z ( config1_decoder3.n91 ) ,
    .I0 ( config1_decoder3.n80 ) ,
    .I1 ( config1_decoder3.n78 ) ) ;
or ( 
    .Z ( config1_decoder3.U112.AB ) ,
    .I0 ( config1_decoder3.n89 ) ,
    .I1 ( config1_decoder3.n85 ) ) ;
and ( 
    .Z ( config1_decoder3.U112.ZN ) ,
    .I0 ( config1_decoder3.U112.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_79 ) ,
    .IN ( config1_decoder3.U112.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U129.AB ) ,
    .I0 ( config1_decoder3.n95 ) ,
    .I1 ( config1_decoder3.n93 ) ) ;
and ( 
    .Z ( config1_decoder3.U129.ZN ) ,
    .I0 ( config1_decoder3.U129.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_66 ) ,
    .IN ( config1_decoder3.U129.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U122.AB ) ,
    .I0 ( config1_decoder3.n82 ) ,
    .I1 ( config1_decoder3.n90 ) ) ;
and ( 
    .Z ( config1_decoder3.U122.ZN ) ,
    .I0 ( config1_decoder3.U122.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_68 ) ,
    .IN ( config1_decoder3.U122.ZN ) ) ;
not ( 
    .O1 ( config1_decoder3.n62 ) ,
    .IN ( masks_hold_reg_4_3 ) ) ;
or ( 
    .Z ( config1_decoder3.U162.AB ) ,
    .I0 ( config1_decoder3.n93 ) ,
    .I1 ( config1_decoder3.n92 ) ) ;
and ( 
    .Z ( config1_decoder3.U162.ZN ) ,
    .I0 ( config1_decoder3.U162.AB ) ,
    .I1 ( config1_decoder3.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_94 ) ,
    .IN ( config1_decoder3.U162.ZN ) ) ;
or ( 
    .Z ( config1_decoder3.U91.AB ) ,
    .I0 ( config1_decoder3.n88 ) ,
    .I1 ( config1_decoder3.n84 ) ) ;
and ( 
    .Z ( config1_decoder3.U91.ZN ) ,
    .I0 ( config1_decoder3.U91.AB ) ,
    .I1 ( config1_decoder3.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_2_23 ) ,
    .IN ( config1_decoder3.U91.ZN ) ) ;
and ( 
    .Z ( config1_decoder1.U199.AB ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config1_decoder1.U199.ZN ) ,
    .I0 ( config1_decoder1.U199.AB ) ,
    .I1 ( config1_decoder1.n1 ) ) ;
not ( 
    .O1 ( config1_decoder1.n2 ) ,
    .IN ( config1_decoder1.U199.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder1.n3 ) ,
    .IN ( config1_decoder1.n2 ) ) ;
buf ( 
    .O1 ( config1_decoder1.n4 ) ,
    .IN ( config1_decoder1.n2 ) ) ;
or ( 
    .Z ( config1_decoder1.U87.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n53 ) ) ;
and ( 
    .Z ( config1_decoder1.U87.ZN ) ,
    .I0 ( config1_decoder1.U87.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_138 ) ,
    .IN ( config1_decoder1.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U59.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n23 ) ) ;
and ( 
    .Z ( config1_decoder1.U59.ZN ) ,
    .I0 ( config1_decoder1.U59.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_66 ) ,
    .IN ( config1_decoder1.U59.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n23 ) ,
    .I0 ( config1_decoder1.n51 ) ,
    .I1 ( config1_decoder1.n36 ) ) ;
nand ( 
    .Z ( config1_decoder1.n25 ) ,
    .I0 ( config1_decoder1.n37 ) ,
    .I1 ( config1_decoder1.n39 ) ) ;
nor ( 
    .Z ( config1_decoder1.n35 ) ,
    .I0 ( masks_hold_reg_0_8 ) ,
    .I1 ( masks_hold_reg_0_9 ) ) ;
not ( 
    .O1 ( config1_decoder1.n63 ) ,
    .IN ( masks_hold_reg_0_5 ) ) ;
or ( 
    .Z ( config1_decoder1.U86.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n54 ) ) ;
and ( 
    .Z ( config1_decoder1.U86.ZN ) ,
    .I0 ( config1_decoder1.U86.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_137 ) ,
    .IN ( config1_decoder1.U86.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n14 ) ,
    .I0 ( config1_decoder1.n65 ) ,
    .I1 ( config1_decoder1.n36 ) ) ;
nand ( 
    .Z ( config1_decoder1.n31 ) ,
    .I0 ( config1_decoder1.n50 ) ,
    .I1 ( config1_decoder1.n64 ) ) ;
or ( 
    .Z ( config1_decoder1.U196.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U196.ZN ) ,
    .I0 ( config1_decoder1.U196.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_105 ) ,
    .IN ( config1_decoder1.U196.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.n58 ) ,
    .IN ( config1_decoder1.n44 ) ) ;
or ( 
    .Z ( config1_decoder1.U164.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U164.ZN ) ,
    .I0 ( config1_decoder1.U164.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_113 ) ,
    .IN ( config1_decoder1.U164.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U191.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U191.ZN ) ,
    .I0 ( config1_decoder1.U191.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_103 ) ,
    .IN ( config1_decoder1.U191.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U159.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n16 ) ) ;
and ( 
    .Z ( config1_decoder1.U159.ZN ) ,
    .I0 ( config1_decoder1.U159.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_96 ) ,
    .IN ( config1_decoder1.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U165.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U165.ZN ) ,
    .I0 ( config1_decoder1.U165.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_107 ) ,
    .IN ( config1_decoder1.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U190.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n42 ) ) ;
and ( 
    .Z ( config1_decoder1.U190.ZN ) ,
    .I0 ( config1_decoder1.U190.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_156 ) ,
    .IN ( config1_decoder1.U190.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U158.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n17 ) ) ;
and ( 
    .Z ( config1_decoder1.U158.ZN ) ,
    .I0 ( config1_decoder1.U158.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_95 ) ,
    .IN ( config1_decoder1.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U193.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n52 ) ) ;
and ( 
    .Z ( config1_decoder1.U193.ZN ) ,
    .I0 ( config1_decoder1.U193.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_147 ) ,
    .IN ( config1_decoder1.U193.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U192.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n49 ) ) ;
and ( 
    .Z ( config1_decoder1.U192.ZN ) ,
    .I0 ( config1_decoder1.U192.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_148 ) ,
    .IN ( config1_decoder1.U192.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U108.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U108.ZN ) ,
    .I0 ( config1_decoder1.U108.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_122 ) ,
    .IN ( config1_decoder1.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U168.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U168.ZN ) ,
    .I0 ( config1_decoder1.U168.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_58 ) ,
    .IN ( config1_decoder1.U168.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n27 ) ,
    .I0 ( config1_decoder1.n55 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config1_decoder1.U109.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U109.ZN ) ,
    .I0 ( config1_decoder1.U109.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_121 ) ,
    .IN ( config1_decoder1.U109.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U169.AB ) ,
    .I0 ( config1_decoder1.n30 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U169.ZN ) ,
    .I0 ( config1_decoder1.U169.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_61 ) ,
    .IN ( config1_decoder1.U169.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U239.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n49 ) ) ;
and ( 
    .Z ( config1_decoder1.U239.ZN ) ,
    .I0 ( config1_decoder1.U239.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_150 ) ,
    .IN ( config1_decoder1.U239.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U41.AB ) ,
    .I0 ( config1_decoder1.n23 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U41.ZN ) ,
    .I0 ( config1_decoder1.U41.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_18 ) ,
    .IN ( config1_decoder1.U41.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U40.AB ) ,
    .I0 ( config1_decoder1.n22 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U40.ZN ) ,
    .I0 ( config1_decoder1.U40.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_19 ) ,
    .IN ( config1_decoder1.U40.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U27.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U27.ZN ) ,
    .I0 ( config1_decoder1.U27.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_59 ) ,
    .IN ( config1_decoder1.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U43.AB ) ,
    .I0 ( config1_decoder1.n24 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U43.ZN ) ,
    .I0 ( config1_decoder1.U43.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_16 ) ,
    .IN ( config1_decoder1.U43.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U26.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n22 ) ) ;
and ( 
    .Z ( config1_decoder1.U26.ZN ) ,
    .I0 ( config1_decoder1.U26.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_11 ) ,
    .IN ( config1_decoder1.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U42.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U42.ZN ) ,
    .I0 ( config1_decoder1.U42.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_17 ) ,
    .IN ( config1_decoder1.U42.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U25.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U25.ZN ) ,
    .I0 ( config1_decoder1.U25.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_31 ) ,
    .IN ( config1_decoder1.U25.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U45.AB ) ,
    .I0 ( config1_decoder1.n31 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U45.ZN ) ,
    .I0 ( config1_decoder1.U45.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_53 ) ,
    .IN ( config1_decoder1.U45.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U24.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U24.ZN ) ,
    .I0 ( config1_decoder1.U24.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_1 ) ,
    .IN ( config1_decoder1.U24.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U44.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U44.ZN ) ,
    .I0 ( config1_decoder1.U44.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_51 ) ,
    .IN ( config1_decoder1.U44.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U23.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n10 ) ) ;
and ( 
    .Z ( config1_decoder1.U23.ZN ) ,
    .I0 ( config1_decoder1.U23.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_9 ) ,
    .IN ( config1_decoder1.U23.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U115.AB ) ,
    .I0 ( config1_decoder1.n22 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U115.ZN ) ,
    .I0 ( config1_decoder1.U115.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_83 ) ,
    .IN ( config1_decoder1.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U207.AB ) ,
    .I0 ( config1_decoder1.n21 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U207.ZN ) ,
    .I0 ( config1_decoder1.U207.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_76 ) ,
    .IN ( config1_decoder1.U207.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U47.AB ) ,
    .I0 ( config1_decoder1.n32 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U47.ZN ) ,
    .I0 ( config1_decoder1.U47.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_52 ) ,
    .IN ( config1_decoder1.U47.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n32 ) ,
    .I0 ( config1_decoder1.n65 ) ,
    .I1 ( config1_decoder1.n58 ) ) ;
or ( 
    .Z ( config1_decoder1.U114.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U114.ZN ) ,
    .I0 ( config1_decoder1.U114.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_86 ) ,
    .IN ( config1_decoder1.U114.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n10 ) ,
    .I0 ( config1_decoder1.n35 ) ,
    .I1 ( config1_decoder1.n55 ) ) ;
or ( 
    .Z ( config1_decoder1.U206.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U206.ZN ) ,
    .I0 ( config1_decoder1.U206.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_119 ) ,
    .IN ( config1_decoder1.U206.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U46.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U46.ZN ) ,
    .I0 ( config1_decoder1.U46.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_50 ) ,
    .IN ( config1_decoder1.U46.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n29 ) ,
    .I0 ( config1_decoder1.n50 ) ,
    .I1 ( config1_decoder1.n65 ) ) ;
or ( 
    .Z ( config1_decoder1.U117.AB ) ,
    .I0 ( config1_decoder1.n20 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U117.ZN ) ,
    .I0 ( config1_decoder1.U117.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_77 ) ,
    .IN ( config1_decoder1.U117.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n28 ) ,
    .I0 ( config1_decoder1.n35 ) ,
    .I1 ( config1_decoder1.n59 ) ) ;
or ( 
    .Z ( config1_decoder1.U173.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U173.ZN ) ,
    .I0 ( config1_decoder1.U173.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_56 ) ,
    .IN ( config1_decoder1.U173.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U205.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n54 ) ) ;
and ( 
    .Z ( config1_decoder1.U205.ZN ) ,
    .I0 ( config1_decoder1.U205.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_139 ) ,
    .IN ( config1_decoder1.U205.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U49.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n42 ) ) ;
and ( 
    .Z ( config1_decoder1.U49.ZN ) ,
    .I0 ( config1_decoder1.U49.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_152 ) ,
    .IN ( config1_decoder1.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U116.AB ) ,
    .I0 ( config1_decoder1.n22 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U116.ZN ) ,
    .I0 ( config1_decoder1.U116.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_75 ) ,
    .IN ( config1_decoder1.U116.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U172.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U172.ZN ) ,
    .I0 ( config1_decoder1.U172.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_57 ) ,
    .IN ( config1_decoder1.U172.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U204.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U204.ZN ) ,
    .I0 ( config1_decoder1.U204.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_112 ) ,
    .IN ( config1_decoder1.U204.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U230.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n14 ) ) ;
and ( 
    .Z ( config1_decoder1.U230.ZN ) ,
    .I0 ( config1_decoder1.U230.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_98 ) ,
    .IN ( config1_decoder1.U230.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U240.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n42 ) ) ;
and ( 
    .Z ( config1_decoder1.U240.ZN ) ,
    .I0 ( config1_decoder1.U240.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_158 ) ,
    .IN ( config1_decoder1.U240.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U90.AB ) ,
    .I0 ( config1_decoder1.n23 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U90.ZN ) ,
    .I0 ( config1_decoder1.U90.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_82 ) ,
    .IN ( config1_decoder1.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U78.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U78.ZN ) ,
    .I0 ( config1_decoder1.U78.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_47 ) ,
    .IN ( config1_decoder1.U78.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U195.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U195.ZN ) ,
    .I0 ( config1_decoder1.U195.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_104 ) ,
    .IN ( config1_decoder1.U195.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U101.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n56 ) ) ;
and ( 
    .Z ( config1_decoder1.U101.ZN ) ,
    .I0 ( config1_decoder1.U101.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_134 ) ,
    .IN ( config1_decoder1.U101.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n42 ) ,
    .I0 ( config1_decoder1.n47 ) ,
    .I1 ( config1_decoder1.n34 ) ) ;
or ( 
    .Z ( config1_decoder1.U161.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U161.ZN ) ,
    .I0 ( config1_decoder1.U161.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_100 ) ,
    .IN ( config1_decoder1.U161.ZN ) ) ;
and ( 
    .Z ( config1_decoder1.n60 ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( config1_decoder1.n62 ) ) ;
or ( 
    .Z ( config1_decoder1.U91.AB ) ,
    .I0 ( config1_decoder1.n21 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U91.ZN ) ,
    .I0 ( config1_decoder1.U91.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_84 ) ,
    .IN ( config1_decoder1.U91.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U79.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n17 ) ) ;
and ( 
    .Z ( config1_decoder1.U79.ZN ) ,
    .I0 ( config1_decoder1.U79.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_39 ) ,
    .IN ( config1_decoder1.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U194.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n52 ) ) ;
and ( 
    .Z ( config1_decoder1.U194.ZN ) ,
    .I0 ( config1_decoder1.U194.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_149 ) ,
    .IN ( config1_decoder1.U194.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U102.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n53 ) ) ;
and ( 
    .Z ( config1_decoder1.U102.ZN ) ,
    .I0 ( config1_decoder1.U102.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_140 ) ,
    .IN ( config1_decoder1.U102.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n43 ) ,
    .I0 ( config1_decoder1.n48 ) ,
    .I1 ( config1_decoder1.n34 ) ) ;
or ( 
    .Z ( config1_decoder1.U166.AB ) ,
    .I0 ( config1_decoder1.n27 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U166.ZN ) ,
    .I0 ( config1_decoder1.U166.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_110 ) ,
    .IN ( config1_decoder1.U166.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U232.AB ) ,
    .I0 ( config1_decoder1.n27 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U232.ZN ) ,
    .I0 ( config1_decoder1.U232.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_108 ) ,
    .IN ( config1_decoder1.U232.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U92.AB ) ,
    .I0 ( config1_decoder1.n20 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U92.ZN ) ,
    .I0 ( config1_decoder1.U92.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_85 ) ,
    .IN ( config1_decoder1.U92.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U197.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U197.ZN ) ,
    .I0 ( config1_decoder1.U197.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_94 ) ,
    .IN ( config1_decoder1.U197.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U103.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n54 ) ) ;
and ( 
    .Z ( config1_decoder1.U103.ZN ) ,
    .I0 ( config1_decoder1.U103.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_141 ) ,
    .IN ( config1_decoder1.U103.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.n50 ) ,
    .IN ( config1_decoder1.n41 ) ) ;
or ( 
    .Z ( config1_decoder1.U48.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n25 ) ) ;
and ( 
    .Z ( config1_decoder1.U48.ZN ) ,
    .I0 ( config1_decoder1.U48.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_7 ) ,
    .IN ( config1_decoder1.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U111.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U111.ZN ) ,
    .I0 ( config1_decoder1.U111.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_123 ) ,
    .IN ( config1_decoder1.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U171.AB ) ,
    .I0 ( config1_decoder1.n29 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U171.ZN ) ,
    .I0 ( config1_decoder1.U171.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_54 ) ,
    .IN ( config1_decoder1.U171.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.n61 ) ,
    .IN ( masks_hold_reg_0_2 ) ) ;
or ( 
    .Z ( config1_decoder1.U110.AB ) ,
    .I0 ( config1_decoder1.n23 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U110.ZN ) ,
    .I0 ( config1_decoder1.U110.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_74 ) ,
    .IN ( config1_decoder1.U110.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U170.AB ) ,
    .I0 ( config1_decoder1.n30 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U170.ZN ) ,
    .I0 ( config1_decoder1.U170.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_60 ) ,
    .IN ( config1_decoder1.U170.ZN ) ) ;
nor ( 
    .Z ( config1_decoder1.n39 ) ,
    .I0 ( masks_hold_reg_0_3 ) ,
    .I1 ( masks_hold_reg_0_4 ) ) ;
or ( 
    .Z ( config1_decoder1.U113.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U113.ZN ) ,
    .I0 ( config1_decoder1.U113.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_78 ) ,
    .IN ( config1_decoder1.U113.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U177.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n21 ) ) ;
and ( 
    .Z ( config1_decoder1.U177.ZN ) ,
    .I0 ( config1_decoder1.U177.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_12 ) ,
    .IN ( config1_decoder1.U177.ZN ) ) ;
nor ( 
    .Z ( config1_decoder1.n59 ) ,
    .I0 ( masks_hold_reg_0_5 ) ,
    .I1 ( masks_hold_reg_0_6 ) ) ;
or ( 
    .Z ( config1_decoder1.U112.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U112.ZN ) ,
    .I0 ( config1_decoder1.U112.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_115 ) ,
    .IN ( config1_decoder1.U112.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U176.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n23 ) ) ;
and ( 
    .Z ( config1_decoder1.U176.ZN ) ,
    .I0 ( config1_decoder1.U176.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_10 ) ,
    .IN ( config1_decoder1.U176.ZN ) ) ;
and ( 
    .Z ( config1_decoder1.U200.ABC ) ,
    .I0 ( config1_decoder1.n59 ) ,
    .I1 ( config1_decoder1.n61 ) ,
    .I2 ( config1_decoder1.n39 ) ) ;
or ( 
    .Z ( config1_decoder1.U200.ZN ) ,
    .I0 ( config1_decoder1.U200.ABC ) ,
    .I1 ( config1_decoder1.n40 ) ) ;
not ( 
    .O1 ( config1_decoder1.n1 ) ,
    .IN ( config1_decoder1.U200.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U175.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U175.ZN ) ,
    .I0 ( config1_decoder1.U175.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_48 ) ,
    .IN ( config1_decoder1.U175.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U174.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U174.ZN ) ,
    .I0 ( config1_decoder1.U174.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_49 ) ,
    .IN ( config1_decoder1.U174.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U29.AB ) ,
    .I0 ( config1_decoder1.n25 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U29.ZN ) ,
    .I0 ( config1_decoder1.U29.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_23 ) ,
    .IN ( config1_decoder1.U29.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U28.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U28.ZN ) ,
    .I0 ( config1_decoder1.U28.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_55 ) ,
    .IN ( config1_decoder1.U28.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U119.AB ) ,
    .I0 ( config1_decoder1.n25 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U119.ZN ) ,
    .I0 ( config1_decoder1.U119.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_71 ) ,
    .IN ( config1_decoder1.U119.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U179.AB ) ,
    .I0 ( config1_decoder1.n22 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U179.ZN ) ,
    .I0 ( config1_decoder1.U179.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_3 ) ,
    .IN ( config1_decoder1.U179.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U5.AB ) ,
    .I0 ( config1_decoder1.n28 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U5.ZN ) ,
    .I0 ( config1_decoder1.U5.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_37 ) ,
    .IN ( config1_decoder1.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U118.AB ) ,
    .I0 ( config1_decoder1.n25 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U118.ZN ) ,
    .I0 ( config1_decoder1.U118.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_79 ) ,
    .IN ( config1_decoder1.U118.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U178.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n20 ) ) ;
and ( 
    .Z ( config1_decoder1.U178.ZN ) ,
    .I0 ( config1_decoder1.U178.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_13 ) ,
    .IN ( config1_decoder1.U178.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U4.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U4.ZN ) ,
    .I0 ( config1_decoder1.U4.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_45 ) ,
    .IN ( config1_decoder1.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U209.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n56 ) ) ;
and ( 
    .Z ( config1_decoder1.U209.ZN ) ,
    .I0 ( config1_decoder1.U209.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_128 ) ,
    .IN ( config1_decoder1.U209.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U7.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n52 ) ) ;
and ( 
    .Z ( config1_decoder1.U7.ZN ) ,
    .I0 ( config1_decoder1.U7.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_143 ) ,
    .IN ( config1_decoder1.U7.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n9 ) ,
    .I0 ( config1_decoder1.n36 ) ,
    .I1 ( config1_decoder1.n37 ) ) ;
or ( 
    .Z ( config1_decoder1.U208.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n49 ) ) ;
and ( 
    .Z ( config1_decoder1.U208.ZN ) ,
    .I0 ( config1_decoder1.U208.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_144 ) ,
    .IN ( config1_decoder1.U208.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U6.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n53 ) ) ;
and ( 
    .Z ( config1_decoder1.U6.ZN ) ,
    .I0 ( config1_decoder1.U6.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_136 ) ,
    .IN ( config1_decoder1.U6.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n16 ) ,
    .I0 ( config1_decoder1.n65 ) ,
    .I1 ( config1_decoder1.n39 ) ) ;
or ( 
    .Z ( config1_decoder1.U1.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U1.ZN ) ,
    .I0 ( config1_decoder1.U1.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_35 ) ,
    .IN ( config1_decoder1.U1.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U3.AB ) ,
    .I0 ( config1_decoder1.n29 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U3.ZN ) ,
    .I0 ( config1_decoder1.U3.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_62 ) ,
    .IN ( config1_decoder1.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U2.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n15 ) ) ;
and ( 
    .Z ( config1_decoder1.U2.ZN ) ,
    .I0 ( config1_decoder1.U2.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_41 ) ,
    .IN ( config1_decoder1.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U9.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n52 ) ) ;
and ( 
    .Z ( config1_decoder1.U9.ZN ) ,
    .I0 ( config1_decoder1.U9.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_145 ) ,
    .IN ( config1_decoder1.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U8.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n49 ) ) ;
and ( 
    .Z ( config1_decoder1.U8.ZN ) ,
    .I0 ( config1_decoder1.U8.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_146 ) ,
    .IN ( config1_decoder1.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U50.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n43 ) ) ;
and ( 
    .Z ( config1_decoder1.U50.ZN ) ,
    .I0 ( config1_decoder1.U50.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_151 ) ,
    .IN ( config1_decoder1.U50.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U51.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n43 ) ) ;
and ( 
    .Z ( config1_decoder1.U51.ZN ) ,
    .I0 ( config1_decoder1.U51.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_153 ) ,
    .IN ( config1_decoder1.U51.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U63.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n22 ) ) ;
and ( 
    .Z ( config1_decoder1.U63.ZN ) ,
    .I0 ( config1_decoder1.U63.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_91 ) ,
    .IN ( config1_decoder1.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U36.AB ) ,
    .I0 ( config1_decoder1.n24 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U36.ZN ) ,
    .I0 ( config1_decoder1.U36.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_24 ) ,
    .IN ( config1_decoder1.U36.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U62.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n20 ) ) ;
and ( 
    .Z ( config1_decoder1.U62.ZN ) ,
    .I0 ( config1_decoder1.U62.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_93 ) ,
    .IN ( config1_decoder1.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U37.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U37.ZN ) ,
    .I0 ( config1_decoder1.U37.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_22 ) ,
    .IN ( config1_decoder1.U37.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U89.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n56 ) ) ;
and ( 
    .Z ( config1_decoder1.U89.ZN ) ,
    .I0 ( config1_decoder1.U89.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_130 ) ,
    .IN ( config1_decoder1.U89.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U61.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n21 ) ) ;
and ( 
    .Z ( config1_decoder1.U61.ZN ) ,
    .I0 ( config1_decoder1.U61.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_68 ) ,
    .IN ( config1_decoder1.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U34.AB ) ,
    .I0 ( config1_decoder1.n23 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U34.ZN ) ,
    .I0 ( config1_decoder1.U34.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_26 ) ,
    .IN ( config1_decoder1.U34.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U88.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n57 ) ) ;
and ( 
    .Z ( config1_decoder1.U88.ZN ) ,
    .I0 ( config1_decoder1.U88.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_129 ) ,
    .IN ( config1_decoder1.U88.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U60.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n21 ) ) ;
and ( 
    .Z ( config1_decoder1.U60.ZN ) ,
    .I0 ( config1_decoder1.U60.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_92 ) ,
    .IN ( config1_decoder1.U60.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U35.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U35.ZN ) ,
    .I0 ( config1_decoder1.U35.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_25 ) ,
    .IN ( config1_decoder1.U35.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U55.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n13 ) ) ;
and ( 
    .Z ( config1_decoder1.U55.ZN ) ,
    .I0 ( config1_decoder1.U55.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_65 ) ,
    .IN ( config1_decoder1.U55.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U67.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U67.ZN ) ,
    .I0 ( config1_decoder1.U67.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_126 ) ,
    .IN ( config1_decoder1.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U32.AB ) ,
    .I0 ( config1_decoder1.n21 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U32.ZN ) ,
    .I0 ( config1_decoder1.U32.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_28 ) ,
    .IN ( config1_decoder1.U32.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n13 ) ,
    .I0 ( masks_hold_reg_0_8 ) ,
    .I1 ( config1_decoder1.n59 ) ) ;
or ( 
    .Z ( config1_decoder1.U56.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n24 ) ) ;
and ( 
    .Z ( config1_decoder1.U56.ZN ) ,
    .I0 ( config1_decoder1.U56.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_88 ) ,
    .IN ( config1_decoder1.U56.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U66.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n25 ) ) ;
and ( 
    .Z ( config1_decoder1.U66.ZN ) ,
    .I0 ( config1_decoder1.U66.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_63 ) ,
    .IN ( config1_decoder1.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U33.AB ) ,
    .I0 ( config1_decoder1.n22 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U33.ZN ) ,
    .I0 ( config1_decoder1.U33.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_27 ) ,
    .IN ( config1_decoder1.U33.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n18 ) ,
    .I0 ( config1_decoder1.n50 ) ,
    .I1 ( config1_decoder1.n51 ) ) ;
nand ( 
    .Z ( config1_decoder1.n41 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( masks_hold_reg_0_3 ) ) ;
nand ( 
    .Z ( config1_decoder1.n26 ) ,
    .I0 ( config1_decoder1.n38 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config1_decoder1.U85.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n54 ) ) ;
and ( 
    .Z ( config1_decoder1.U85.ZN ) ,
    .I0 ( config1_decoder1.U85.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_135 ) ,
    .IN ( config1_decoder1.U85.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U57.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n24 ) ) ;
and ( 
    .Z ( config1_decoder1.U57.ZN ) ,
    .I0 ( config1_decoder1.U57.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_64 ) ,
    .IN ( config1_decoder1.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U65.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n25 ) ) ;
and ( 
    .Z ( config1_decoder1.U65.ZN ) ,
    .I0 ( config1_decoder1.U65.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_87 ) ,
    .IN ( config1_decoder1.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U30.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U30.ZN ) ,
    .I0 ( config1_decoder1.U30.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_30 ) ,
    .IN ( config1_decoder1.U30.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U188.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n43 ) ) ;
and ( 
    .Z ( config1_decoder1.U188.ZN ) ,
    .I0 ( config1_decoder1.U188.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_155 ) ,
    .IN ( config1_decoder1.U188.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n21 ) ,
    .I0 ( config1_decoder1.n51 ) ,
    .I1 ( config1_decoder1.n58 ) ) ;
nand ( 
    .Z ( config1_decoder1.n30 ) ,
    .I0 ( config1_decoder1.n34 ) ,
    .I1 ( config1_decoder1.n35 ) ) ;
nor ( 
    .Z ( config1_decoder1.n36 ) ,
    .I0 ( config1_decoder1.n66 ) ,
    .I1 ( masks_hold_reg_0_4 ) ) ;
or ( 
    .Z ( config1_decoder1.U84.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U84.ZN ) ,
    .I0 ( config1_decoder1.U84.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_34 ) ,
    .IN ( config1_decoder1.U84.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U58.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n23 ) ) ;
and ( 
    .Z ( config1_decoder1.U58.ZN ) ,
    .I0 ( config1_decoder1.U58.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_90 ) ,
    .IN ( config1_decoder1.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U64.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n22 ) ) ;
and ( 
    .Z ( config1_decoder1.U64.ZN ) ,
    .I0 ( config1_decoder1.U64.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_67 ) ,
    .IN ( config1_decoder1.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U31.AB ) ,
    .I0 ( config1_decoder1.n20 ) ,
    .I1 ( config1_decoder1.n30 ) ) ;
and ( 
    .Z ( config1_decoder1.U31.ZN ) ,
    .I0 ( config1_decoder1.U31.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_29 ) ,
    .IN ( config1_decoder1.U31.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U189.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U189.ZN ) ,
    .I0 ( config1_decoder1.U189.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_102 ) ,
    .IN ( config1_decoder1.U189.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n12 ) ,
    .I0 ( config1_decoder1.n58 ) ,
    .I1 ( config1_decoder1.n64 ) ) ;
nand ( 
    .Z ( config1_decoder1.n33 ) ,
    .I0 ( config1_decoder1.n38 ) ,
    .I1 ( config1_decoder1.n35 ) ) ;
nor ( 
    .Z ( config1_decoder1.n55 ) ,
    .I0 ( config1_decoder1.n63 ) ,
    .I1 ( masks_hold_reg_0_6 ) ) ;
not ( 
    .O1 ( config1_decoder1.n66 ) ,
    .IN ( masks_hold_reg_0_3 ) ) ;
or ( 
    .Z ( config1_decoder1.U167.AB ) ,
    .I0 ( config1_decoder1.n27 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U167.ZN ) ,
    .I0 ( config1_decoder1.U167.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_109 ) ,
    .IN ( config1_decoder1.U167.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U233.AB ) ,
    .I0 ( config1_decoder1.n12 ) ,
    .I1 ( config1_decoder1.n13 ) ) ;
and ( 
    .Z ( config1_decoder1.U233.ZN ) ,
    .I0 ( config1_decoder1.U233.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_99 ) ,
    .IN ( config1_decoder1.U233.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U93.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n18 ) ) ;
and ( 
    .Z ( config1_decoder1.U93.ZN ) ,
    .I0 ( config1_decoder1.U93.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_70 ) ,
    .IN ( config1_decoder1.U93.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.U213.BN ) ,
    .IN ( masks_hold_reg_0_6 ) ) ;
nor ( 
    .Z ( config1_decoder1.n38 ) ,
    .I0 ( config1_decoder1.U213.BN ) ,
    .I1 ( masks_hold_reg_0_5 ) ) ;
nor ( 
    .Z ( config1_decoder1.n51 ) ,
    .I0 ( config1_decoder1.n61 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
or ( 
    .Z ( config1_decoder1.U81.AB ) ,
    .I0 ( config1_decoder1.n28 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U81.ZN ) ,
    .I0 ( config1_decoder1.U81.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_38 ) ,
    .IN ( config1_decoder1.U81.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U69.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U69.ZN ) ,
    .I0 ( config1_decoder1.U69.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_124 ) ,
    .IN ( config1_decoder1.U69.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U184.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n18 ) ) ;
and ( 
    .Z ( config1_decoder1.U184.ZN ) ,
    .I0 ( config1_decoder1.U184.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_14 ) ,
    .IN ( config1_decoder1.U184.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n15 ) ,
    .I0 ( config1_decoder1.n64 ) ,
    .I1 ( config1_decoder1.n36 ) ) ;
not ( 
    .O1 ( config1_decoder1.n46 ) ,
    .IN ( config1_decoder1.n39 ) ) ;
or ( 
    .Z ( config1_decoder1.U210.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n20 ) ) ;
and ( 
    .Z ( config1_decoder1.U210.ZN ) ,
    .I0 ( config1_decoder1.U210.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_69 ) ,
    .IN ( config1_decoder1.U210.ZN ) ) ;
nor ( 
    .Z ( config1_decoder1.n37 ) ,
    .I0 ( masks_hold_reg_0_2 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
or ( 
    .Z ( config1_decoder1.U80.AB ) ,
    .I0 ( config1_decoder1.n28 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U80.ZN ) ,
    .I0 ( config1_decoder1.U80.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_36 ) ,
    .IN ( config1_decoder1.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U68.AB ) ,
    .I0 ( config1_decoder1.n26 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U68.ZN ) ,
    .I0 ( config1_decoder1.U68.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_118 ) ,
    .IN ( config1_decoder1.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U185.AB ) ,
    .I0 ( config1_decoder1.n20 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U185.ZN ) ,
    .I0 ( config1_decoder1.U185.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_5 ) ,
    .IN ( config1_decoder1.U185.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n24 ) ,
    .I0 ( config1_decoder1.n51 ) ,
    .I1 ( config1_decoder1.n39 ) ) ;
not ( 
    .O1 ( config1_decoder1.n45 ) ,
    .IN ( config1_decoder1.n36 ) ) ;
or ( 
    .Z ( config1_decoder1.U211.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n53 ) ) ;
and ( 
    .Z ( config1_decoder1.U211.ZN ) ,
    .I0 ( config1_decoder1.U211.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_142 ) ,
    .IN ( config1_decoder1.U211.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.U223.BN ) ,
    .IN ( config1_decoder1.n60 ) ) ;
nor ( 
    .Z ( config1_decoder1.n48 ) ,
    .I0 ( config1_decoder1.U223.BN ) ,
    .I1 ( masks_hold_reg_0_2 ) ) ;
or ( 
    .Z ( config1_decoder1.U83.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U83.ZN ) ,
    .I0 ( config1_decoder1.U83.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_32 ) ,
    .IN ( config1_decoder1.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U186.AB ) ,
    .I0 ( config1_decoder1.n21 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U186.ZN ) ,
    .I0 ( config1_decoder1.U186.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_4 ) ,
    .IN ( config1_decoder1.U186.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n17 ) ,
    .I0 ( config1_decoder1.n64 ) ,
    .I1 ( config1_decoder1.n39 ) ) ;
nand ( 
    .Z ( config1_decoder1.n57 ) ,
    .I0 ( config1_decoder1.n48 ) ,
    .I1 ( config1_decoder1.n59 ) ) ;
nor ( 
    .Z ( config1_decoder1.n64 ) ,
    .I0 ( config1_decoder1.n62 ) ,
    .I1 ( masks_hold_reg_0_2 ) ) ;
or ( 
    .Z ( config1_decoder1.U82.AB ) ,
    .I0 ( config1_decoder1.n15 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U82.ZN ) ,
    .I0 ( config1_decoder1.U82.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_33 ) ,
    .IN ( config1_decoder1.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U187.AB ) ,
    .I0 ( config1_decoder1.n18 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U187.ZN ) ,
    .I0 ( config1_decoder1.U187.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_6 ) ,
    .IN ( config1_decoder1.U187.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n56 ) ,
    .I0 ( config1_decoder1.n47 ) ,
    .I1 ( config1_decoder1.n59 ) ) ;
or ( 
    .Z ( config1_decoder1.U38.AB ) ,
    .I0 ( config1_decoder1.n20 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U38.ZN ) ,
    .I0 ( config1_decoder1.U38.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_21 ) ,
    .IN ( config1_decoder1.U38.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U180.AB ) ,
    .I0 ( config1_decoder1.n24 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U180.ZN ) ,
    .I0 ( config1_decoder1.U180.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_0 ) ,
    .IN ( config1_decoder1.U180.ZN ) ) ;
nor ( 
    .Z ( config1_decoder1.n65 ) ,
    .I0 ( config1_decoder1.n61 ) ,
    .I1 ( config1_decoder1.n62 ) ) ;
or ( 
    .Z ( config1_decoder1.U39.AB ) ,
    .I0 ( config1_decoder1.n21 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U39.ZN ) ,
    .I0 ( config1_decoder1.U39.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_20 ) ,
    .IN ( config1_decoder1.U39.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U181.AB ) ,
    .I0 ( config1_decoder1.n23 ) ,
    .I1 ( config1_decoder1.n28 ) ) ;
and ( 
    .Z ( config1_decoder1.U181.ZN ) ,
    .I0 ( config1_decoder1.U181.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_2 ) ,
    .IN ( config1_decoder1.U181.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.U149.BN ) ,
    .IN ( config1_decoder1.n60 ) ) ;
nor ( 
    .Z ( config1_decoder1.n47 ) ,
    .I0 ( config1_decoder1.U149.BN ) ,
    .I1 ( config1_decoder1.n61 ) ) ;
or ( 
    .Z ( config1_decoder1.U182.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n24 ) ) ;
and ( 
    .Z ( config1_decoder1.U182.ZN ) ,
    .I0 ( config1_decoder1.U182.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_8 ) ,
    .IN ( config1_decoder1.U182.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U183.AB ) ,
    .I0 ( config1_decoder1.n25 ) ,
    .I1 ( config1_decoder1.n33 ) ) ;
and ( 
    .Z ( config1_decoder1.U183.ZN ) ,
    .I0 ( config1_decoder1.U183.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_15 ) ,
    .IN ( config1_decoder1.U183.ZN ) ) ;
not ( 
    .O1 ( config1_decoder1.n62 ) ,
    .IN ( masks_hold_reg_0_7 ) ) ;
nand ( 
    .Z ( config1_decoder1.n44 ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( config1_decoder1.n66 ) ) ;
nand ( 
    .Z ( config1_decoder1.n40 ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( masks_hold_reg_0_7 ) ) ;
nand ( 
    .Z ( config1_decoder1.n20 ) ,
    .I0 ( config1_decoder1.n50 ) ,
    .I1 ( config1_decoder1.n37 ) ) ;
not ( 
    .O1 ( config1_decoder1.U219.BN ) ,
    .IN ( masks_hold_reg_0_6 ) ) ;
nor ( 
    .Z ( config1_decoder1.n34 ) ,
    .I0 ( config1_decoder1.U219.BN ) ,
    .I1 ( config1_decoder1.n63 ) ) ;
nand ( 
    .Z ( config1_decoder1.n22 ) ,
    .I0 ( config1_decoder1.n58 ) ,
    .I1 ( config1_decoder1.n37 ) ) ;
or ( 
    .Z ( config1_decoder1.U72.AB ) ,
    .I0 ( config1_decoder1.n26 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U72.ZN ) ,
    .I0 ( config1_decoder1.U72.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_117 ) ,
    .IN ( config1_decoder1.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U73.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n16 ) ) ;
and ( 
    .Z ( config1_decoder1.U73.ZN ) ,
    .I0 ( config1_decoder1.U73.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_40 ) ,
    .IN ( config1_decoder1.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U98.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n56 ) ) ;
and ( 
    .Z ( config1_decoder1.U98.ZN ) ,
    .I0 ( config1_decoder1.U98.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_132 ) ,
    .IN ( config1_decoder1.U98.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U70.AB ) ,
    .I0 ( config1_decoder1.n26 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U70.ZN ) ,
    .I0 ( config1_decoder1.U70.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_116 ) ,
    .IN ( config1_decoder1.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U99.AB ) ,
    .I0 ( config1_decoder1.n44 ) ,
    .I1 ( config1_decoder1.n57 ) ) ;
and ( 
    .Z ( config1_decoder1.U99.ZN ) ,
    .I0 ( config1_decoder1.U99.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_131 ) ,
    .IN ( config1_decoder1.U99.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U71.AB ) ,
    .I0 ( config1_decoder1.n19 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U71.ZN ) ,
    .I0 ( config1_decoder1.U71.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_125 ) ,
    .IN ( config1_decoder1.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U76.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n32 ) ) ;
and ( 
    .Z ( config1_decoder1.U76.ZN ) ,
    .I0 ( config1_decoder1.U76.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_44 ) ,
    .IN ( config1_decoder1.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U77.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n29 ) ) ;
and ( 
    .Z ( config1_decoder1.U77.ZN ) ,
    .I0 ( config1_decoder1.U77.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_46 ) ,
    .IN ( config1_decoder1.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U104.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U104.ZN ) ,
    .I0 ( config1_decoder1.U104.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_81 ) ,
    .IN ( config1_decoder1.U104.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U94.AB ) ,
    .I0 ( config1_decoder1.n24 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U94.ZN ) ,
    .I0 ( config1_decoder1.U94.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_72 ) ,
    .IN ( config1_decoder1.U94.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U74.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n14 ) ) ;
and ( 
    .Z ( config1_decoder1.U74.ZN ) ,
    .I0 ( config1_decoder1.U74.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_42 ) ,
    .IN ( config1_decoder1.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U105.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U105.ZN ) ,
    .I0 ( config1_decoder1.U105.AB ) ,
    .I1 ( config1_decoder1.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_89 ) ,
    .IN ( config1_decoder1.U105.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n49 ) ,
    .I0 ( config1_decoder1.n47 ) ,
    .I1 ( config1_decoder1.n38 ) ) ;
nand ( 
    .Z ( config1_decoder1.n19 ) ,
    .I0 ( config1_decoder1.n34 ) ,
    .I1 ( masks_hold_reg_0_8 ) ) ;
or ( 
    .Z ( config1_decoder1.U243.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n43 ) ) ;
and ( 
    .Z ( config1_decoder1.U243.ZN ) ,
    .I0 ( config1_decoder1.U243.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_157 ) ,
    .IN ( config1_decoder1.U243.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U95.AB ) ,
    .I0 ( config1_decoder1.n9 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U95.ZN ) ,
    .I0 ( config1_decoder1.U95.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_73 ) ,
    .IN ( config1_decoder1.U95.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U75.AB ) ,
    .I0 ( config1_decoder1.n10 ) ,
    .I1 ( config1_decoder1.n12 ) ) ;
and ( 
    .Z ( config1_decoder1.U75.ZN ) ,
    .I0 ( config1_decoder1.U75.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_43 ) ,
    .IN ( config1_decoder1.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U106.AB ) ,
    .I0 ( config1_decoder1.n16 ) ,
    .I1 ( config1_decoder1.n19 ) ) ;
and ( 
    .Z ( config1_decoder1.U106.ZN ) ,
    .I0 ( config1_decoder1.U106.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_120 ) ,
    .IN ( config1_decoder1.U106.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n52 ) ,
    .I0 ( config1_decoder1.n48 ) ,
    .I1 ( config1_decoder1.n38 ) ) ;
or ( 
    .Z ( config1_decoder1.U162.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n31 ) ) ;
and ( 
    .Z ( config1_decoder1.U162.ZN ) ,
    .I0 ( config1_decoder1.U162.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_101 ) ,
    .IN ( config1_decoder1.U162.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U236.AB ) ,
    .I0 ( config1_decoder1.n45 ) ,
    .I1 ( config1_decoder1.n42 ) ) ;
and ( 
    .Z ( config1_decoder1.U236.ZN ) ,
    .I0 ( config1_decoder1.U236.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_154 ) ,
    .IN ( config1_decoder1.U236.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U242.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n27 ) ) ;
and ( 
    .Z ( config1_decoder1.U242.ZN ) ,
    .I0 ( config1_decoder1.U242.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_106 ) ,
    .IN ( config1_decoder1.U242.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U96.AB ) ,
    .I0 ( config1_decoder1.n17 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U96.ZN ) ,
    .I0 ( config1_decoder1.U96.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_111 ) ,
    .IN ( config1_decoder1.U96.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U107.AB ) ,
    .I0 ( config1_decoder1.n24 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U107.ZN ) ,
    .I0 ( config1_decoder1.U107.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_80 ) ,
    .IN ( config1_decoder1.U107.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n54 ) ,
    .I0 ( config1_decoder1.n48 ) ,
    .I1 ( config1_decoder1.n55 ) ) ;
or ( 
    .Z ( config1_decoder1.U163.AB ) ,
    .I0 ( config1_decoder1.n14 ) ,
    .I1 ( config1_decoder1.n26 ) ) ;
and ( 
    .Z ( config1_decoder1.U163.ZN ) ,
    .I0 ( config1_decoder1.U163.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_114 ) ,
    .IN ( config1_decoder1.U163.ZN ) ) ;
nand ( 
    .Z ( config1_onehot_decoded_masks_0_159 ) ,
    .I0 ( config1_decoder1.n2 ) ,
    .I1 ( config1_decoder1.n40 ) ) ;
or ( 
    .Z ( config1_decoder1.U97.AB ) ,
    .I0 ( config1_decoder1.n46 ) ,
    .I1 ( config1_decoder1.n57 ) ) ;
and ( 
    .Z ( config1_decoder1.U97.ZN ) ,
    .I0 ( config1_decoder1.U97.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_127 ) ,
    .IN ( config1_decoder1.U97.ZN ) ) ;
or ( 
    .Z ( config1_decoder1.U100.AB ) ,
    .I0 ( config1_decoder1.n41 ) ,
    .I1 ( config1_decoder1.n57 ) ) ;
and ( 
    .Z ( config1_decoder1.U100.ZN ) ,
    .I0 ( config1_decoder1.U100.AB ) ,
    .I1 ( config1_decoder1.n3 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_133 ) ,
    .IN ( config1_decoder1.U100.ZN ) ) ;
nand ( 
    .Z ( config1_decoder1.n53 ) ,
    .I0 ( config1_decoder1.n47 ) ,
    .I1 ( config1_decoder1.n55 ) ) ;
or ( 
    .Z ( config1_decoder1.U160.AB ) ,
    .I0 ( config1_decoder1.n13 ) ,
    .I1 ( config1_decoder1.n15 ) ) ;
and ( 
    .Z ( config1_decoder1.U160.ZN ) ,
    .I0 ( config1_decoder1.U160.AB ) ,
    .I1 ( config1_decoder1.n4 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_0_97 ) ,
    .IN ( config1_decoder1.U160.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder6.n2 ) ,
    .IN ( config1_decoder6.n1 ) ) ;
nand ( 
    .Z ( config1_decoder6.n71 ) ,
    .I0 ( config1_decoder6.n70 ) ,
    .I1 ( config1_decoder6.n76 ) ) ;
or ( 
    .Z ( config1_decoder6.U111.AB ) ,
    .I0 ( config1_decoder6.n93 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U111.ZN ) ,
    .I0 ( config1_decoder6.U111.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_78 ) ,
    .IN ( config1_decoder6.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U107.AB ) ,
    .I0 ( config1_decoder6.n89 ) ,
    .I1 ( config1_decoder6.n88 ) ) ;
and ( 
    .Z ( config1_decoder6.U107.ZN ) ,
    .I0 ( config1_decoder6.U107.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_87 ) ,
    .IN ( config1_decoder6.U107.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U135.AB ) ,
    .I0 ( config1_decoder6.n97 ) ,
    .I1 ( config1_decoder6.n98 ) ) ;
and ( 
    .Z ( config1_decoder6.U135.ZN ) ,
    .I0 ( config1_decoder6.U135.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_97 ) ,
    .IN ( config1_decoder6.U135.ZN ) ) ;
nor ( 
    .Z ( config1_decoder6.n77 ) ,
    .I0 ( config1_decoder6.n62 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
or ( 
    .Z ( config1_decoder6.U151.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n89 ) ) ;
and ( 
    .Z ( config1_decoder6.U151.ZN ) ,
    .I0 ( config1_decoder6.U151.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_71 ) ,
    .IN ( config1_decoder6.U151.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U59.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U59.ZN ) ,
    .I0 ( config1_decoder6.U59.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_39 ) ,
    .IN ( config1_decoder6.U59.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U49.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U49.ZN ) ,
    .I0 ( config1_decoder6.U49.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_21 ) ,
    .IN ( config1_decoder6.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U75.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U75.ZN ) ,
    .I0 ( config1_decoder6.U75.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_19 ) ,
    .IN ( config1_decoder6.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U65.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U65.ZN ) ,
    .I0 ( config1_decoder6.U65.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_40 ) ,
    .IN ( config1_decoder6.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U12.AB ) ,
    .I0 ( config1_decoder6.n83 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U12.ZN ) ,
    .I0 ( config1_decoder6.U12.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_14 ) ,
    .IN ( config1_decoder6.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n81 ) ,
    .I0 ( config1_decoder6.n79 ) ,
    .I1 ( config1_decoder6.n64 ) ) ;
nand ( 
    .Z ( config1_decoder6.n91 ) ,
    .I0 ( config1_decoder6.n80 ) ,
    .I1 ( config1_decoder6.n78 ) ) ;
nand ( 
    .Z ( config1_decoder6.n93 ) ,
    .I0 ( config1_decoder6.n80 ) ,
    .I1 ( config1_decoder6.n79 ) ) ;
nor ( 
    .Z ( config1_decoder6.n80 ) ,
    .I0 ( config1_decoder6.n75 ) ,
    .I1 ( masks_hold_reg_9_9 ) ) ;
nor ( 
    .Z ( config1_decoder6.n66 ) ,
    .I0 ( config1_decoder6.n65 ) ,
    .I1 ( masks_hold_reg_10_9 ) ) ;
or ( 
    .Z ( config1_decoder6.U155.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n90 ) ) ;
and ( 
    .Z ( config1_decoder6.U155.ZN ) ,
    .I0 ( config1_decoder6.U155.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_64 ) ,
    .IN ( config1_decoder6.U155.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U143.AB ) ,
    .I0 ( config1_decoder6.n91 ) ,
    .I1 ( config1_decoder6.n88 ) ) ;
and ( 
    .Z ( config1_decoder6.U143.ZN ) ,
    .I0 ( config1_decoder6.U143.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_89 ) ,
    .IN ( config1_decoder6.U143.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U163.AB ) ,
    .I0 ( config1_decoder6.n98 ) ,
    .I1 ( config1_decoder6.n96 ) ) ;
and ( 
    .Z ( config1_decoder6.U163.ZN ) ,
    .I0 ( config1_decoder6.U163.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_96 ) ,
    .IN ( config1_decoder6.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U92.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U92.ZN ) ,
    .I0 ( config1_decoder6.U92.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_27 ) ,
    .IN ( config1_decoder6.U92.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U80.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U80.ZN ) ,
    .I0 ( config1_decoder6.U80.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_7 ) ,
    .IN ( config1_decoder6.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U48.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n82 ) ) ;
and ( 
    .Z ( config1_decoder6.U48.ZN ) ,
    .I0 ( config1_decoder6.U48.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_5 ) ,
    .IN ( config1_decoder6.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U64.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U64.ZN ) ,
    .I0 ( config1_decoder6.U64.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_41 ) ,
    .IN ( config1_decoder6.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U13.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U13.ZN ) ,
    .I0 ( config1_decoder6.U13.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_15 ) ,
    .IN ( config1_decoder6.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n87 ) ,
    .I0 ( config1_decoder6.n77 ) ,
    .I1 ( config1_decoder6.n64 ) ) ;
nand ( 
    .Z ( config1_decoder6.n104 ) ,
    .I0 ( config1_decoder6.n64 ) ,
    .I1 ( config1_decoder6.n78 ) ) ;
nor ( 
    .Z ( config1_decoder6.n70 ) ,
    .I0 ( config1_decoder6.n69 ) ,
    .I1 ( masks_hold_reg_9_10 ) ) ;
nand ( 
    .Z ( config1_decoder6.n86 ) ,
    .I0 ( config1_decoder6.n66 ) ,
    .I1 ( masks_hold_reg_10_8 ) ) ;
or ( 
    .Z ( config1_decoder6.U154.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n90 ) ) ;
and ( 
    .Z ( config1_decoder6.U154.ZN ) ,
    .I0 ( config1_decoder6.U154.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_68 ) ,
    .IN ( config1_decoder6.U154.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U144.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n89 ) ) ;
and ( 
    .Z ( config1_decoder6.U144.ZN ) ,
    .I0 ( config1_decoder6.U144.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_67 ) ,
    .IN ( config1_decoder6.U144.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U160.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U160.ZN ) ,
    .I0 ( config1_decoder6.U160.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_62 ) ,
    .IN ( config1_decoder6.U160.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n79 ) ,
    .IN ( config1_decoder6.n99 ) ) ;
or ( 
    .Z ( config1_decoder6.U98.AB ) ,
    .I0 ( config1_decoder6.n97 ) ,
    .I1 ( config1_decoder6.n101 ) ) ;
and ( 
    .Z ( config1_decoder6.U98.ZN ) ,
    .I0 ( config1_decoder6.U98.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_101 ) ,
    .IN ( config1_decoder6.U98.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U83.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U83.ZN ) ,
    .I0 ( config1_decoder6.U83.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_3 ) ,
    .IN ( config1_decoder6.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U50.AB ) ,
    .I0 ( config1_decoder6.n87 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U50.ZN ) ,
    .I0 ( config1_decoder6.U50.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_20 ) ,
    .IN ( config1_decoder6.U50.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n89 ) ,
    .I0 ( config1_decoder6.n80 ) ,
    .I1 ( config1_decoder6.n76 ) ) ;
nand ( 
    .Z ( config1_decoder6.n1 ) ,
    .I0 ( config1_decoder6.n94 ) ,
    .I1 ( config1_decoder6.n60 ) ) ;
or ( 
    .Z ( config1_decoder6.U157.AB ) ,
    .I0 ( config1_decoder6.n93 ) ,
    .I1 ( config1_decoder6.n92 ) ) ;
and ( 
    .Z ( config1_decoder6.U157.ZN ) ,
    .I0 ( config1_decoder6.U157.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_94 ) ,
    .IN ( config1_decoder6.U157.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U145.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n89 ) ) ;
and ( 
    .Z ( config1_decoder6.U145.ZN ) ,
    .I0 ( config1_decoder6.U145.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_63 ) ,
    .IN ( config1_decoder6.U145.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U161.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n93 ) ) ;
and ( 
    .Z ( config1_decoder6.U161.ZN ) ,
    .I0 ( config1_decoder6.U161.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_66 ) ,
    .IN ( config1_decoder6.U161.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U82.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n87 ) ) ;
and ( 
    .Z ( config1_decoder6.U82.ZN ) ,
    .I0 ( config1_decoder6.U82.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_0 ) ,
    .IN ( config1_decoder6.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U89.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U89.ZN ) ,
    .I0 ( config1_decoder6.U89.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_49 ) ,
    .IN ( config1_decoder6.U89.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.U51.BN ) ,
    .IN ( config1_decoder6.n103 ) ) ;
nand ( 
    .Z ( config1_decoder6.n63 ) ,
    .I0 ( config1_decoder6.U51.BN ) ,
    .I1 ( config1_decoder6.n94 ) ) ;
nor ( 
    .Z ( config1_decoder6.n94 ) ,
    .I0 ( config1_decoder6.n75 ) ,
    .I1 ( config1_decoder6.n69 ) ) ;
or ( 
    .Z ( config1_decoder6.U78.AB ) ,
    .I0 ( config1_decoder6.n90 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U78.ZN ) ,
    .I0 ( config1_decoder6.U78.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_76 ) ,
    .IN ( config1_decoder6.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n90 ) ,
    .I0 ( config1_decoder6.n80 ) ,
    .I1 ( config1_decoder6.n77 ) ) ;
nor ( 
    .Z ( config1_decoder6.n61 ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( masks_hold_reg_10_10 ) ) ;
or ( 
    .Z ( config1_decoder6.U156.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n93 ) ) ;
and ( 
    .Z ( config1_decoder6.U156.ZN ) ,
    .I0 ( config1_decoder6.U156.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_70 ) ,
    .IN ( config1_decoder6.U156.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U146.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n91 ) ) ;
and ( 
    .Z ( config1_decoder6.U146.ZN ) ,
    .I0 ( config1_decoder6.U146.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_69 ) ,
    .IN ( config1_decoder6.U146.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U5.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U5.ZN ) ,
    .I0 ( config1_decoder6.U5.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_34 ) ,
    .IN ( config1_decoder6.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U88.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U88.ZN ) ,
    .I0 ( config1_decoder6.U88.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_55 ) ,
    .IN ( config1_decoder6.U88.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U52.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n87 ) ) ;
and ( 
    .Z ( config1_decoder6.U52.ZN ) ,
    .I0 ( config1_decoder6.U52.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_24 ) ,
    .IN ( config1_decoder6.U52.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n84 ) ,
    .I0 ( config1_decoder6.n76 ) ,
    .I1 ( config1_decoder6.n64 ) ) ;
or ( 
    .Z ( config1_decoder6.U79.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n87 ) ) ;
and ( 
    .Z ( config1_decoder6.U79.ZN ) ,
    .I0 ( config1_decoder6.U79.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_4 ) ,
    .IN ( config1_decoder6.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U72.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n87 ) ) ;
and ( 
    .Z ( config1_decoder6.U72.ZN ) ,
    .I0 ( config1_decoder6.U72.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_28 ) ,
    .IN ( config1_decoder6.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U69.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U69.ZN ) ,
    .I0 ( config1_decoder6.U69.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_48 ) ,
    .IN ( config1_decoder6.U69.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n82 ) ,
    .I0 ( config1_decoder6.n61 ) ,
    .I1 ( masks_hold_reg_10_8 ) ) ;
nand ( 
    .Z ( config1_decoder6.n88 ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( config1_decoder6.n67 ) ,
    .I2 ( masks_hold_reg_10_10 ) ) ;
or ( 
    .Z ( config1_decoder6.U159.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n90 ) ) ;
and ( 
    .Z ( config1_decoder6.U159.ZN ) ,
    .I0 ( config1_decoder6.U159.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_92 ) ,
    .IN ( config1_decoder6.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U147.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n91 ) ) ;
and ( 
    .Z ( config1_decoder6.U147.ZN ) ,
    .I0 ( config1_decoder6.U147.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_93 ) ,
    .IN ( config1_decoder6.U147.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U9.AB ) ,
    .I0 ( config1_decoder6.n83 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U9.ZN ) ,
    .I0 ( config1_decoder6.U9.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_44 ) ,
    .IN ( config1_decoder6.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U4.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U4.ZN ) ,
    .I0 ( config1_decoder6.U4.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_32 ) ,
    .IN ( config1_decoder6.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U53.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n87 ) ) ;
and ( 
    .Z ( config1_decoder6.U53.ZN ) ,
    .I0 ( config1_decoder6.U53.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_8 ) ,
    .IN ( config1_decoder6.U53.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.U43.BN ) ,
    .IN ( config1_decoder6.n82 ) ) ;
nand ( 
    .Z ( config1_decoder6.n101 ) ,
    .I0 ( config1_decoder6.U43.BN ) ,
    .I1 ( config1_decoder6.n94 ) ) ;
or ( 
    .Z ( config1_decoder6.U73.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U73.ZN ) ,
    .I0 ( config1_decoder6.U73.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_30 ) ,
    .IN ( config1_decoder6.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U68.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U68.ZN ) ,
    .I0 ( config1_decoder6.U68.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_51 ) ,
    .IN ( config1_decoder6.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U63.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U63.ZN ) ,
    .I0 ( config1_decoder6.U63.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_31 ) ,
    .IN ( config1_decoder6.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U14.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n95 ) ) ;
and ( 
    .Z ( config1_decoder6.U14.ZN ) ,
    .I0 ( config1_decoder6.U14.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_1 ) ,
    .IN ( config1_decoder6.U14.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n103 ) ,
    .I0 ( config1_decoder6.n67 ) ,
    .I1 ( config1_decoder6.n65 ) ,
    .I2 ( masks_hold_reg_10_9 ) ) ;
nand ( 
    .Z ( config1_decoder6.n92 ) ,
    .I0 ( masks_hold_reg_10_10 ) ,
    .I1 ( config1_decoder6.n68 ) ) ;
or ( 
    .Z ( config1_decoder6.U108.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n89 ) ) ;
and ( 
    .Z ( config1_decoder6.U108.ZN ) ,
    .I0 ( config1_decoder6.U108.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_91 ) ,
    .IN ( config1_decoder6.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U105.AB ) ,
    .I0 ( config1_decoder6.n91 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U105.ZN ) ,
    .I0 ( config1_decoder6.U105.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_85 ) ,
    .IN ( config1_decoder6.U105.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U137.AB ) ,
    .I0 ( config1_decoder6.n96 ) ,
    .I1 ( config1_decoder6.n63 ) ) ;
and ( 
    .Z ( config1_decoder6.U137.ZN ) ,
    .I0 ( config1_decoder6.U137.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_104 ) ,
    .IN ( config1_decoder6.U137.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U158.AB ) ,
    .I0 ( config1_decoder6.n90 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U158.ZN ) ,
    .I0 ( config1_decoder6.U158.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_80 ) ,
    .IN ( config1_decoder6.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U148.AB ) ,
    .I0 ( config1_decoder6.n89 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U148.ZN ) ,
    .I0 ( config1_decoder6.U148.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_79 ) ,
    .IN ( config1_decoder6.U148.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U164.AB ) ,
    .I0 ( config1_decoder6.n97 ) ,
    .I1 ( config1_decoder6.n63 ) ) ;
and ( 
    .Z ( config1_decoder6.U164.ZN ) ,
    .I0 ( config1_decoder6.U164.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_105 ) ,
    .IN ( config1_decoder6.U164.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n100 ) ,
    .IN ( config1_decoder6.n76 ) ) ;
or ( 
    .Z ( config1_decoder6.U8.AB ) ,
    .I0 ( config1_decoder6.n83 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U8.ZN ) ,
    .I0 ( config1_decoder6.U8.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_45 ) ,
    .IN ( config1_decoder6.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U7.AB ) ,
    .I0 ( config1_decoder6.n83 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U7.ZN ) ,
    .I0 ( config1_decoder6.U7.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_46 ) ,
    .IN ( config1_decoder6.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U54.AB ) ,
    .I0 ( config1_decoder6.n87 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U54.ZN ) ,
    .I0 ( config1_decoder6.U54.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_16 ) ,
    .IN ( config1_decoder6.U54.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n95 ) ,
    .I0 ( config1_decoder6.n61 ) ,
    .I1 ( config1_decoder6.n67 ) ) ;
or ( 
    .Z ( config1_decoder6.U70.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U70.ZN ) ,
    .I0 ( config1_decoder6.U70.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_22 ) ,
    .IN ( config1_decoder6.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U62.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U62.ZN ) ,
    .I0 ( config1_decoder6.U62.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_38 ) ,
    .IN ( config1_decoder6.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U15.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U15.ZN ) ,
    .I0 ( config1_decoder6.U15.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_13 ) ,
    .IN ( config1_decoder6.U15.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n67 ) ,
    .IN ( masks_hold_reg_10_8 ) ) ;
or ( 
    .Z ( config1_decoder6.U109.AB ) ,
    .I0 ( config1_decoder6.n93 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U109.ZN ) ,
    .I0 ( config1_decoder6.U109.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_82 ) ,
    .IN ( config1_decoder6.U109.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U106.AB ) ,
    .I0 ( config1_decoder6.n91 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U106.ZN ) ,
    .I0 ( config1_decoder6.U106.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_77 ) ,
    .IN ( config1_decoder6.U106.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U136.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U136.ZN ) ,
    .I0 ( config1_decoder6.U136.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_58 ) ,
    .IN ( config1_decoder6.U136.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n65 ) ,
    .IN ( masks_hold_reg_10_10 ) ) ;
or ( 
    .Z ( config1_decoder6.U149.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U149.ZN ) ,
    .I0 ( config1_decoder6.U149.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_61 ) ,
    .IN ( config1_decoder6.U149.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U165.AB ) ,
    .I0 ( config1_decoder6.n100 ) ,
    .I1 ( config1_decoder6.n63 ) ) ;
and ( 
    .Z ( config1_decoder6.U165.ZN ) ,
    .I0 ( config1_decoder6.U165.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_103 ) ,
    .IN ( config1_decoder6.U165.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n96 ) ,
    .IN ( config1_decoder6.n77 ) ) ;
or ( 
    .Z ( config1_decoder6.U6.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U6.ZN ) ,
    .I0 ( config1_decoder6.U6.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_47 ) ,
    .IN ( config1_decoder6.U6.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U85.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U85.ZN ) ,
    .I0 ( config1_decoder6.U85.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_59 ) ,
    .IN ( config1_decoder6.U85.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n78 ) ,
    .IN ( config1_decoder6.n97 ) ) ;
or ( 
    .Z ( config1_decoder6.U45.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n88 ) ) ;
and ( 
    .Z ( config1_decoder6.U45.ZN ) ,
    .I0 ( config1_decoder6.U45.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_25 ) ,
    .IN ( config1_decoder6.U45.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U71.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U71.ZN ) ,
    .I0 ( config1_decoder6.U71.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_10 ) ,
    .IN ( config1_decoder6.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U61.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U61.ZN ) ,
    .I0 ( config1_decoder6.U61.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_36 ) ,
    .IN ( config1_decoder6.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U16.AB ) ,
    .I0 ( config1_decoder6.n87 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U16.ZN ) ,
    .I0 ( config1_decoder6.U16.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_12 ) ,
    .IN ( config1_decoder6.U16.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U96.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U96.ZN ) ,
    .I0 ( config1_decoder6.U96.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_2 ) ,
    .IN ( config1_decoder6.U96.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.U1.BN ) ,
    .IN ( config1_decoder6.n95 ) ) ;
nand ( 
    .Z ( config1_decoder6.n98 ) ,
    .I0 ( config1_decoder6.U1.BN ) ,
    .I1 ( config1_decoder6.n94 ) ) ;
or ( 
    .Z ( config1_decoder6.U84.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U84.ZN ) ,
    .I0 ( config1_decoder6.U84.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_57 ) ,
    .IN ( config1_decoder6.U84.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U56.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U56.ZN ) ,
    .I0 ( config1_decoder6.U56.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_26 ) ,
    .IN ( config1_decoder6.U56.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n83 ) ,
    .I0 ( config1_decoder6.n68 ) ,
    .I1 ( config1_decoder6.n65 ) ) ;
or ( 
    .Z ( config1_decoder6.U76.AB ) ,
    .I0 ( config1_decoder6.n89 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U76.ZN ) ,
    .I0 ( config1_decoder6.U76.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_83 ) ,
    .IN ( config1_decoder6.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U60.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U60.ZN ) ,
    .I0 ( config1_decoder6.U60.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_37 ) ,
    .IN ( config1_decoder6.U60.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U17.AB ) ,
    .I0 ( config1_decoder6.n84 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U17.ZN ) ,
    .I0 ( config1_decoder6.U17.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_11 ) ,
    .IN ( config1_decoder6.U17.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n72 ) ,
    .I0 ( config1_decoder6.n70 ) ,
    .I1 ( config1_decoder6.n77 ) ) ;
or ( 
    .Z ( config1_decoder6.U27.AB ) ,
    .I0 ( config1_decoder6.n91 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U27.ZN ) ,
    .I0 ( config1_decoder6.U27.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_81 ) ,
    .IN ( config1_decoder6.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U110.AB ) ,
    .I0 ( config1_decoder6.n93 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U110.ZN ) ,
    .I0 ( config1_decoder6.U110.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_86 ) ,
    .IN ( config1_decoder6.U110.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n69 ) ,
    .IN ( masks_hold_reg_9_9 ) ) ;
or ( 
    .Z ( config1_decoder6.U134.AB ) ,
    .I0 ( config1_decoder6.n101 ) ,
    .I1 ( config1_decoder6.n96 ) ) ;
and ( 
    .Z ( config1_decoder6.U134.ZN ) ,
    .I0 ( config1_decoder6.U134.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_100 ) ,
    .IN ( config1_decoder6.U134.ZN ) ) ;
nor ( 
    .Z ( config1_decoder6.n76 ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
or ( 
    .Z ( config1_decoder6.U150.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n91 ) ) ;
and ( 
    .Z ( config1_decoder6.U150.ZN ) ,
    .I0 ( config1_decoder6.U150.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_65 ) ,
    .IN ( config1_decoder6.U150.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U140.AB ) ,
    .I0 ( config1_decoder6.n101 ) ,
    .I1 ( config1_decoder6.n100 ) ) ;
and ( 
    .Z ( config1_decoder6.U140.ZN ) ,
    .I0 ( config1_decoder6.U140.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_99 ) ,
    .IN ( config1_decoder6.U140.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U97.AB ) ,
    .I0 ( config1_decoder6.n92 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U97.ZN ) ,
    .I0 ( config1_decoder6.U97.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_60 ) ,
    .IN ( config1_decoder6.U97.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U87.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U87.ZN ) ,
    .I0 ( config1_decoder6.U87.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_56 ) ,
    .IN ( config1_decoder6.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U57.AB ) ,
    .I0 ( config1_decoder6.n88 ) ,
    .I1 ( config1_decoder6.n84 ) ) ;
and ( 
    .Z ( config1_decoder6.U57.ZN ) ,
    .I0 ( config1_decoder6.U57.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_23 ) ,
    .IN ( config1_decoder6.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U47.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n103 ) ) ;
and ( 
    .Z ( config1_decoder6.U47.ZN ) ,
    .I0 ( config1_decoder6.U47.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_9 ) ,
    .IN ( config1_decoder6.U47.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U77.AB ) ,
    .I0 ( config1_decoder6.n89 ) ,
    .I1 ( config1_decoder6.n83 ) ) ;
and ( 
    .Z ( config1_decoder6.U77.ZN ) ,
    .I0 ( config1_decoder6.U77.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_75 ) ,
    .IN ( config1_decoder6.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U67.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n72 ) ) ;
and ( 
    .Z ( config1_decoder6.U67.ZN ) ,
    .I0 ( config1_decoder6.U67.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_52 ) ,
    .IN ( config1_decoder6.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U10.AB ) ,
    .I0 ( config1_decoder6.n83 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U10.ZN ) ,
    .I0 ( config1_decoder6.U10.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_43 ) ,
    .IN ( config1_decoder6.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n85 ) ,
    .I0 ( config1_decoder6.n66 ) ,
    .I1 ( config1_decoder6.n67 ) ) ;
or ( 
    .Z ( config1_decoder6.U26.AB ) ,
    .I0 ( config1_decoder6.n90 ) ,
    .I1 ( config1_decoder6.n86 ) ) ;
and ( 
    .Z ( config1_decoder6.U26.ZN ) ,
    .I0 ( config1_decoder6.U26.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_84 ) ,
    .IN ( config1_decoder6.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U113.AB ) ,
    .I0 ( config1_decoder6.n90 ) ,
    .I1 ( config1_decoder6.n88 ) ) ;
and ( 
    .Z ( config1_decoder6.U113.ZN ) ,
    .I0 ( config1_decoder6.U113.AB ) ,
    .I1 ( config1_decoder6.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_88 ) ,
    .IN ( config1_decoder6.U113.ZN ) ) ;
not ( 
    .O1 ( config1_decoder6.n75 ) ,
    .IN ( masks_hold_reg_9_10 ) ) ;
not ( 
    .O1 ( config1_decoder6.n62 ) ,
    .IN ( masks_hold_reg_10_6 ) ) ;
nor ( 
    .Z ( config1_decoder6.n64 ) ,
    .I0 ( masks_hold_reg_9_9 ) ,
    .I1 ( masks_hold_reg_9_10 ) ) ;
nand ( 
    .Z ( config1_decoder6.n97 ) ,
    .I0 ( masks_hold_reg_10_7 ) ,
    .I1 ( config1_decoder6.n62 ) ) ;
or ( 
    .Z ( config1_decoder6.U153.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n93 ) ) ;
and ( 
    .Z ( config1_decoder6.U153.ZN ) ,
    .I0 ( config1_decoder6.U153.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_74 ) ,
    .IN ( config1_decoder6.U153.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U141.AB ) ,
    .I0 ( config1_decoder6.n99 ) ,
    .I1 ( config1_decoder6.n98 ) ) ;
and ( 
    .Z ( config1_decoder6.U141.ZN ) ,
    .I0 ( config1_decoder6.U141.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_98 ) ,
    .IN ( config1_decoder6.U141.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U90.AB ) ,
    .I0 ( config1_decoder6.n99 ) ,
    .I1 ( config1_decoder6.n101 ) ) ;
and ( 
    .Z ( config1_decoder6.U90.ZN ) ,
    .I0 ( config1_decoder6.U90.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_102 ) ,
    .IN ( config1_decoder6.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U3.AB ) ,
    .I0 ( config1_decoder6.n95 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U3.ZN ) ,
    .I0 ( config1_decoder6.U3.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_33 ) ,
    .IN ( config1_decoder6.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U86.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n73 ) ) ;
and ( 
    .Z ( config1_decoder6.U86.ZN ) ,
    .I0 ( config1_decoder6.U86.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_53 ) ,
    .IN ( config1_decoder6.U86.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U58.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n71 ) ) ;
and ( 
    .Z ( config1_decoder6.U58.ZN ) ,
    .I0 ( config1_decoder6.U58.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_35 ) ,
    .IN ( config1_decoder6.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U46.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n92 ) ) ;
and ( 
    .Z ( config1_decoder6.U46.ZN ) ,
    .I0 ( config1_decoder6.U46.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_29 ) ,
    .IN ( config1_decoder6.U46.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U74.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U74.ZN ) ,
    .I0 ( config1_decoder6.U74.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_18 ) ,
    .IN ( config1_decoder6.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U66.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U66.ZN ) ,
    .I0 ( config1_decoder6.U66.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_42 ) ,
    .IN ( config1_decoder6.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U11.AB ) ,
    .I0 ( config1_decoder6.n85 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U11.ZN ) ,
    .I0 ( config1_decoder6.U11.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_50 ) ,
    .IN ( config1_decoder6.U11.ZN ) ) ;
nand ( 
    .Z ( config1_decoder6.n73 ) ,
    .I0 ( config1_decoder6.n70 ) ,
    .I1 ( config1_decoder6.n78 ) ) ;
nand ( 
    .Z ( config1_decoder6.n74 ) ,
    .I0 ( config1_decoder6.n70 ) ,
    .I1 ( config1_decoder6.n79 ) ) ;
or ( 
    .Z ( config1_decoder6.U112.AB ) ,
    .I0 ( config1_decoder6.n93 ) ,
    .I1 ( config1_decoder6.n88 ) ) ;
and ( 
    .Z ( config1_decoder6.U112.ZN ) ,
    .I0 ( config1_decoder6.U112.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_90 ) ,
    .IN ( config1_decoder6.U112.ZN ) ) ;
and ( 
    .Z ( config1_decoder6.n68 ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( masks_hold_reg_10_8 ) ) ;
nand ( 
    .Z ( config1_decoder6.n99 ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( masks_hold_reg_10_7 ) ) ;
and ( 
    .Z ( config1_decoder6.U122.AB ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( config1_decoder6.n79 ) ) ;
or ( 
    .Z ( config1_decoder6.n60 ) ,
    .I0 ( config1_decoder6.U122.AB ) ,
    .I1 ( config1_decoder6.n68 ) ,
    .I2 ( masks_hold_reg_10_10 ) ) ;
or ( 
    .Z ( config1_decoder6.U152.AB ) ,
    .I0 ( config1_decoder6.n100 ) ,
    .I1 ( config1_decoder6.n98 ) ) ;
and ( 
    .Z ( config1_decoder6.U152.ZN ) ,
    .I0 ( config1_decoder6.U152.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_95 ) ,
    .IN ( config1_decoder6.U152.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U142.AB ) ,
    .I0 ( config1_decoder6.n86 ) ,
    .I1 ( config1_decoder6.n74 ) ) ;
and ( 
    .Z ( config1_decoder6.U142.ZN ) ,
    .I0 ( config1_decoder6.U142.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_54 ) ,
    .IN ( config1_decoder6.U142.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U162.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n90 ) ) ;
and ( 
    .Z ( config1_decoder6.U162.ZN ) ,
    .I0 ( config1_decoder6.U162.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_72 ) ,
    .IN ( config1_decoder6.U162.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U91.AB ) ,
    .I0 ( config1_decoder6.n103 ) ,
    .I1 ( config1_decoder6.n91 ) ) ;
and ( 
    .Z ( config1_decoder6.U91.ZN ) ,
    .I0 ( config1_decoder6.U91.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_73 ) ,
    .IN ( config1_decoder6.U91.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U2.AB ) ,
    .I0 ( config1_decoder6.n104 ) ,
    .I1 ( config1_decoder6.n85 ) ) ;
and ( 
    .Z ( config1_decoder6.U2.ZN ) ,
    .I0 ( config1_decoder6.U2.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_17 ) ,
    .IN ( config1_decoder6.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder6.U81.AB ) ,
    .I0 ( config1_decoder6.n82 ) ,
    .I1 ( config1_decoder6.n81 ) ) ;
and ( 
    .Z ( config1_decoder6.U81.ZN ) ,
    .I0 ( config1_decoder6.U81.AB ) ,
    .I1 ( config1_decoder6.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_5_6 ) ,
    .IN ( config1_decoder6.U81.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder7.n2 ) ,
    .IN ( config1_decoder7.n1 ) ) ;
or ( 
    .Z ( config1_decoder7.U110.AB ) ,
    .I0 ( config1_decoder7.n89 ) ,
    .I1 ( config1_decoder7.n88 ) ) ;
and ( 
    .Z ( config1_decoder7.U110.ZN ) ,
    .I0 ( config1_decoder7.U110.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_87 ) ,
    .IN ( config1_decoder7.U110.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n96 ) ,
    .IN ( config1_decoder7.n77 ) ) ;
nand ( 
    .Z ( config1_decoder7.n99 ) ,
    .I0 ( masks_hold_reg_12_7 ) ,
    .I1 ( masks_hold_reg_12_8 ) ) ;
nor ( 
    .Z ( config1_decoder7.n77 ) ,
    .I0 ( config1_decoder7.n62 ) ,
    .I1 ( masks_hold_reg_12_8 ) ) ;
nand ( 
    .Z ( config1_decoder7.n86 ) ,
    .I0 ( config1_decoder7.n66 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
or ( 
    .Z ( config1_decoder7.U150.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n91 ) ) ;
and ( 
    .Z ( config1_decoder7.U150.ZN ) ,
    .I0 ( config1_decoder7.U150.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_69 ) ,
    .IN ( config1_decoder7.U150.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n62 ) ,
    .IN ( masks_hold_reg_12_7 ) ) ;
or ( 
    .Z ( config1_decoder7.U97.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U97.ZN ) ,
    .I0 ( config1_decoder7.U97.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_27 ) ,
    .IN ( config1_decoder7.U97.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U87.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U87.ZN ) ,
    .I0 ( config1_decoder7.U87.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_59 ) ,
    .IN ( config1_decoder7.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U57.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U57.ZN ) ,
    .I0 ( config1_decoder7.U57.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_23 ) ,
    .IN ( config1_decoder7.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U47.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U47.ZN ) ,
    .I0 ( config1_decoder7.U47.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_21 ) ,
    .IN ( config1_decoder7.U47.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U13.AB ) ,
    .I0 ( config1_decoder7.n83 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U13.ZN ) ,
    .I0 ( config1_decoder7.U13.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_14 ) ,
    .IN ( config1_decoder7.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n90 ) ,
    .I0 ( config1_decoder7.n80 ) ,
    .I1 ( config1_decoder7.n77 ) ) ;
or ( 
    .Z ( config1_decoder7.U28.AB ) ,
    .I0 ( config1_decoder7.n91 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U28.ZN ) ,
    .I0 ( config1_decoder7.U28.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_81 ) ,
    .IN ( config1_decoder7.U28.ZN ) ) ;
nor ( 
    .Z ( config1_decoder7.n66 ) ,
    .I0 ( config1_decoder7.n65 ) ,
    .I1 ( masks_hold_reg_12_10 ) ) ;
or ( 
    .Z ( config1_decoder7.U120.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n90 ) ) ;
and ( 
    .Z ( config1_decoder7.U120.ZN ) ,
    .I0 ( config1_decoder7.U120.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_92 ) ,
    .IN ( config1_decoder7.U120.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U154.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n89 ) ) ;
and ( 
    .Z ( config1_decoder7.U154.ZN ) ,
    .I0 ( config1_decoder7.U154.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_71 ) ,
    .IN ( config1_decoder7.U154.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n69 ) ,
    .IN ( masks_hold_reg_11_10 ) ) ;
or ( 
    .Z ( config1_decoder7.U160.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U160.ZN ) ,
    .I0 ( config1_decoder7.U160.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_62 ) ,
    .IN ( config1_decoder7.U160.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U93.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U93.ZN ) ,
    .I0 ( config1_decoder7.U93.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_49 ) ,
    .IN ( config1_decoder7.U93.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n79 ) ,
    .IN ( config1_decoder7.n99 ) ) ;
or ( 
    .Z ( config1_decoder7.U83.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U83.ZN ) ,
    .I0 ( config1_decoder7.U83.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_3 ) ,
    .IN ( config1_decoder7.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U50.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n92 ) ) ;
and ( 
    .Z ( config1_decoder7.U50.ZN ) ,
    .I0 ( config1_decoder7.U50.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_29 ) ,
    .IN ( config1_decoder7.U50.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n95 ) ,
    .I0 ( config1_decoder7.n61 ) ,
    .I1 ( config1_decoder7.n67 ) ) ;
nand ( 
    .Z ( config1_decoder7.n88 ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( config1_decoder7.n67 ) ,
    .I2 ( masks_hold_reg_11_9 ) ) ;
or ( 
    .Z ( config1_decoder7.U157.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n90 ) ) ;
and ( 
    .Z ( config1_decoder7.U157.ZN ) ,
    .I0 ( config1_decoder7.U157.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_64 ) ,
    .IN ( config1_decoder7.U157.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n75 ) ,
    .IN ( masks_hold_reg_10_0 ) ) ;
or ( 
    .Z ( config1_decoder7.U81.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U81.ZN ) ,
    .I0 ( config1_decoder7.U81.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_7 ) ,
    .IN ( config1_decoder7.U81.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n78 ) ,
    .IN ( config1_decoder7.n97 ) ) ;
or ( 
    .Z ( config1_decoder7.U49.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n103 ) ) ;
and ( 
    .Z ( config1_decoder7.U49.ZN ) ,
    .I0 ( config1_decoder7.U49.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_9 ) ,
    .IN ( config1_decoder7.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U75.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U75.ZN ) ,
    .I0 ( config1_decoder7.U75.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_31 ) ,
    .IN ( config1_decoder7.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U65.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U65.ZN ) ,
    .I0 ( config1_decoder7.U65.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_41 ) ,
    .IN ( config1_decoder7.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U12.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U12.ZN ) ,
    .I0 ( config1_decoder7.U12.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_50 ) ,
    .IN ( config1_decoder7.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n72 ) ,
    .I0 ( config1_decoder7.n70 ) ,
    .I1 ( config1_decoder7.n77 ) ) ;
nand ( 
    .Z ( config1_decoder7.n89 ) ,
    .I0 ( config1_decoder7.n80 ) ,
    .I1 ( config1_decoder7.n76 ) ) ;
nand ( 
    .Z ( config1_decoder7.n104 ) ,
    .I0 ( config1_decoder7.n64 ) ,
    .I1 ( config1_decoder7.n78 ) ) ;
nand ( 
    .Z ( config1_decoder7.n82 ) ,
    .I0 ( config1_decoder7.n61 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
not ( 
    .O1 ( config1_decoder7.n67 ) ,
    .IN ( masks_hold_reg_12_9 ) ) ;
or ( 
    .Z ( config1_decoder7.U155.AB ) ,
    .I0 ( config1_decoder7.n100 ) ,
    .I1 ( config1_decoder7.n98 ) ) ;
and ( 
    .Z ( config1_decoder7.U155.ZN ) ,
    .I0 ( config1_decoder7.U155.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_95 ) ,
    .IN ( config1_decoder7.U155.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U143.AB ) ,
    .I0 ( config1_decoder7.n96 ) ,
    .I1 ( config1_decoder7.n63 ) ) ;
and ( 
    .Z ( config1_decoder7.U143.ZN ) ,
    .I0 ( config1_decoder7.U143.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_104 ) ,
    .IN ( config1_decoder7.U143.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U163.AB ) ,
    .I0 ( config1_decoder7.n98 ) ,
    .I1 ( config1_decoder7.n96 ) ) ;
and ( 
    .Z ( config1_decoder7.U163.ZN ) ,
    .I0 ( config1_decoder7.U163.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_96 ) ,
    .IN ( config1_decoder7.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U92.AB ) ,
    .I0 ( config1_decoder7.n97 ) ,
    .I1 ( config1_decoder7.n101 ) ) ;
and ( 
    .Z ( config1_decoder7.U92.ZN ) ,
    .I0 ( config1_decoder7.U92.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_101 ) ,
    .IN ( config1_decoder7.U92.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U80.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n87 ) ) ;
and ( 
    .Z ( config1_decoder7.U80.ZN ) ,
    .I0 ( config1_decoder7.U80.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_4 ) ,
    .IN ( config1_decoder7.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U48.AB ) ,
    .I0 ( config1_decoder7.n87 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U48.ZN ) ,
    .I0 ( config1_decoder7.U48.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_20 ) ,
    .IN ( config1_decoder7.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U64.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U64.ZN ) ,
    .I0 ( config1_decoder7.U64.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_38 ) ,
    .IN ( config1_decoder7.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U161.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n93 ) ) ;
and ( 
    .Z ( config1_decoder7.U161.ZN ) ,
    .I0 ( config1_decoder7.U161.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_66 ) ,
    .IN ( config1_decoder7.U161.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.n100 ) ,
    .IN ( config1_decoder7.n76 ) ) ;
or ( 
    .Z ( config1_decoder7.U82.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U82.ZN ) ,
    .I0 ( config1_decoder7.U82.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_6 ) ,
    .IN ( config1_decoder7.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U89.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U89.ZN ) ,
    .I0 ( config1_decoder7.U89.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_56 ) ,
    .IN ( config1_decoder7.U89.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.U51.BN ) ,
    .IN ( config1_decoder7.n103 ) ) ;
nand ( 
    .Z ( config1_decoder7.n63 ) ,
    .I0 ( config1_decoder7.U51.BN ) ,
    .I1 ( config1_decoder7.n94 ) ) ;
nand ( 
    .Z ( config1_decoder7.n81 ) ,
    .I0 ( config1_decoder7.n79 ) ,
    .I1 ( config1_decoder7.n64 ) ) ;
or ( 
    .Z ( config1_decoder7.U78.AB ) ,
    .I0 ( config1_decoder7.n89 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U78.ZN ) ,
    .I0 ( config1_decoder7.U78.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_75 ) ,
    .IN ( config1_decoder7.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n93 ) ,
    .I0 ( config1_decoder7.n80 ) ,
    .I1 ( config1_decoder7.n79 ) ) ;
or ( 
    .Z ( config1_decoder7.U115.AB ) ,
    .I0 ( config1_decoder7.n93 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U115.ZN ) ,
    .I0 ( config1_decoder7.U115.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_78 ) ,
    .IN ( config1_decoder7.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U156.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n90 ) ) ;
and ( 
    .Z ( config1_decoder7.U156.ZN ) ,
    .I0 ( config1_decoder7.U156.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_68 ) ,
    .IN ( config1_decoder7.U156.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U146.AB ) ,
    .I0 ( config1_decoder7.n97 ) ,
    .I1 ( config1_decoder7.n98 ) ) ;
and ( 
    .Z ( config1_decoder7.U146.ZN ) ,
    .I0 ( config1_decoder7.U146.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_97 ) ,
    .IN ( config1_decoder7.U146.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U5.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U5.ZN ) ,
    .I0 ( config1_decoder7.U5.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_32 ) ,
    .IN ( config1_decoder7.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U88.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U88.ZN ) ,
    .I0 ( config1_decoder7.U88.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_53 ) ,
    .IN ( config1_decoder7.U88.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U52.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n87 ) ) ;
and ( 
    .Z ( config1_decoder7.U52.ZN ) ,
    .I0 ( config1_decoder7.U52.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_24 ) ,
    .IN ( config1_decoder7.U52.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n73 ) ,
    .I0 ( config1_decoder7.n70 ) ,
    .I1 ( config1_decoder7.n78 ) ) ;
or ( 
    .Z ( config1_decoder7.U79.AB ) ,
    .I0 ( config1_decoder7.n90 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U79.ZN ) ,
    .I0 ( config1_decoder7.U79.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_76 ) ,
    .IN ( config1_decoder7.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U72.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U72.ZN ) ,
    .I0 ( config1_decoder7.U72.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_10 ) ,
    .IN ( config1_decoder7.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U69.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U69.ZN ) ,
    .I0 ( config1_decoder7.U69.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_52 ) ,
    .IN ( config1_decoder7.U69.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U119.AB ) ,
    .I0 ( config1_decoder7.n90 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U119.ZN ) ,
    .I0 ( config1_decoder7.U119.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_80 ) ,
    .IN ( config1_decoder7.U119.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U114.AB ) ,
    .I0 ( config1_decoder7.n93 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U114.ZN ) ,
    .I0 ( config1_decoder7.U114.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_86 ) ,
    .IN ( config1_decoder7.U114.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U159.AB ) ,
    .I0 ( config1_decoder7.n93 ) ,
    .I1 ( config1_decoder7.n92 ) ) ;
and ( 
    .Z ( config1_decoder7.U159.ZN ) ,
    .I0 ( config1_decoder7.U159.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_94 ) ,
    .IN ( config1_decoder7.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U147.AB ) ,
    .I0 ( config1_decoder7.n99 ) ,
    .I1 ( config1_decoder7.n98 ) ) ;
and ( 
    .Z ( config1_decoder7.U147.ZN ) ,
    .I0 ( config1_decoder7.U147.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_98 ) ,
    .IN ( config1_decoder7.U147.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U9.AB ) ,
    .I0 ( config1_decoder7.n83 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U9.ZN ) ,
    .I0 ( config1_decoder7.U9.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_45 ) ,
    .IN ( config1_decoder7.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U4.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U4.ZN ) ,
    .I0 ( config1_decoder7.U4.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_33 ) ,
    .IN ( config1_decoder7.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U53.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n87 ) ) ;
and ( 
    .Z ( config1_decoder7.U53.ZN ) ,
    .I0 ( config1_decoder7.U53.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_8 ) ,
    .IN ( config1_decoder7.U53.ZN ) ) ;
nor ( 
    .Z ( config1_decoder7.n94 ) ,
    .I0 ( config1_decoder7.n75 ) ,
    .I1 ( config1_decoder7.n69 ) ) ;
or ( 
    .Z ( config1_decoder7.U73.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n87 ) ) ;
and ( 
    .Z ( config1_decoder7.U73.ZN ) ,
    .I0 ( config1_decoder7.U73.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_28 ) ,
    .IN ( config1_decoder7.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U68.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U68.ZN ) ,
    .I0 ( config1_decoder7.U68.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_54 ) ,
    .IN ( config1_decoder7.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U63.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U63.ZN ) ,
    .I0 ( config1_decoder7.U63.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_36 ) ,
    .IN ( config1_decoder7.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U14.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U14.ZN ) ,
    .I0 ( config1_decoder7.U14.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_15 ) ,
    .IN ( config1_decoder7.U14.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U118.AB ) ,
    .I0 ( config1_decoder7.n90 ) ,
    .I1 ( config1_decoder7.n88 ) ) ;
and ( 
    .Z ( config1_decoder7.U118.ZN ) ,
    .I0 ( config1_decoder7.U118.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_88 ) ,
    .IN ( config1_decoder7.U118.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U117.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n93 ) ) ;
and ( 
    .Z ( config1_decoder7.U117.ZN ) ,
    .I0 ( config1_decoder7.U117.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_74 ) ,
    .IN ( config1_decoder7.U117.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U108.AB ) ,
    .I0 ( config1_decoder7.n91 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U108.ZN ) ,
    .I0 ( config1_decoder7.U108.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_77 ) ,
    .IN ( config1_decoder7.U108.ZN ) ) ;
nor ( 
    .Z ( config1_decoder7.n80 ) ,
    .I0 ( config1_decoder7.n75 ) ,
    .I1 ( masks_hold_reg_11_10 ) ) ;
or ( 
    .Z ( config1_decoder7.U158.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n93 ) ) ;
and ( 
    .Z ( config1_decoder7.U158.ZN ) ,
    .I0 ( config1_decoder7.U158.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_70 ) ,
    .IN ( config1_decoder7.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U148.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n89 ) ) ;
and ( 
    .Z ( config1_decoder7.U148.ZN ) ,
    .I0 ( config1_decoder7.U148.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_67 ) ,
    .IN ( config1_decoder7.U148.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U164.AB ) ,
    .I0 ( config1_decoder7.n97 ) ,
    .I1 ( config1_decoder7.n63 ) ) ;
and ( 
    .Z ( config1_decoder7.U164.ZN ) ,
    .I0 ( config1_decoder7.U164.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_105 ) ,
    .IN ( config1_decoder7.U164.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U94.AB ) ,
    .I0 ( config1_decoder7.n99 ) ,
    .I1 ( config1_decoder7.n101 ) ) ;
and ( 
    .Z ( config1_decoder7.U94.ZN ) ,
    .I0 ( config1_decoder7.U94.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_102 ) ,
    .IN ( config1_decoder7.U94.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U8.AB ) ,
    .I0 ( config1_decoder7.n83 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U8.ZN ) ,
    .I0 ( config1_decoder7.U8.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_46 ) ,
    .IN ( config1_decoder7.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U7.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U7.ZN ) ,
    .I0 ( config1_decoder7.U7.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_47 ) ,
    .IN ( config1_decoder7.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U54.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n87 ) ) ;
and ( 
    .Z ( config1_decoder7.U54.ZN ) ,
    .I0 ( config1_decoder7.U54.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_0 ) ,
    .IN ( config1_decoder7.U54.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n84 ) ,
    .I0 ( config1_decoder7.n76 ) ,
    .I1 ( config1_decoder7.n64 ) ) ;
or ( 
    .Z ( config1_decoder7.U70.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U70.ZN ) ,
    .I0 ( config1_decoder7.U70.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_51 ) ,
    .IN ( config1_decoder7.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U62.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U62.ZN ) ,
    .I0 ( config1_decoder7.U62.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_37 ) ,
    .IN ( config1_decoder7.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U15.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U15.ZN ) ,
    .I0 ( config1_decoder7.U15.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_13 ) ,
    .IN ( config1_decoder7.U15.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U116.AB ) ,
    .I0 ( config1_decoder7.n93 ) ,
    .I1 ( config1_decoder7.n88 ) ) ;
and ( 
    .Z ( config1_decoder7.U116.ZN ) ,
    .I0 ( config1_decoder7.U116.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_90 ) ,
    .IN ( config1_decoder7.U116.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U109.AB ) ,
    .I0 ( config1_decoder7.n91 ) ,
    .I1 ( config1_decoder7.n88 ) ) ;
and ( 
    .Z ( config1_decoder7.U109.ZN ) ,
    .I0 ( config1_decoder7.U109.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_89 ) ,
    .IN ( config1_decoder7.U109.ZN ) ) ;
and ( 
    .Z ( config1_decoder7.n68 ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( masks_hold_reg_12_9 ) ) ;
nand ( 
    .Z ( config1_decoder7.n92 ) ,
    .I0 ( masks_hold_reg_11_9 ) ,
    .I1 ( config1_decoder7.n68 ) ) ;
or ( 
    .Z ( config1_decoder7.U149.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n89 ) ) ;
and ( 
    .Z ( config1_decoder7.U149.ZN ) ,
    .I0 ( config1_decoder7.U149.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_63 ) ,
    .IN ( config1_decoder7.U149.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U165.AB ) ,
    .I0 ( config1_decoder7.n100 ) ,
    .I1 ( config1_decoder7.n63 ) ) ;
and ( 
    .Z ( config1_decoder7.U165.ZN ) ,
    .I0 ( config1_decoder7.U165.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_103 ) ,
    .IN ( config1_decoder7.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U95.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n91 ) ) ;
and ( 
    .Z ( config1_decoder7.U95.ZN ) ,
    .I0 ( config1_decoder7.U95.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_73 ) ,
    .IN ( config1_decoder7.U95.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U6.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U6.ZN ) ,
    .I0 ( config1_decoder7.U6.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_34 ) ,
    .IN ( config1_decoder7.U6.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U85.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U85.ZN ) ,
    .I0 ( config1_decoder7.U85.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_57 ) ,
    .IN ( config1_decoder7.U85.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U55.AB ) ,
    .I0 ( config1_decoder7.n87 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U55.ZN ) ,
    .I0 ( config1_decoder7.U55.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_16 ) ,
    .IN ( config1_decoder7.U55.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.U45.BN ) ,
    .IN ( config1_decoder7.n82 ) ) ;
nand ( 
    .Z ( config1_decoder7.n101 ) ,
    .I0 ( config1_decoder7.U45.BN ) ,
    .I1 ( config1_decoder7.n94 ) ) ;
or ( 
    .Z ( config1_decoder7.U71.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U71.ZN ) ,
    .I0 ( config1_decoder7.U71.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_22 ) ,
    .IN ( config1_decoder7.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U61.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U61.ZN ) ,
    .I0 ( config1_decoder7.U61.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_39 ) ,
    .IN ( config1_decoder7.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U16.AB ) ,
    .I0 ( config1_decoder7.n87 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U16.ZN ) ,
    .I0 ( config1_decoder7.U16.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_12 ) ,
    .IN ( config1_decoder7.U16.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n85 ) ,
    .I0 ( config1_decoder7.n66 ) ,
    .I1 ( config1_decoder7.n67 ) ) ;
or ( 
    .Z ( config1_decoder7.U111.AB ) ,
    .I0 ( config1_decoder7.n89 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U111.ZN ) ,
    .I0 ( config1_decoder7.U111.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_79 ) ,
    .IN ( config1_decoder7.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U107.AB ) ,
    .I0 ( config1_decoder7.n91 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U107.ZN ) ,
    .I0 ( config1_decoder7.U107.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_85 ) ,
    .IN ( config1_decoder7.U107.ZN ) ) ;
nor ( 
    .Z ( config1_decoder7.n64 ) ,
    .I0 ( masks_hold_reg_11_10 ) ,
    .I1 ( masks_hold_reg_10_0 ) ) ;
not ( 
    .O1 ( config1_decoder7.n65 ) ,
    .IN ( masks_hold_reg_11_9 ) ) ;
or ( 
    .Z ( config1_decoder7.U151.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n91 ) ) ;
and ( 
    .Z ( config1_decoder7.U151.ZN ) ,
    .I0 ( config1_decoder7.U151.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_93 ) ,
    .IN ( config1_decoder7.U151.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U96.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n82 ) ) ;
and ( 
    .Z ( config1_decoder7.U96.ZN ) ,
    .I0 ( config1_decoder7.U96.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_5 ) ,
    .IN ( config1_decoder7.U96.ZN ) ) ;
not ( 
    .O1 ( config1_decoder7.U1.BN ) ,
    .IN ( config1_decoder7.n95 ) ) ;
nand ( 
    .Z ( config1_decoder7.n98 ) ,
    .I0 ( config1_decoder7.U1.BN ) ,
    .I1 ( config1_decoder7.n94 ) ) ;
or ( 
    .Z ( config1_decoder7.U84.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U84.ZN ) ,
    .I0 ( config1_decoder7.U84.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_2 ) ,
    .IN ( config1_decoder7.U84.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U56.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U56.ZN ) ,
    .I0 ( config1_decoder7.U56.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_26 ) ,
    .IN ( config1_decoder7.U56.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n83 ) ,
    .I0 ( config1_decoder7.n68 ) ,
    .I1 ( config1_decoder7.n65 ) ) ;
or ( 
    .Z ( config1_decoder7.U76.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U76.ZN ) ,
    .I0 ( config1_decoder7.U76.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_18 ) ,
    .IN ( config1_decoder7.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U60.AB ) ,
    .I0 ( config1_decoder7.n82 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U60.ZN ) ,
    .I0 ( config1_decoder7.U60.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_35 ) ,
    .IN ( config1_decoder7.U60.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U17.AB ) ,
    .I0 ( config1_decoder7.n84 ) ,
    .I1 ( config1_decoder7.n83 ) ) ;
and ( 
    .Z ( config1_decoder7.U17.ZN ) ,
    .I0 ( config1_decoder7.U17.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_11 ) ,
    .IN ( config1_decoder7.U17.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n74 ) ,
    .I0 ( config1_decoder7.n70 ) ,
    .I1 ( config1_decoder7.n79 ) ) ;
or ( 
    .Z ( config1_decoder7.U27.AB ) ,
    .I0 ( config1_decoder7.n89 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U27.ZN ) ,
    .I0 ( config1_decoder7.U27.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_83 ) ,
    .IN ( config1_decoder7.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U77.AB ) ,
    .I0 ( config1_decoder7.n86 ) ,
    .I1 ( config1_decoder7.n84 ) ) ;
and ( 
    .Z ( config1_decoder7.U77.ZN ) ,
    .I0 ( config1_decoder7.U77.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_19 ) ,
    .IN ( config1_decoder7.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U67.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U67.ZN ) ,
    .I0 ( config1_decoder7.U67.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_42 ) ,
    .IN ( config1_decoder7.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U10.AB ) ,
    .I0 ( config1_decoder7.n83 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U10.ZN ) ,
    .I0 ( config1_decoder7.U10.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_44 ) ,
    .IN ( config1_decoder7.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n91 ) ,
    .I0 ( config1_decoder7.n80 ) ,
    .I1 ( config1_decoder7.n78 ) ) ;
or ( 
    .Z ( config1_decoder7.U26.AB ) ,
    .I0 ( config1_decoder7.n90 ) ,
    .I1 ( config1_decoder7.n86 ) ) ;
and ( 
    .Z ( config1_decoder7.U26.ZN ) ,
    .I0 ( config1_decoder7.U26.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_84 ) ,
    .IN ( config1_decoder7.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U113.AB ) ,
    .I0 ( config1_decoder7.n93 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U113.ZN ) ,
    .I0 ( config1_decoder7.U113.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_82 ) ,
    .IN ( config1_decoder7.U113.ZN ) ) ;
nor ( 
    .Z ( config1_decoder7.n70 ) ,
    .I0 ( config1_decoder7.n69 ) ,
    .I1 ( masks_hold_reg_10_0 ) ) ;
nor ( 
    .Z ( config1_decoder7.n76 ) ,
    .I0 ( masks_hold_reg_12_7 ) ,
    .I1 ( masks_hold_reg_12_8 ) ) ;
nand ( 
    .Z ( config1_decoder7.n1 ) ,
    .I0 ( config1_decoder7.n94 ) ,
    .I1 ( config1_decoder7.n60 ) ) ;
nand ( 
    .Z ( config1_decoder7.n103 ) ,
    .I0 ( config1_decoder7.n67 ) ,
    .I1 ( config1_decoder7.n65 ) ,
    .I2 ( masks_hold_reg_12_10 ) ) ;
or ( 
    .Z ( config1_decoder7.U153.AB ) ,
    .I0 ( config1_decoder7.n95 ) ,
    .I1 ( config1_decoder7.n91 ) ) ;
and ( 
    .Z ( config1_decoder7.U153.ZN ) ,
    .I0 ( config1_decoder7.U153.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_65 ) ,
    .IN ( config1_decoder7.U153.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U141.AB ) ,
    .I0 ( config1_decoder7.n101 ) ,
    .I1 ( config1_decoder7.n96 ) ) ;
and ( 
    .Z ( config1_decoder7.U141.ZN ) ,
    .I0 ( config1_decoder7.U141.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_100 ) ,
    .IN ( config1_decoder7.U141.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U90.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U90.ZN ) ,
    .I0 ( config1_decoder7.U90.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_55 ) ,
    .IN ( config1_decoder7.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U3.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n85 ) ) ;
and ( 
    .Z ( config1_decoder7.U3.ZN ) ,
    .I0 ( config1_decoder7.U3.AB ) ,
    .I1 ( config1_decoder7.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_17 ) ,
    .IN ( config1_decoder7.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U86.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U86.ZN ) ,
    .I0 ( config1_decoder7.U86.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_60 ) ,
    .IN ( config1_decoder7.U86.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U58.AB ) ,
    .I0 ( config1_decoder7.n88 ) ,
    .I1 ( config1_decoder7.n74 ) ) ;
and ( 
    .Z ( config1_decoder7.U58.ZN ) ,
    .I0 ( config1_decoder7.U58.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_58 ) ,
    .IN ( config1_decoder7.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U46.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n88 ) ) ;
and ( 
    .Z ( config1_decoder7.U46.ZN ) ,
    .I0 ( config1_decoder7.U46.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_25 ) ,
    .IN ( config1_decoder7.U46.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U74.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n81 ) ) ;
and ( 
    .Z ( config1_decoder7.U74.ZN ) ,
    .I0 ( config1_decoder7.U74.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_30 ) ,
    .IN ( config1_decoder7.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U66.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U66.ZN ) ,
    .I0 ( config1_decoder7.U66.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_40 ) ,
    .IN ( config1_decoder7.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U11.AB ) ,
    .I0 ( config1_decoder7.n83 ) ,
    .I1 ( config1_decoder7.n71 ) ) ;
and ( 
    .Z ( config1_decoder7.U11.ZN ) ,
    .I0 ( config1_decoder7.U11.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_43 ) ,
    .IN ( config1_decoder7.U11.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n71 ) ,
    .I0 ( config1_decoder7.n70 ) ,
    .I1 ( config1_decoder7.n76 ) ) ;
nand ( 
    .Z ( config1_decoder7.n87 ) ,
    .I0 ( config1_decoder7.n77 ) ,
    .I1 ( config1_decoder7.n64 ) ) ;
or ( 
    .Z ( config1_decoder7.U112.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n89 ) ) ;
and ( 
    .Z ( config1_decoder7.U112.ZN ) ,
    .I0 ( config1_decoder7.U112.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_91 ) ,
    .IN ( config1_decoder7.U112.ZN ) ) ;
nand ( 
    .Z ( config1_decoder7.n97 ) ,
    .I0 ( masks_hold_reg_12_8 ) ,
    .I1 ( config1_decoder7.n62 ) ) ;
and ( 
    .Z ( config1_decoder7.U129.AB ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( config1_decoder7.n79 ) ) ;
or ( 
    .Z ( config1_decoder7.n60 ) ,
    .I0 ( config1_decoder7.U129.AB ) ,
    .I1 ( config1_decoder7.n68 ) ,
    .I2 ( masks_hold_reg_11_9 ) ) ;
nor ( 
    .Z ( config1_decoder7.n61 ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( masks_hold_reg_11_9 ) ) ;
or ( 
    .Z ( config1_decoder7.U152.AB ) ,
    .I0 ( config1_decoder7.n92 ) ,
    .I1 ( config1_decoder7.n73 ) ) ;
and ( 
    .Z ( config1_decoder7.U152.ZN ) ,
    .I0 ( config1_decoder7.U152.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_61 ) ,
    .IN ( config1_decoder7.U152.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U142.AB ) ,
    .I0 ( config1_decoder7.n101 ) ,
    .I1 ( config1_decoder7.n100 ) ) ;
and ( 
    .Z ( config1_decoder7.U142.ZN ) ,
    .I0 ( config1_decoder7.U142.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_99 ) ,
    .IN ( config1_decoder7.U142.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U162.AB ) ,
    .I0 ( config1_decoder7.n103 ) ,
    .I1 ( config1_decoder7.n90 ) ) ;
and ( 
    .Z ( config1_decoder7.U162.ZN ) ,
    .I0 ( config1_decoder7.U162.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_72 ) ,
    .IN ( config1_decoder7.U162.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U91.AB ) ,
    .I0 ( config1_decoder7.n85 ) ,
    .I1 ( config1_decoder7.n72 ) ) ;
and ( 
    .Z ( config1_decoder7.U91.ZN ) ,
    .I0 ( config1_decoder7.U91.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_48 ) ,
    .IN ( config1_decoder7.U91.ZN ) ) ;
or ( 
    .Z ( config1_decoder7.U2.AB ) ,
    .I0 ( config1_decoder7.n104 ) ,
    .I1 ( config1_decoder7.n95 ) ) ;
and ( 
    .Z ( config1_decoder7.U2.ZN ) ,
    .I0 ( config1_decoder7.U2.AB ) ,
    .I1 ( config1_decoder7.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_6_1 ) ,
    .IN ( config1_decoder7.U2.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder4.n2 ) ,
    .IN ( config1_decoder4.n1 ) ) ;
nand ( 
    .Z ( config1_decoder4.n103 ) ,
    .I0 ( config1_decoder4.n67 ) ,
    .I1 ( config1_decoder4.n65 ) ,
    .I2 ( masks_hold_reg_6_7 ) ) ;
or ( 
    .Z ( config1_decoder4.U113.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n89 ) ) ;
and ( 
    .Z ( config1_decoder4.U113.ZN ) ,
    .I0 ( config1_decoder4.U113.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_71 ) ,
    .IN ( config1_decoder4.U113.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n76 ) ,
    .I0 ( masks_hold_reg_6_4 ) ,
    .I1 ( masks_hold_reg_6_5 ) ) ;
nand ( 
    .Z ( config1_decoder4.n86 ) ,
    .I0 ( config1_decoder4.n66 ) ,
    .I1 ( masks_hold_reg_6_6 ) ) ;
nand ( 
    .Z ( config1_decoder4.n92 ) ,
    .I0 ( masks_hold_reg_6_8 ) ,
    .I1 ( config1_decoder4.n68 ) ) ;
or ( 
    .Z ( config1_decoder4.U125.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U125.ZN ) ,
    .I0 ( config1_decoder4.U125.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_62 ) ,
    .IN ( config1_decoder4.U125.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U153.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n82 ) ) ;
and ( 
    .Z ( config1_decoder4.U153.ZN ) ,
    .I0 ( config1_decoder4.U153.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_5 ) ,
    .IN ( config1_decoder4.U153.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n77 ) ,
    .I0 ( config1_decoder4.n62 ) ,
    .I1 ( masks_hold_reg_6_5 ) ) ;
or ( 
    .Z ( config1_decoder4.U90.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U90.ZN ) ,
    .I0 ( config1_decoder4.U90.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_27 ) ,
    .IN ( config1_decoder4.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U3.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U3.ZN ) ,
    .I0 ( config1_decoder4.U3.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_33 ) ,
    .IN ( config1_decoder4.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U86.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U86.ZN ) ,
    .I0 ( config1_decoder4.U86.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_49 ) ,
    .IN ( config1_decoder4.U86.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U58.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U58.ZN ) ,
    .I0 ( config1_decoder4.U58.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_38 ) ,
    .IN ( config1_decoder4.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U46.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n88 ) ) ;
and ( 
    .Z ( config1_decoder4.U46.ZN ) ,
    .I0 ( config1_decoder4.U46.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_25 ) ,
    .IN ( config1_decoder4.U46.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U74.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n87 ) ) ;
and ( 
    .Z ( config1_decoder4.U74.ZN ) ,
    .I0 ( config1_decoder4.U74.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_4 ) ,
    .IN ( config1_decoder4.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U66.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U66.ZN ) ,
    .I0 ( config1_decoder4.U66.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_22 ) ,
    .IN ( config1_decoder4.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U11.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U11.ZN ) ,
    .I0 ( config1_decoder4.U11.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_50 ) ,
    .IN ( config1_decoder4.U11.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U13.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U13.ZN ) ,
    .I0 ( config1_decoder4.U13.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_15 ) ,
    .IN ( config1_decoder4.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n91 ) ,
    .I0 ( config1_decoder4.n80 ) ,
    .I1 ( config1_decoder4.n78 ) ) ;
or ( 
    .Z ( config1_decoder4.U28.AB ) ,
    .I0 ( config1_decoder4.n89 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U28.ZN ) ,
    .I0 ( config1_decoder4.U28.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_75 ) ,
    .IN ( config1_decoder4.U28.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n67 ) ,
    .IN ( masks_hold_reg_6_6 ) ) ;
or ( 
    .Z ( config1_decoder4.U120.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n90 ) ) ;
and ( 
    .Z ( config1_decoder4.U120.ZN ) ,
    .I0 ( config1_decoder4.U120.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_64 ) ,
    .IN ( config1_decoder4.U120.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U154.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n95 ) ) ;
and ( 
    .Z ( config1_decoder4.U154.ZN ) ,
    .I0 ( config1_decoder4.U154.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_1 ) ,
    .IN ( config1_decoder4.U154.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n80 ) ,
    .I0 ( config1_decoder4.n75 ) ,
    .I1 ( masks_hold_reg_6_9 ) ) ;
or ( 
    .Z ( config1_decoder4.U160.AB ) ,
    .I0 ( config1_decoder4.n100 ) ,
    .I1 ( config1_decoder4.n98 ) ) ;
and ( 
    .Z ( config1_decoder4.U160.ZN ) ,
    .I0 ( config1_decoder4.U160.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_95 ) ,
    .IN ( config1_decoder4.U160.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n100 ) ,
    .IN ( config1_decoder4.n76 ) ) ;
or ( 
    .Z ( config1_decoder4.U83.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U83.ZN ) ,
    .I0 ( config1_decoder4.U83.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_55 ) ,
    .IN ( config1_decoder4.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U50.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U50.ZN ) ,
    .I0 ( config1_decoder4.U50.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_21 ) ,
    .IN ( config1_decoder4.U50.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n93 ) ,
    .I0 ( config1_decoder4.n80 ) ,
    .I1 ( config1_decoder4.n79 ) ) ;
or ( 
    .Z ( config1_decoder4.U121.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n93 ) ) ;
and ( 
    .Z ( config1_decoder4.U121.ZN ) ,
    .I0 ( config1_decoder4.U121.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_70 ) ,
    .IN ( config1_decoder4.U121.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U157.AB ) ,
    .I0 ( config1_decoder4.n101 ) ,
    .I1 ( config1_decoder4.n96 ) ) ;
and ( 
    .Z ( config1_decoder4.U157.ZN ) ,
    .I0 ( config1_decoder4.U157.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_100 ) ,
    .IN ( config1_decoder4.U157.ZN ) ) ;
and ( 
    .Z ( config1_decoder4.n68 ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( masks_hold_reg_6_6 ) ) ;
or ( 
    .Z ( config1_decoder4.U161.AB ) ,
    .I0 ( config1_decoder4.n93 ) ,
    .I1 ( config1_decoder4.n92 ) ) ;
and ( 
    .Z ( config1_decoder4.U161.ZN ) ,
    .I0 ( config1_decoder4.U161.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_94 ) ,
    .IN ( config1_decoder4.U161.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U82.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U82.ZN ) ,
    .I0 ( config1_decoder4.U82.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_56 ) ,
    .IN ( config1_decoder4.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U89.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U89.ZN ) ,
    .I0 ( config1_decoder4.U89.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_23 ) ,
    .IN ( config1_decoder4.U89.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U51.AB ) ,
    .I0 ( config1_decoder4.n87 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U51.ZN ) ,
    .I0 ( config1_decoder4.U51.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_20 ) ,
    .IN ( config1_decoder4.U51.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n84 ) ,
    .I0 ( config1_decoder4.n76 ) ,
    .I1 ( config1_decoder4.n64 ) ) ;
or ( 
    .Z ( config1_decoder4.U78.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U78.ZN ) ,
    .I0 ( config1_decoder4.U78.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_58 ) ,
    .IN ( config1_decoder4.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n89 ) ,
    .I0 ( config1_decoder4.n80 ) ,
    .I1 ( config1_decoder4.n76 ) ) ;
or ( 
    .Z ( config1_decoder4.U115.AB ) ,
    .I0 ( config1_decoder4.n93 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U115.ZN ) ,
    .I0 ( config1_decoder4.U115.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_86 ) ,
    .IN ( config1_decoder4.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U156.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U156.ZN ) ,
    .I0 ( config1_decoder4.U156.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_54 ) ,
    .IN ( config1_decoder4.U156.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n75 ) ,
    .IN ( masks_hold_reg_6_10 ) ) ;
or ( 
    .Z ( config1_decoder4.U5.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U5.ZN ) ,
    .I0 ( config1_decoder4.U5.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_34 ) ,
    .IN ( config1_decoder4.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U88.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n91 ) ) ;
and ( 
    .Z ( config1_decoder4.U88.ZN ) ,
    .I0 ( config1_decoder4.U88.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_73 ) ,
    .IN ( config1_decoder4.U88.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U52.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n87 ) ) ;
and ( 
    .Z ( config1_decoder4.U52.ZN ) ,
    .I0 ( config1_decoder4.U52.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_24 ) ,
    .IN ( config1_decoder4.U52.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n81 ) ,
    .I0 ( config1_decoder4.n79 ) ,
    .I1 ( config1_decoder4.n64 ) ) ;
or ( 
    .Z ( config1_decoder4.U79.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U79.ZN ) ,
    .I0 ( config1_decoder4.U79.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_60 ) ,
    .IN ( config1_decoder4.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U72.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U72.ZN ) ,
    .I0 ( config1_decoder4.U72.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_18 ) ,
    .IN ( config1_decoder4.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U69.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U69.ZN ) ,
    .I0 ( config1_decoder4.U69.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_30 ) ,
    .IN ( config1_decoder4.U69.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U119.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n90 ) ) ;
and ( 
    .Z ( config1_decoder4.U119.ZN ) ,
    .I0 ( config1_decoder4.U119.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_68 ) ,
    .IN ( config1_decoder4.U119.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n79 ) ,
    .IN ( config1_decoder4.n99 ) ) ;
or ( 
    .Z ( config1_decoder4.U2.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U2.ZN ) ,
    .I0 ( config1_decoder4.U2.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_17 ) ,
    .IN ( config1_decoder4.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U81.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U81.ZN ) ,
    .I0 ( config1_decoder4.U81.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_53 ) ,
    .IN ( config1_decoder4.U81.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U59.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U59.ZN ) ,
    .I0 ( config1_decoder4.U59.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_41 ) ,
    .IN ( config1_decoder4.U59.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.U49.BN ) ,
    .IN ( config1_decoder4.n103 ) ) ;
nand ( 
    .Z ( config1_decoder4.n63 ) ,
    .I0 ( config1_decoder4.U49.BN ) ,
    .I1 ( config1_decoder4.n94 ) ) ;
or ( 
    .Z ( config1_decoder4.U75.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U75.ZN ) ,
    .I0 ( config1_decoder4.U75.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_7 ) ,
    .IN ( config1_decoder4.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U65.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U65.ZN ) ,
    .I0 ( config1_decoder4.U65.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_26 ) ,
    .IN ( config1_decoder4.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U12.AB ) ,
    .I0 ( config1_decoder4.n83 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U12.ZN ) ,
    .I0 ( config1_decoder4.U12.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_14 ) ,
    .IN ( config1_decoder4.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n73 ) ,
    .I0 ( config1_decoder4.n70 ) ,
    .I1 ( config1_decoder4.n78 ) ) ;
nand ( 
    .Z ( config1_decoder4.n90 ) ,
    .I0 ( config1_decoder4.n80 ) ,
    .I1 ( config1_decoder4.n77 ) ) ;
nand ( 
    .Z ( config1_decoder4.n104 ) ,
    .I0 ( config1_decoder4.n64 ) ,
    .I1 ( config1_decoder4.n78 ) ) ;
or ( 
    .Z ( config1_decoder4.U103.AB ) ,
    .I0 ( config1_decoder4.n91 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U103.ZN ) ,
    .I0 ( config1_decoder4.U103.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_85 ) ,
    .IN ( config1_decoder4.U103.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U123.AB ) ,
    .I0 ( config1_decoder4.n90 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U123.ZN ) ,
    .I0 ( config1_decoder4.U123.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_80 ) ,
    .IN ( config1_decoder4.U123.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U155.AB ) ,
    .I0 ( config1_decoder4.n99 ) ,
    .I1 ( config1_decoder4.n98 ) ) ;
and ( 
    .Z ( config1_decoder4.U155.ZN ) ,
    .I0 ( config1_decoder4.U155.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_98 ) ,
    .IN ( config1_decoder4.U155.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n99 ) ,
    .I0 ( masks_hold_reg_6_4 ) ,
    .I1 ( masks_hold_reg_6_5 ) ) ;
or ( 
    .Z ( config1_decoder4.U163.AB ) ,
    .I0 ( config1_decoder4.n98 ) ,
    .I1 ( config1_decoder4.n96 ) ) ;
and ( 
    .Z ( config1_decoder4.U163.ZN ) ,
    .I0 ( config1_decoder4.U163.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_96 ) ,
    .IN ( config1_decoder4.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U92.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U92.ZN ) ,
    .I0 ( config1_decoder4.U92.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_19 ) ,
    .IN ( config1_decoder4.U92.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U80.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U80.ZN ) ,
    .I0 ( config1_decoder4.U80.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_59 ) ,
    .IN ( config1_decoder4.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U48.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n103 ) ) ;
and ( 
    .Z ( config1_decoder4.U48.ZN ) ,
    .I0 ( config1_decoder4.U48.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_9 ) ,
    .IN ( config1_decoder4.U48.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n78 ) ,
    .IN ( config1_decoder4.n97 ) ) ;
or ( 
    .Z ( config1_decoder4.U114.AB ) ,
    .I0 ( config1_decoder4.n93 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U114.ZN ) ,
    .I0 ( config1_decoder4.U114.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_82 ) ,
    .IN ( config1_decoder4.U114.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U104.AB ) ,
    .I0 ( config1_decoder4.n91 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U104.ZN ) ,
    .I0 ( config1_decoder4.U104.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_77 ) ,
    .IN ( config1_decoder4.U104.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U159.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U159.ZN ) ,
    .I0 ( config1_decoder4.U159.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_61 ) ,
    .IN ( config1_decoder4.U159.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n62 ) ,
    .IN ( masks_hold_reg_6_4 ) ) ;
or ( 
    .Z ( config1_decoder4.U9.AB ) ,
    .I0 ( config1_decoder4.n83 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U9.ZN ) ,
    .I0 ( config1_decoder4.U9.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_44 ) ,
    .IN ( config1_decoder4.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U4.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U4.ZN ) ,
    .I0 ( config1_decoder4.U4.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_32 ) ,
    .IN ( config1_decoder4.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U53.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n87 ) ) ;
and ( 
    .Z ( config1_decoder4.U53.ZN ) ,
    .I0 ( config1_decoder4.U53.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_8 ) ,
    .IN ( config1_decoder4.U53.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n95 ) ,
    .I0 ( config1_decoder4.n61 ) ,
    .I1 ( config1_decoder4.n67 ) ) ;
or ( 
    .Z ( config1_decoder4.U73.AB ) ,
    .I0 ( config1_decoder4.n90 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U73.ZN ) ,
    .I0 ( config1_decoder4.U73.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_76 ) ,
    .IN ( config1_decoder4.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U68.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n87 ) ) ;
and ( 
    .Z ( config1_decoder4.U68.ZN ) ,
    .I0 ( config1_decoder4.U68.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_28 ) ,
    .IN ( config1_decoder4.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U63.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U63.ZN ) ,
    .I0 ( config1_decoder4.U63.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_51 ) ,
    .IN ( config1_decoder4.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U14.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U14.ZN ) ,
    .I0 ( config1_decoder4.U14.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_13 ) ,
    .IN ( config1_decoder4.U14.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U118.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n93 ) ) ;
and ( 
    .Z ( config1_decoder4.U118.ZN ) ,
    .I0 ( config1_decoder4.U118.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_74 ) ,
    .IN ( config1_decoder4.U118.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U117.AB ) ,
    .I0 ( config1_decoder4.n93 ) ,
    .I1 ( config1_decoder4.n88 ) ) ;
and ( 
    .Z ( config1_decoder4.U117.ZN ) ,
    .I0 ( config1_decoder4.U117.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_90 ) ,
    .IN ( config1_decoder4.U117.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U108.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n91 ) ) ;
and ( 
    .Z ( config1_decoder4.U108.ZN ) ,
    .I0 ( config1_decoder4.U108.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_69 ) ,
    .IN ( config1_decoder4.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U105.AB ) ,
    .I0 ( config1_decoder4.n91 ) ,
    .I1 ( config1_decoder4.n88 ) ) ;
and ( 
    .Z ( config1_decoder4.U105.ZN ) ,
    .I0 ( config1_decoder4.U105.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_89 ) ,
    .IN ( config1_decoder4.U105.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n64 ) ,
    .I0 ( masks_hold_reg_6_9 ) ,
    .I1 ( masks_hold_reg_6_10 ) ) ;
or ( 
    .Z ( config1_decoder4.U158.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n91 ) ) ;
and ( 
    .Z ( config1_decoder4.U158.ZN ) ,
    .I0 ( config1_decoder4.U158.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_93 ) ,
    .IN ( config1_decoder4.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U148.AB ) ,
    .I0 ( config1_decoder4.n97 ) ,
    .I1 ( config1_decoder4.n98 ) ) ;
and ( 
    .Z ( config1_decoder4.U148.ZN ) ,
    .I0 ( config1_decoder4.U148.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_97 ) ,
    .IN ( config1_decoder4.U148.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U164.AB ) ,
    .I0 ( config1_decoder4.n97 ) ,
    .I1 ( config1_decoder4.n63 ) ) ;
and ( 
    .Z ( config1_decoder4.U164.ZN ) ,
    .I0 ( config1_decoder4.U164.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_105 ) ,
    .IN ( config1_decoder4.U164.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n96 ) ,
    .IN ( config1_decoder4.n77 ) ) ;
or ( 
    .Z ( config1_decoder4.U8.AB ) ,
    .I0 ( config1_decoder4.n83 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U8.ZN ) ,
    .I0 ( config1_decoder4.U8.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_45 ) ,
    .IN ( config1_decoder4.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U7.AB ) ,
    .I0 ( config1_decoder4.n83 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U7.ZN ) ,
    .I0 ( config1_decoder4.U7.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_46 ) ,
    .IN ( config1_decoder4.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U54.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U54.ZN ) ,
    .I0 ( config1_decoder4.U54.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_35 ) ,
    .IN ( config1_decoder4.U54.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n94 ) ,
    .I0 ( config1_decoder4.n75 ) ,
    .I1 ( config1_decoder4.n69 ) ) ;
or ( 
    .Z ( config1_decoder4.U70.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U70.ZN ) ,
    .I0 ( config1_decoder4.U70.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_31 ) ,
    .IN ( config1_decoder4.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U62.AB ) ,
    .I0 ( config1_decoder4.n86 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U62.ZN ) ,
    .I0 ( config1_decoder4.U62.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_52 ) ,
    .IN ( config1_decoder4.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U15.AB ) ,
    .I0 ( config1_decoder4.n87 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U15.ZN ) ,
    .I0 ( config1_decoder4.U15.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_12 ) ,
    .IN ( config1_decoder4.U15.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U116.AB ) ,
    .I0 ( config1_decoder4.n93 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U116.ZN ) ,
    .I0 ( config1_decoder4.U116.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_78 ) ,
    .IN ( config1_decoder4.U116.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U109.AB ) ,
    .I0 ( config1_decoder4.n89 ) ,
    .I1 ( config1_decoder4.n88 ) ) ;
and ( 
    .Z ( config1_decoder4.U109.ZN ) ,
    .I0 ( config1_decoder4.U109.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_87 ) ,
    .IN ( config1_decoder4.U109.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U106.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n89 ) ) ;
and ( 
    .Z ( config1_decoder4.U106.ZN ) ,
    .I0 ( config1_decoder4.U106.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_67 ) ,
    .IN ( config1_decoder4.U106.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.n65 ) ,
    .IN ( masks_hold_reg_6_8 ) ) ;
or ( 
    .Z ( config1_decoder4.U126.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n93 ) ) ;
and ( 
    .Z ( config1_decoder4.U126.ZN ) ,
    .I0 ( config1_decoder4.U126.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_66 ) ,
    .IN ( config1_decoder4.U126.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U149.AB ) ,
    .I0 ( config1_decoder4.n101 ) ,
    .I1 ( config1_decoder4.n100 ) ) ;
and ( 
    .Z ( config1_decoder4.U149.ZN ) ,
    .I0 ( config1_decoder4.U149.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_99 ) ,
    .IN ( config1_decoder4.U149.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U165.AB ) ,
    .I0 ( config1_decoder4.n100 ) ,
    .I1 ( config1_decoder4.n63 ) ) ;
and ( 
    .Z ( config1_decoder4.U165.ZN ) ,
    .I0 ( config1_decoder4.U165.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_103 ) ,
    .IN ( config1_decoder4.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U95.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U95.ZN ) ,
    .I0 ( config1_decoder4.U95.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_6 ) ,
    .IN ( config1_decoder4.U95.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U6.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U6.ZN ) ,
    .I0 ( config1_decoder4.U6.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_47 ) ,
    .IN ( config1_decoder4.U6.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U85.AB ) ,
    .I0 ( config1_decoder4.n97 ) ,
    .I1 ( config1_decoder4.n101 ) ) ;
and ( 
    .Z ( config1_decoder4.U85.ZN ) ,
    .I0 ( config1_decoder4.U85.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_101 ) ,
    .IN ( config1_decoder4.U85.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U55.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U55.ZN ) ,
    .I0 ( config1_decoder4.U55.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_39 ) ,
    .IN ( config1_decoder4.U55.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n83 ) ,
    .I0 ( config1_decoder4.n68 ) ,
    .I1 ( config1_decoder4.n65 ) ) ;
or ( 
    .Z ( config1_decoder4.U71.AB ) ,
    .I0 ( config1_decoder4.n87 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U71.ZN ) ,
    .I0 ( config1_decoder4.U71.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_16 ) ,
    .IN ( config1_decoder4.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U61.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n74 ) ) ;
and ( 
    .Z ( config1_decoder4.U61.ZN ) ,
    .I0 ( config1_decoder4.U61.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_42 ) ,
    .IN ( config1_decoder4.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U16.AB ) ,
    .I0 ( config1_decoder4.n84 ) ,
    .I1 ( config1_decoder4.n83 ) ) ;
and ( 
    .Z ( config1_decoder4.U16.ZN ) ,
    .I0 ( config1_decoder4.U16.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_11 ) ,
    .IN ( config1_decoder4.U16.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n74 ) ,
    .I0 ( config1_decoder4.n70 ) ,
    .I1 ( config1_decoder4.n79 ) ) ;
or ( 
    .Z ( config1_decoder4.U111.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n89 ) ) ;
and ( 
    .Z ( config1_decoder4.U111.ZN ) ,
    .I0 ( config1_decoder4.U111.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_91 ) ,
    .IN ( config1_decoder4.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U107.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n89 ) ) ;
and ( 
    .Z ( config1_decoder4.U107.ZN ) ,
    .I0 ( config1_decoder4.U107.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_63 ) ,
    .IN ( config1_decoder4.U107.ZN ) ) ;
and ( 
    .Z ( config1_decoder4.U135.AB ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( config1_decoder4.n79 ) ) ;
or ( 
    .Z ( config1_decoder4.n60 ) ,
    .I0 ( config1_decoder4.U135.AB ) ,
    .I1 ( config1_decoder4.n68 ) ,
    .I2 ( masks_hold_reg_6_8 ) ) ;
nand ( 
    .Z ( config1_decoder4.n88 ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( config1_decoder4.n67 ) ,
    .I2 ( masks_hold_reg_6_8 ) ) ;
not ( 
    .O1 ( config1_decoder4.n69 ) ,
    .IN ( masks_hold_reg_6_9 ) ) ;
or ( 
    .Z ( config1_decoder4.U96.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n84 ) ) ;
and ( 
    .Z ( config1_decoder4.U96.ZN ) ,
    .I0 ( config1_decoder4.U96.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_3 ) ,
    .IN ( config1_decoder4.U96.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.U1.BN ) ,
    .IN ( config1_decoder4.n95 ) ) ;
nand ( 
    .Z ( config1_decoder4.n98 ) ,
    .I0 ( config1_decoder4.U1.BN ) ,
    .I1 ( config1_decoder4.n94 ) ) ;
or ( 
    .Z ( config1_decoder4.U84.AB ) ,
    .I0 ( config1_decoder4.n85 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U84.ZN ) ,
    .I0 ( config1_decoder4.U84.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_48 ) ,
    .IN ( config1_decoder4.U84.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U56.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U56.ZN ) ,
    .I0 ( config1_decoder4.U56.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_37 ) ,
    .IN ( config1_decoder4.U56.ZN ) ) ;
not ( 
    .O1 ( config1_decoder4.U44.BN ) ,
    .IN ( config1_decoder4.n82 ) ) ;
nand ( 
    .Z ( config1_decoder4.n101 ) ,
    .I0 ( config1_decoder4.U44.BN ) ,
    .I1 ( config1_decoder4.n94 ) ) ;
or ( 
    .Z ( config1_decoder4.U76.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n87 ) ) ;
and ( 
    .Z ( config1_decoder4.U76.ZN ) ,
    .I0 ( config1_decoder4.U76.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_0 ) ,
    .IN ( config1_decoder4.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U60.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U60.ZN ) ,
    .I0 ( config1_decoder4.U60.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_40 ) ,
    .IN ( config1_decoder4.U60.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n71 ) ,
    .I0 ( config1_decoder4.n70 ) ,
    .I1 ( config1_decoder4.n76 ) ) ;
or ( 
    .Z ( config1_decoder4.U27.AB ) ,
    .I0 ( config1_decoder4.n89 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U27.ZN ) ,
    .I0 ( config1_decoder4.U27.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_83 ) ,
    .IN ( config1_decoder4.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U110.AB ) ,
    .I0 ( config1_decoder4.n89 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U110.ZN ) ,
    .I0 ( config1_decoder4.U110.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_79 ) ,
    .IN ( config1_decoder4.U110.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n66 ) ,
    .I0 ( config1_decoder4.n65 ) ,
    .I1 ( masks_hold_reg_6_7 ) ) ;
nand ( 
    .Z ( config1_decoder4.n1 ) ,
    .I0 ( config1_decoder4.n94 ) ,
    .I1 ( config1_decoder4.n60 ) ) ;
or ( 
    .Z ( config1_decoder4.U124.AB ) ,
    .I0 ( config1_decoder4.n92 ) ,
    .I1 ( config1_decoder4.n90 ) ) ;
and ( 
    .Z ( config1_decoder4.U124.ZN ) ,
    .I0 ( config1_decoder4.U124.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_92 ) ,
    .IN ( config1_decoder4.U124.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U150.AB ) ,
    .I0 ( config1_decoder4.n96 ) ,
    .I1 ( config1_decoder4.n63 ) ) ;
and ( 
    .Z ( config1_decoder4.U150.ZN ) ,
    .I0 ( config1_decoder4.U150.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_104 ) ,
    .IN ( config1_decoder4.U150.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n97 ) ,
    .I0 ( masks_hold_reg_6_5 ) ,
    .I1 ( config1_decoder4.n62 ) ) ;
or ( 
    .Z ( config1_decoder4.U87.AB ) ,
    .I0 ( config1_decoder4.n99 ) ,
    .I1 ( config1_decoder4.n101 ) ) ;
and ( 
    .Z ( config1_decoder4.U87.ZN ) ,
    .I0 ( config1_decoder4.U87.AB ) ,
    .I1 ( config1_decoder4.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_102 ) ,
    .IN ( config1_decoder4.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U57.AB ) ,
    .I0 ( config1_decoder4.n82 ) ,
    .I1 ( config1_decoder4.n72 ) ) ;
and ( 
    .Z ( config1_decoder4.U57.ZN ) ,
    .I0 ( config1_decoder4.U57.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_36 ) ,
    .IN ( config1_decoder4.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U47.AB ) ,
    .I0 ( config1_decoder4.n104 ) ,
    .I1 ( config1_decoder4.n92 ) ) ;
and ( 
    .Z ( config1_decoder4.U47.ZN ) ,
    .I0 ( config1_decoder4.U47.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_29 ) ,
    .IN ( config1_decoder4.U47.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U77.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U77.ZN ) ,
    .I0 ( config1_decoder4.U77.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_2 ) ,
    .IN ( config1_decoder4.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U67.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n81 ) ) ;
and ( 
    .Z ( config1_decoder4.U67.ZN ) ,
    .I0 ( config1_decoder4.U67.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_10 ) ,
    .IN ( config1_decoder4.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U10.AB ) ,
    .I0 ( config1_decoder4.n83 ) ,
    .I1 ( config1_decoder4.n71 ) ) ;
and ( 
    .Z ( config1_decoder4.U10.ZN ) ,
    .I0 ( config1_decoder4.U10.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_43 ) ,
    .IN ( config1_decoder4.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n87 ) ,
    .I0 ( config1_decoder4.n77 ) ,
    .I1 ( config1_decoder4.n64 ) ) ;
or ( 
    .Z ( config1_decoder4.U26.AB ) ,
    .I0 ( config1_decoder4.n90 ) ,
    .I1 ( config1_decoder4.n86 ) ) ;
and ( 
    .Z ( config1_decoder4.U26.ZN ) ,
    .I0 ( config1_decoder4.U26.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_84 ) ,
    .IN ( config1_decoder4.U26.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n72 ) ,
    .I0 ( config1_decoder4.n70 ) ,
    .I1 ( config1_decoder4.n77 ) ) ;
nand ( 
    .Z ( config1_decoder4.n85 ) ,
    .I0 ( config1_decoder4.n66 ) ,
    .I1 ( config1_decoder4.n67 ) ) ;
or ( 
    .Z ( config1_decoder4.U25.AB ) ,
    .I0 ( config1_decoder4.n91 ) ,
    .I1 ( config1_decoder4.n85 ) ) ;
and ( 
    .Z ( config1_decoder4.U25.ZN ) ,
    .I0 ( config1_decoder4.U25.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_81 ) ,
    .IN ( config1_decoder4.U25.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U112.AB ) ,
    .I0 ( config1_decoder4.n95 ) ,
    .I1 ( config1_decoder4.n91 ) ) ;
and ( 
    .Z ( config1_decoder4.U112.ZN ) ,
    .I0 ( config1_decoder4.U112.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_65 ) ,
    .IN ( config1_decoder4.U112.ZN ) ) ;
nand ( 
    .Z ( config1_decoder4.n82 ) ,
    .I0 ( config1_decoder4.n61 ) ,
    .I1 ( masks_hold_reg_6_6 ) ) ;
nor ( 
    .Z ( config1_decoder4.n61 ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( masks_hold_reg_6_8 ) ) ;
or ( 
    .Z ( config1_decoder4.U122.AB ) ,
    .I0 ( config1_decoder4.n90 ) ,
    .I1 ( config1_decoder4.n88 ) ) ;
and ( 
    .Z ( config1_decoder4.U122.ZN ) ,
    .I0 ( config1_decoder4.U122.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_88 ) ,
    .IN ( config1_decoder4.U122.ZN ) ) ;
or ( 
    .Z ( config1_decoder4.U152.AB ) ,
    .I0 ( config1_decoder4.n88 ) ,
    .I1 ( config1_decoder4.n73 ) ) ;
and ( 
    .Z ( config1_decoder4.U152.ZN ) ,
    .I0 ( config1_decoder4.U152.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_57 ) ,
    .IN ( config1_decoder4.U152.ZN ) ) ;
nor ( 
    .Z ( config1_decoder4.n70 ) ,
    .I0 ( config1_decoder4.n69 ) ,
    .I1 ( masks_hold_reg_6_10 ) ) ;
or ( 
    .Z ( config1_decoder4.U162.AB ) ,
    .I0 ( config1_decoder4.n103 ) ,
    .I1 ( config1_decoder4.n90 ) ) ;
and ( 
    .Z ( config1_decoder4.U162.ZN ) ,
    .I0 ( config1_decoder4.U162.AB ) ,
    .I1 ( config1_decoder4.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_3_72 ) ,
    .IN ( config1_decoder4.U162.ZN ) ) ;
buf ( 
    .O1 ( config1_decoder5.n2 ) ,
    .IN ( config1_decoder5.n1 ) ) ;
nand ( 
    .Z ( config1_decoder5.n97 ) ,
    .I0 ( masks_hold_reg_8_6 ) ,
    .I1 ( config1_decoder5.n62 ) ) ;
nand ( 
    .Z ( config1_decoder5.n103 ) ,
    .I0 ( config1_decoder5.n67 ) ,
    .I1 ( config1_decoder5.n65 ) ,
    .I2 ( masks_hold_reg_8_8 ) ) ;
or ( 
    .Z ( config1_decoder5.U152.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n89 ) ) ;
and ( 
    .Z ( config1_decoder5.U152.ZN ) ,
    .I0 ( config1_decoder5.U152.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_71 ) ,
    .IN ( config1_decoder5.U152.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U142.AB ) ,
    .I0 ( config1_decoder5.n97 ) ,
    .I1 ( config1_decoder5.n98 ) ) ;
and ( 
    .Z ( config1_decoder5.U142.ZN ) ,
    .I0 ( config1_decoder5.U142.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_97 ) ,
    .IN ( config1_decoder5.U142.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U162.AB ) ,
    .I0 ( config1_decoder5.n98 ) ,
    .I1 ( config1_decoder5.n96 ) ) ;
and ( 
    .Z ( config1_decoder5.U162.ZN ) ,
    .I0 ( config1_decoder5.U162.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_96 ) ,
    .IN ( config1_decoder5.U162.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U91.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U91.ZN ) ,
    .I0 ( config1_decoder5.U91.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_55 ) ,
    .IN ( config1_decoder5.U91.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U2.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U2.ZN ) ,
    .I0 ( config1_decoder5.U2.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_17 ) ,
    .IN ( config1_decoder5.U2.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U81.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U81.ZN ) ,
    .I0 ( config1_decoder5.U81.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_7 ) ,
    .IN ( config1_decoder5.U81.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U59.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U59.ZN ) ,
    .I0 ( config1_decoder5.U59.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_37 ) ,
    .IN ( config1_decoder5.U59.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U49.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n103 ) ) ;
and ( 
    .Z ( config1_decoder5.U49.ZN ) ,
    .I0 ( config1_decoder5.U49.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_9 ) ,
    .IN ( config1_decoder5.U49.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U75.AB ) ,
    .I0 ( config1_decoder5.n87 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U75.ZN ) ,
    .I0 ( config1_decoder5.U75.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_16 ) ,
    .IN ( config1_decoder5.U75.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U65.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U65.ZN ) ,
    .I0 ( config1_decoder5.U65.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_58 ) ,
    .IN ( config1_decoder5.U65.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U12.AB ) ,
    .I0 ( config1_decoder5.n83 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U12.ZN ) ,
    .I0 ( config1_decoder5.U12.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_14 ) ,
    .IN ( config1_decoder5.U12.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n73 ) ,
    .I0 ( config1_decoder5.n70 ) ,
    .I1 ( config1_decoder5.n78 ) ) ;
nand ( 
    .Z ( config1_decoder5.n90 ) ,
    .I0 ( config1_decoder5.n80 ) ,
    .I1 ( config1_decoder5.n77 ) ) ;
or ( 
    .Z ( config1_decoder5.U13.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U13.ZN ) ,
    .I0 ( config1_decoder5.U13.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_15 ) ,
    .IN ( config1_decoder5.U13.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n91 ) ,
    .I0 ( config1_decoder5.n80 ) ,
    .I1 ( config1_decoder5.n78 ) ) ;
or ( 
    .Z ( config1_decoder5.U28.AB ) ,
    .I0 ( config1_decoder5.n89 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U28.ZN ) ,
    .I0 ( config1_decoder5.U28.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_83 ) ,
    .IN ( config1_decoder5.U28.ZN ) ) ;
nor ( 
    .Z ( config1_decoder5.n77 ) ,
    .I0 ( config1_decoder5.n62 ) ,
    .I1 ( masks_hold_reg_8_6 ) ) ;
not ( 
    .O1 ( config1_decoder5.n67 ) ,
    .IN ( masks_hold_reg_8_7 ) ) ;
or ( 
    .Z ( config1_decoder5.U154.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n90 ) ) ;
and ( 
    .Z ( config1_decoder5.U154.ZN ) ,
    .I0 ( config1_decoder5.U154.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_68 ) ,
    .IN ( config1_decoder5.U154.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U144.AB ) ,
    .I0 ( config1_decoder5.n91 ) ,
    .I1 ( config1_decoder5.n88 ) ) ;
and ( 
    .Z ( config1_decoder5.U144.ZN ) ,
    .I0 ( config1_decoder5.U144.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_89 ) ,
    .IN ( config1_decoder5.U144.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U160.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n93 ) ) ;
and ( 
    .Z ( config1_decoder5.U160.ZN ) ,
    .I0 ( config1_decoder5.U160.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_66 ) ,
    .IN ( config1_decoder5.U160.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U93.AB ) ,
    .I0 ( config1_decoder5.n97 ) ,
    .I1 ( config1_decoder5.n101 ) ) ;
and ( 
    .Z ( config1_decoder5.U93.ZN ) ,
    .I0 ( config1_decoder5.U93.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_101 ) ,
    .IN ( config1_decoder5.U93.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U98.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U98.ZN ) ,
    .I0 ( config1_decoder5.U98.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_27 ) ,
    .IN ( config1_decoder5.U98.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U83.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n87 ) ) ;
and ( 
    .Z ( config1_decoder5.U83.ZN ) ,
    .I0 ( config1_decoder5.U83.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_0 ) ,
    .IN ( config1_decoder5.U83.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U50.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U50.ZN ) ,
    .I0 ( config1_decoder5.U50.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_21 ) ,
    .IN ( config1_decoder5.U50.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n93 ) ,
    .I0 ( config1_decoder5.n80 ) ,
    .I1 ( config1_decoder5.n79 ) ) ;
nand ( 
    .Z ( config1_decoder5.n82 ) ,
    .I0 ( config1_decoder5.n61 ) ,
    .I1 ( masks_hold_reg_8_7 ) ) ;
or ( 
    .Z ( config1_decoder5.U157.AB ) ,
    .I0 ( config1_decoder5.n93 ) ,
    .I1 ( config1_decoder5.n92 ) ) ;
and ( 
    .Z ( config1_decoder5.U157.ZN ) ,
    .I0 ( config1_decoder5.U157.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_94 ) ,
    .IN ( config1_decoder5.U157.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U145.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n89 ) ) ;
and ( 
    .Z ( config1_decoder5.U145.ZN ) ,
    .I0 ( config1_decoder5.U145.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_67 ) ,
    .IN ( config1_decoder5.U145.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U161.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n90 ) ) ;
and ( 
    .Z ( config1_decoder5.U161.ZN ) ,
    .I0 ( config1_decoder5.U161.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_72 ) ,
    .IN ( config1_decoder5.U161.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n100 ) ,
    .IN ( config1_decoder5.n76 ) ) ;
or ( 
    .Z ( config1_decoder5.U82.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U82.ZN ) ,
    .I0 ( config1_decoder5.U82.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_6 ) ,
    .IN ( config1_decoder5.U82.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U89.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U89.ZN ) ,
    .I0 ( config1_decoder5.U89.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_53 ) ,
    .IN ( config1_decoder5.U89.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U51.AB ) ,
    .I0 ( config1_decoder5.n87 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U51.ZN ) ,
    .I0 ( config1_decoder5.U51.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_20 ) ,
    .IN ( config1_decoder5.U51.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n84 ) ,
    .I0 ( config1_decoder5.n76 ) ,
    .I1 ( config1_decoder5.n64 ) ) ;
or ( 
    .Z ( config1_decoder5.U78.AB ) ,
    .I0 ( config1_decoder5.n89 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U78.ZN ) ,
    .I0 ( config1_decoder5.U78.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_75 ) ,
    .IN ( config1_decoder5.U78.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n89 ) ,
    .I0 ( config1_decoder5.n80 ) ,
    .I1 ( config1_decoder5.n76 ) ) ;
or ( 
    .Z ( config1_decoder5.U115.AB ) ,
    .I0 ( config1_decoder5.n90 ) ,
    .I1 ( config1_decoder5.n88 ) ) ;
and ( 
    .Z ( config1_decoder5.U115.ZN ) ,
    .I0 ( config1_decoder5.U115.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_88 ) ,
    .IN ( config1_decoder5.U115.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U156.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n93 ) ) ;
and ( 
    .Z ( config1_decoder5.U156.ZN ) ,
    .I0 ( config1_decoder5.U156.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_70 ) ,
    .IN ( config1_decoder5.U156.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U146.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n89 ) ) ;
and ( 
    .Z ( config1_decoder5.U146.ZN ) ,
    .I0 ( config1_decoder5.U146.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_63 ) ,
    .IN ( config1_decoder5.U146.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U5.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U5.ZN ) ,
    .I0 ( config1_decoder5.U5.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_34 ) ,
    .IN ( config1_decoder5.U5.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U88.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U88.ZN ) ,
    .I0 ( config1_decoder5.U88.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_59 ) ,
    .IN ( config1_decoder5.U88.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.U52.BN ) ,
    .IN ( config1_decoder5.n103 ) ) ;
nand ( 
    .Z ( config1_decoder5.n63 ) ,
    .I0 ( config1_decoder5.U52.BN ) ,
    .I1 ( config1_decoder5.n94 ) ) ;
nand ( 
    .Z ( config1_decoder5.n81 ) ,
    .I0 ( config1_decoder5.n79 ) ,
    .I1 ( config1_decoder5.n64 ) ) ;
or ( 
    .Z ( config1_decoder5.U79.AB ) ,
    .I0 ( config1_decoder5.n90 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U79.ZN ) ,
    .I0 ( config1_decoder5.U79.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_76 ) ,
    .IN ( config1_decoder5.U79.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U72.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n87 ) ) ;
and ( 
    .Z ( config1_decoder5.U72.ZN ) ,
    .I0 ( config1_decoder5.U72.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_28 ) ,
    .IN ( config1_decoder5.U72.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U69.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U69.ZN ) ,
    .I0 ( config1_decoder5.U69.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_26 ) ,
    .IN ( config1_decoder5.U69.ZN ) ) ;
nor ( 
    .Z ( config1_decoder5.n61 ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( masks_hold_reg_8_9 ) ) ;
or ( 
    .Z ( config1_decoder5.U114.AB ) ,
    .I0 ( config1_decoder5.n93 ) ,
    .I1 ( config1_decoder5.n88 ) ) ;
and ( 
    .Z ( config1_decoder5.U114.ZN ) ,
    .I0 ( config1_decoder5.U114.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_90 ) ,
    .IN ( config1_decoder5.U114.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U159.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U159.ZN ) ,
    .I0 ( config1_decoder5.U159.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_62 ) ,
    .IN ( config1_decoder5.U159.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U147.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n91 ) ) ;
and ( 
    .Z ( config1_decoder5.U147.ZN ) ,
    .I0 ( config1_decoder5.U147.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_69 ) ,
    .IN ( config1_decoder5.U147.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U9.AB ) ,
    .I0 ( config1_decoder5.n83 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U9.ZN ) ,
    .I0 ( config1_decoder5.U9.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_44 ) ,
    .IN ( config1_decoder5.U9.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U4.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U4.ZN ) ,
    .I0 ( config1_decoder5.U4.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_32 ) ,
    .IN ( config1_decoder5.U4.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U53.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n87 ) ) ;
and ( 
    .Z ( config1_decoder5.U53.ZN ) ,
    .I0 ( config1_decoder5.U53.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_24 ) ,
    .IN ( config1_decoder5.U53.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n95 ) ,
    .I0 ( config1_decoder5.n61 ) ,
    .I1 ( config1_decoder5.n67 ) ) ;
or ( 
    .Z ( config1_decoder5.U73.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U73.ZN ) ,
    .I0 ( config1_decoder5.U73.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_30 ) ,
    .IN ( config1_decoder5.U73.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U68.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U68.ZN ) ,
    .I0 ( config1_decoder5.U68.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_51 ) ,
    .IN ( config1_decoder5.U68.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U63.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U63.ZN ) ,
    .I0 ( config1_decoder5.U63.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_40 ) ,
    .IN ( config1_decoder5.U63.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U14.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U14.ZN ) ,
    .I0 ( config1_decoder5.U14.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_13 ) ,
    .IN ( config1_decoder5.U14.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n92 ) ,
    .I0 ( masks_hold_reg_8_9 ) ,
    .I1 ( config1_decoder5.n68 ) ) ;
nand ( 
    .Z ( config1_decoder5.n88 ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( config1_decoder5.n67 ) ,
    .I2 ( masks_hold_reg_8_9 ) ) ;
or ( 
    .Z ( config1_decoder5.U108.AB ) ,
    .I0 ( config1_decoder5.n91 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U108.ZN ) ,
    .I0 ( config1_decoder5.U108.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_85 ) ,
    .IN ( config1_decoder5.U108.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U137.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n93 ) ) ;
and ( 
    .Z ( config1_decoder5.U137.ZN ) ,
    .I0 ( config1_decoder5.U137.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_74 ) ,
    .IN ( config1_decoder5.U137.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U158.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n90 ) ) ;
and ( 
    .Z ( config1_decoder5.U158.ZN ) ,
    .I0 ( config1_decoder5.U158.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_92 ) ,
    .IN ( config1_decoder5.U158.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U148.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n91 ) ) ;
and ( 
    .Z ( config1_decoder5.U148.ZN ) ,
    .I0 ( config1_decoder5.U148.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_93 ) ,
    .IN ( config1_decoder5.U148.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U164.AB ) ,
    .I0 ( config1_decoder5.n97 ) ,
    .I1 ( config1_decoder5.n63 ) ) ;
and ( 
    .Z ( config1_decoder5.U164.ZN ) ,
    .I0 ( config1_decoder5.U164.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_105 ) ,
    .IN ( config1_decoder5.U164.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U94.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U94.ZN ) ,
    .I0 ( config1_decoder5.U94.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_49 ) ,
    .IN ( config1_decoder5.U94.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n104 ) ,
    .I0 ( config1_decoder5.n64 ) ,
    .I1 ( config1_decoder5.n78 ) ) ;
nand ( 
    .Z ( config1_decoder5.n99 ) ,
    .I0 ( masks_hold_reg_8_5 ) ,
    .I1 ( masks_hold_reg_8_6 ) ) ;
nand ( 
    .Z ( config1_decoder5.n86 ) ,
    .I0 ( config1_decoder5.n66 ) ,
    .I1 ( masks_hold_reg_8_7 ) ) ;
or ( 
    .Z ( config1_decoder5.U155.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n90 ) ) ;
and ( 
    .Z ( config1_decoder5.U155.ZN ) ,
    .I0 ( config1_decoder5.U155.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_64 ) ,
    .IN ( config1_decoder5.U155.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U143.AB ) ,
    .I0 ( config1_decoder5.n101 ) ,
    .I1 ( config1_decoder5.n96 ) ) ;
and ( 
    .Z ( config1_decoder5.U143.ZN ) ,
    .I0 ( config1_decoder5.U143.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_100 ) ,
    .IN ( config1_decoder5.U143.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U163.AB ) ,
    .I0 ( config1_decoder5.n96 ) ,
    .I1 ( config1_decoder5.n63 ) ) ;
and ( 
    .Z ( config1_decoder5.U163.ZN ) ,
    .I0 ( config1_decoder5.U163.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_104 ) ,
    .IN ( config1_decoder5.U163.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U92.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U92.ZN ) ,
    .I0 ( config1_decoder5.U92.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_48 ) ,
    .IN ( config1_decoder5.U92.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U80.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n87 ) ) ;
and ( 
    .Z ( config1_decoder5.U80.ZN ) ,
    .I0 ( config1_decoder5.U80.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_4 ) ,
    .IN ( config1_decoder5.U80.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U48.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n82 ) ) ;
and ( 
    .Z ( config1_decoder5.U48.ZN ) ,
    .I0 ( config1_decoder5.U48.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_5 ) ,
    .IN ( config1_decoder5.U48.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U64.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U64.ZN ) ,
    .I0 ( config1_decoder5.U64.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_42 ) ,
    .IN ( config1_decoder5.U64.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U8.AB ) ,
    .I0 ( config1_decoder5.n83 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U8.ZN ) ,
    .I0 ( config1_decoder5.U8.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_45 ) ,
    .IN ( config1_decoder5.U8.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U7.AB ) ,
    .I0 ( config1_decoder5.n83 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U7.ZN ) ,
    .I0 ( config1_decoder5.U7.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_46 ) ,
    .IN ( config1_decoder5.U7.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U54.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n87 ) ) ;
and ( 
    .Z ( config1_decoder5.U54.ZN ) ,
    .I0 ( config1_decoder5.U54.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_8 ) ,
    .IN ( config1_decoder5.U54.ZN ) ) ;
nor ( 
    .Z ( config1_decoder5.n94 ) ,
    .I0 ( config1_decoder5.n75 ) ,
    .I1 ( config1_decoder5.n69 ) ) ;
or ( 
    .Z ( config1_decoder5.U70.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U70.ZN ) ,
    .I0 ( config1_decoder5.U70.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_22 ) ,
    .IN ( config1_decoder5.U70.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U62.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U62.ZN ) ,
    .I0 ( config1_decoder5.U62.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_41 ) ,
    .IN ( config1_decoder5.U62.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U15.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n95 ) ) ;
and ( 
    .Z ( config1_decoder5.U15.ZN ) ,
    .I0 ( config1_decoder5.U15.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_1 ) ,
    .IN ( config1_decoder5.U15.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U116.AB ) ,
    .I0 ( config1_decoder5.n90 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U116.ZN ) ,
    .I0 ( config1_decoder5.U116.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_80 ) ,
    .IN ( config1_decoder5.U116.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U109.AB ) ,
    .I0 ( config1_decoder5.n89 ) ,
    .I1 ( config1_decoder5.n88 ) ) ;
and ( 
    .Z ( config1_decoder5.U109.ZN ) ,
    .I0 ( config1_decoder5.U109.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_87 ) ,
    .IN ( config1_decoder5.U109.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n62 ) ,
    .IN ( masks_hold_reg_8_5 ) ) ;
and ( 
    .Z ( config1_decoder5.U126.AB ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( config1_decoder5.n79 ) ) ;
or ( 
    .Z ( config1_decoder5.n60 ) ,
    .I0 ( config1_decoder5.U126.AB ) ,
    .I1 ( config1_decoder5.n68 ) ,
    .I2 ( masks_hold_reg_8_9 ) ) ;
or ( 
    .Z ( config1_decoder5.U149.AB ) ,
    .I0 ( config1_decoder5.n89 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U149.ZN ) ,
    .I0 ( config1_decoder5.U149.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_79 ) ,
    .IN ( config1_decoder5.U149.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U165.AB ) ,
    .I0 ( config1_decoder5.n100 ) ,
    .I1 ( config1_decoder5.n63 ) ) ;
and ( 
    .Z ( config1_decoder5.U165.ZN ) ,
    .I0 ( config1_decoder5.U165.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_103 ) ,
    .IN ( config1_decoder5.U165.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U95.AB ) ,
    .I0 ( config1_decoder5.n99 ) ,
    .I1 ( config1_decoder5.n101 ) ) ;
and ( 
    .Z ( config1_decoder5.U95.ZN ) ,
    .I0 ( config1_decoder5.U95.AB ) ,
    .I1 ( config1_decoder5.n1 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_102 ) ,
    .IN ( config1_decoder5.U95.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U6.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U6.ZN ) ,
    .I0 ( config1_decoder5.U6.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_47 ) ,
    .IN ( config1_decoder5.U6.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U85.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U85.ZN ) ,
    .I0 ( config1_decoder5.U85.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_2 ) ,
    .IN ( config1_decoder5.U85.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n79 ) ,
    .IN ( config1_decoder5.n99 ) ) ;
nand ( 
    .Z ( config1_decoder5.n83 ) ,
    .I0 ( config1_decoder5.n68 ) ,
    .I1 ( config1_decoder5.n65 ) ) ;
or ( 
    .Z ( config1_decoder5.U71.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U71.ZN ) ,
    .I0 ( config1_decoder5.U71.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_10 ) ,
    .IN ( config1_decoder5.U71.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U61.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U61.ZN ) ,
    .I0 ( config1_decoder5.U61.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_38 ) ,
    .IN ( config1_decoder5.U61.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U16.AB ) ,
    .I0 ( config1_decoder5.n87 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U16.ZN ) ,
    .I0 ( config1_decoder5.U16.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_12 ) ,
    .IN ( config1_decoder5.U16.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n74 ) ,
    .I0 ( config1_decoder5.n70 ) ,
    .I1 ( config1_decoder5.n79 ) ) ;
or ( 
    .Z ( config1_decoder5.U111.AB ) ,
    .I0 ( config1_decoder5.n93 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U111.ZN ) ,
    .I0 ( config1_decoder5.U111.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_82 ) ,
    .IN ( config1_decoder5.U111.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U107.AB ) ,
    .I0 ( config1_decoder5.n91 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U107.ZN ) ,
    .I0 ( config1_decoder5.U107.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_77 ) ,
    .IN ( config1_decoder5.U107.ZN ) ) ;
and ( 
    .Z ( config1_decoder5.n68 ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( masks_hold_reg_8_7 ) ) ;
not ( 
    .O1 ( config1_decoder5.n65 ) ,
    .IN ( masks_hold_reg_8_9 ) ) ;
or ( 
    .Z ( config1_decoder5.U151.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n91 ) ) ;
and ( 
    .Z ( config1_decoder5.U151.ZN ) ,
    .I0 ( config1_decoder5.U151.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_65 ) ,
    .IN ( config1_decoder5.U151.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U96.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n91 ) ) ;
and ( 
    .Z ( config1_decoder5.U96.ZN ) ,
    .I0 ( config1_decoder5.U96.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_73 ) ,
    .IN ( config1_decoder5.U96.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.U1.BN ) ,
    .IN ( config1_decoder5.n95 ) ) ;
nand ( 
    .Z ( config1_decoder5.n98 ) ,
    .I0 ( config1_decoder5.U1.BN ) ,
    .I1 ( config1_decoder5.n94 ) ) ;
or ( 
    .Z ( config1_decoder5.U84.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U84.ZN ) ,
    .I0 ( config1_decoder5.U84.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_3 ) ,
    .IN ( config1_decoder5.U84.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n78 ) ,
    .IN ( config1_decoder5.n97 ) ) ;
not ( 
    .O1 ( config1_decoder5.U44.BN ) ,
    .IN ( config1_decoder5.n82 ) ) ;
nand ( 
    .Z ( config1_decoder5.n101 ) ,
    .I0 ( config1_decoder5.U44.BN ) ,
    .I1 ( config1_decoder5.n94 ) ) ;
or ( 
    .Z ( config1_decoder5.U76.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n81 ) ) ;
and ( 
    .Z ( config1_decoder5.U76.ZN ) ,
    .I0 ( config1_decoder5.U76.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_18 ) ,
    .IN ( config1_decoder5.U76.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U60.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U60.ZN ) ,
    .I0 ( config1_decoder5.U60.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_36 ) ,
    .IN ( config1_decoder5.U60.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U17.AB ) ,
    .I0 ( config1_decoder5.n84 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U17.ZN ) ,
    .I0 ( config1_decoder5.U17.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_11 ) ,
    .IN ( config1_decoder5.U17.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n71 ) ,
    .I0 ( config1_decoder5.n70 ) ,
    .I1 ( config1_decoder5.n76 ) ) ;
or ( 
    .Z ( config1_decoder5.U27.AB ) ,
    .I0 ( config1_decoder5.n90 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U27.ZN ) ,
    .I0 ( config1_decoder5.U27.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_84 ) ,
    .IN ( config1_decoder5.U27.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U110.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n89 ) ) ;
and ( 
    .Z ( config1_decoder5.U110.ZN ) ,
    .I0 ( config1_decoder5.U110.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_91 ) ,
    .IN ( config1_decoder5.U110.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n96 ) ,
    .IN ( config1_decoder5.n77 ) ) ;
not ( 
    .O1 ( config1_decoder5.n75 ) ,
    .IN ( masks_hold_reg_7_9 ) ) ;
nor ( 
    .Z ( config1_decoder5.n80 ) ,
    .I0 ( config1_decoder5.n75 ) ,
    .I1 ( masks_hold_reg_8_10 ) ) ;
nor ( 
    .Z ( config1_decoder5.n76 ) ,
    .I0 ( masks_hold_reg_8_5 ) ,
    .I1 ( masks_hold_reg_8_6 ) ) ;
or ( 
    .Z ( config1_decoder5.U150.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U150.ZN ) ,
    .I0 ( config1_decoder5.U150.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_61 ) ,
    .IN ( config1_decoder5.U150.ZN ) ) ;
not ( 
    .O1 ( config1_decoder5.n69 ) ,
    .IN ( masks_hold_reg_8_10 ) ) ;
or ( 
    .Z ( config1_decoder5.U97.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U97.ZN ) ,
    .I0 ( config1_decoder5.U97.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_23 ) ,
    .IN ( config1_decoder5.U97.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U87.AB ) ,
    .I0 ( config1_decoder5.n92 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U87.ZN ) ,
    .I0 ( config1_decoder5.U87.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_60 ) ,
    .IN ( config1_decoder5.U87.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U57.AB ) ,
    .I0 ( config1_decoder5.n82 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U57.ZN ) ,
    .I0 ( config1_decoder5.U57.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_35 ) ,
    .IN ( config1_decoder5.U57.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U47.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n92 ) ) ;
and ( 
    .Z ( config1_decoder5.U47.ZN ) ,
    .I0 ( config1_decoder5.U47.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_29 ) ,
    .IN ( config1_decoder5.U47.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U77.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n84 ) ) ;
and ( 
    .Z ( config1_decoder5.U77.ZN ) ,
    .I0 ( config1_decoder5.U77.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_19 ) ,
    .IN ( config1_decoder5.U77.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U67.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U67.ZN ) ,
    .I0 ( config1_decoder5.U67.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_52 ) ,
    .IN ( config1_decoder5.U67.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U10.AB ) ,
    .I0 ( config1_decoder5.n83 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U10.ZN ) ,
    .I0 ( config1_decoder5.U10.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_43 ) ,
    .IN ( config1_decoder5.U10.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n87 ) ,
    .I0 ( config1_decoder5.n77 ) ,
    .I1 ( config1_decoder5.n64 ) ) ;
or ( 
    .Z ( config1_decoder5.U26.AB ) ,
    .I0 ( config1_decoder5.n91 ) ,
    .I1 ( config1_decoder5.n85 ) ) ;
and ( 
    .Z ( config1_decoder5.U26.ZN ) ,
    .I0 ( config1_decoder5.U26.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_81 ) ,
    .IN ( config1_decoder5.U26.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U113.AB ) ,
    .I0 ( config1_decoder5.n93 ) ,
    .I1 ( config1_decoder5.n83 ) ) ;
and ( 
    .Z ( config1_decoder5.U113.ZN ) ,
    .I0 ( config1_decoder5.U113.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_78 ) ,
    .IN ( config1_decoder5.U113.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U138.AB ) ,
    .I0 ( config1_decoder5.n99 ) ,
    .I1 ( config1_decoder5.n98 ) ) ;
and ( 
    .Z ( config1_decoder5.U138.ZN ) ,
    .I0 ( config1_decoder5.U138.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_98 ) ,
    .IN ( config1_decoder5.U138.ZN ) ) ;
nor ( 
    .Z ( config1_decoder5.n70 ) ,
    .I0 ( config1_decoder5.n69 ) ,
    .I1 ( masks_hold_reg_7_9 ) ) ;
nor ( 
    .Z ( config1_decoder5.n66 ) ,
    .I0 ( config1_decoder5.n65 ) ,
    .I1 ( masks_hold_reg_8_8 ) ) ;
nand ( 
    .Z ( config1_decoder5.n1 ) ,
    .I0 ( config1_decoder5.n94 ) ,
    .I1 ( config1_decoder5.n60 ) ) ;
or ( 
    .Z ( config1_decoder5.U153.AB ) ,
    .I0 ( config1_decoder5.n100 ) ,
    .I1 ( config1_decoder5.n98 ) ) ;
and ( 
    .Z ( config1_decoder5.U153.ZN ) ,
    .I0 ( config1_decoder5.U153.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_95 ) ,
    .IN ( config1_decoder5.U153.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U141.AB ) ,
    .I0 ( config1_decoder5.n101 ) ,
    .I1 ( config1_decoder5.n100 ) ) ;
and ( 
    .Z ( config1_decoder5.U141.ZN ) ,
    .I0 ( config1_decoder5.U141.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_99 ) ,
    .IN ( config1_decoder5.U141.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U90.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n72 ) ) ;
and ( 
    .Z ( config1_decoder5.U90.ZN ) ,
    .I0 ( config1_decoder5.U90.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_56 ) ,
    .IN ( config1_decoder5.U90.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U3.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U3.ZN ) ,
    .I0 ( config1_decoder5.U3.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_33 ) ,
    .IN ( config1_decoder5.U3.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U86.AB ) ,
    .I0 ( config1_decoder5.n88 ) ,
    .I1 ( config1_decoder5.n73 ) ) ;
and ( 
    .Z ( config1_decoder5.U86.ZN ) ,
    .I0 ( config1_decoder5.U86.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_57 ) ,
    .IN ( config1_decoder5.U86.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U58.AB ) ,
    .I0 ( config1_decoder5.n103 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U58.ZN ) ,
    .I0 ( config1_decoder5.U58.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_39 ) ,
    .IN ( config1_decoder5.U58.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U46.AB ) ,
    .I0 ( config1_decoder5.n104 ) ,
    .I1 ( config1_decoder5.n88 ) ) ;
and ( 
    .Z ( config1_decoder5.U46.ZN ) ,
    .I0 ( config1_decoder5.U46.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_25 ) ,
    .IN ( config1_decoder5.U46.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U74.AB ) ,
    .I0 ( config1_decoder5.n95 ) ,
    .I1 ( config1_decoder5.n71 ) ) ;
and ( 
    .Z ( config1_decoder5.U74.ZN ) ,
    .I0 ( config1_decoder5.U74.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_31 ) ,
    .IN ( config1_decoder5.U74.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U66.AB ) ,
    .I0 ( config1_decoder5.n86 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U66.ZN ) ,
    .I0 ( config1_decoder5.U66.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_54 ) ,
    .IN ( config1_decoder5.U66.ZN ) ) ;
or ( 
    .Z ( config1_decoder5.U11.AB ) ,
    .I0 ( config1_decoder5.n85 ) ,
    .I1 ( config1_decoder5.n74 ) ) ;
and ( 
    .Z ( config1_decoder5.U11.ZN ) ,
    .I0 ( config1_decoder5.U11.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_50 ) ,
    .IN ( config1_decoder5.U11.ZN ) ) ;
nand ( 
    .Z ( config1_decoder5.n72 ) ,
    .I0 ( config1_decoder5.n70 ) ,
    .I1 ( config1_decoder5.n77 ) ) ;
nand ( 
    .Z ( config1_decoder5.n85 ) ,
    .I0 ( config1_decoder5.n66 ) ,
    .I1 ( config1_decoder5.n67 ) ) ;
or ( 
    .Z ( config1_decoder5.U112.AB ) ,
    .I0 ( config1_decoder5.n93 ) ,
    .I1 ( config1_decoder5.n86 ) ) ;
and ( 
    .Z ( config1_decoder5.U112.ZN ) ,
    .I0 ( config1_decoder5.U112.AB ) ,
    .I1 ( config1_decoder5.n2 ) ) ;
not ( 
    .O1 ( config1_onehot_decoded_masks_4_86 ) ,
    .IN ( config1_decoder5.U112.ZN ) ) ;
nor ( 
    .Z ( config1_decoder5.n64 ) ,
    .I0 ( masks_hold_reg_8_10 ) ,
    .I1 ( masks_hold_reg_7_9 ) ) ;
buf ( 
    .O1 ( n36 ) ,
    .IN ( masks_shift_reg_7_5 ) ) ;
buf ( 
    .O1 ( n35 ) ,
    .IN ( masks_shift_reg_4_4 ) ) ;
and ( 
    .Z ( U1022.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_10 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1022.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_10 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1022.EF ) ,
    .I0 ( xor_decoded_masks_11_10 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_10 ) ,
    .I0 ( U1022.AB ) ,
    .I1 ( U1022.CD ) ,
    .I2 ( U1022.EF ) ) ;
and ( 
    .Z ( U1080.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_26 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1080.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_26 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1080.EF ) ,
    .I0 ( xor_decoded_masks_11_26 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_26 ) ,
    .I0 ( U1080.AB ) ,
    .I1 ( U1080.CD ) ,
    .I2 ( U1080.EF ) ) ;
and ( 
    .Z ( U1018.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_24 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1018.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_24 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1018.EF ) ,
    .I0 ( xor_decoded_masks_11_24 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_24 ) ,
    .I0 ( U1018.AB ) ,
    .I1 ( U1018.CD ) ,
    .I2 ( U1018.EF ) ) ;
not ( 
    .O1 ( n39 ) ,
    .IN ( n37 ) ) ;
buf ( 
    .O1 ( n64 ) ,
    .IN ( n57 ) ) ;
buf ( 
    .O1 ( n65 ) ,
    .IN ( n57 ) ) ;
buf ( 
    .O1 ( n63 ) ,
    .IN ( n57 ) ) ;
buf ( 
    .O1 ( n57 ) ,
    .IN ( n1 ) ) ;
and ( 
    .Z ( U370.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_16 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U370.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_16 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U370.EF ) ,
    .I0 ( xor_decoded_masks_11_16 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_16 ) ,
    .I0 ( U370.AB ) ,
    .I1 ( U370.CD ) ,
    .I2 ( U370.EF ) ) ;
and ( 
    .Z ( U1292.AB ) ,
    .I0 ( masks_hold_reg_8_0 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U1292.CD ) ,
    .I0 ( config1_xor_encoded_masks_97 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_97 ) ,
    .I0 ( U1292.AB ) ,
    .I1 ( U1292.CD ) ) ;
and ( 
    .Z ( U399.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_30 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U399.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_30 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U399.EF ) ,
    .I0 ( xor_decoded_masks_11_30 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_30 ) ,
    .I0 ( U399.AB ) ,
    .I1 ( U399.CD ) ,
    .I2 ( U399.EF ) ) ;
and ( 
    .Z ( U398.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_28 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U398.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_28 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U398.EF ) ,
    .I0 ( xor_decoded_masks_11_28 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_28 ) ,
    .I0 ( U398.AB ) ,
    .I1 ( U398.CD ) ,
    .I2 ( U398.EF ) ) ;
and ( 
    .Z ( U884.AB ) ,
    .I0 ( masks_hold_reg_1_10 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U884.CD ) ,
    .I0 ( config1_xor_encoded_masks_10 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_10 ) ,
    .I0 ( U884.AB ) ,
    .I1 ( U884.CD ) ) ;
and ( 
    .Z ( U804.AB ) ,
    .I0 ( masks_hold_reg_12_3 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U804.CD ) ,
    .I0 ( config1_xor_encoded_masks_138 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_138 ) ,
    .I0 ( U804.AB ) ,
    .I1 ( U804.CD ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2801 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I1 ) ) ;
buf ( 
    .O1 ( n78 ) ,
    .IN ( masks_shift_reg_2_3 ) ) ;
buf ( 
    .O1 ( n77 ) ,
    .IN ( masks_shift_reg_9_8 ) ) ;
buf ( 
    .O1 ( n80 ) ,
    .IN ( masks_shift_reg_4_5 ) ) ;
buf ( 
    .O1 ( n81 ) ,
    .IN ( masks_shift_reg_4_1 ) ) ;
buf ( 
    .O1 ( n82 ) ,
    .IN ( masks_shift_reg_4_2 ) ) ;
buf ( 
    .O1 ( n83 ) ,
    .IN ( masks_shift_reg_4_3 ) ) ;
buf ( 
    .O1 ( n84 ) ,
    .IN ( masks_shift_reg_2_6 ) ) ;
buf ( 
    .O1 ( n85 ) ,
    .IN ( masks_shift_reg_2_5 ) ) ;
buf ( 
    .O1 ( n87 ) ,
    .IN ( masks_shift_reg_3_8 ) ) ;
buf ( 
    .O1 ( n88 ) ,
    .IN ( masks_shift_reg_4_6 ) ) ;
buf ( 
    .O1 ( n89 ) ,
    .IN ( masks_shift_reg_4_7 ) ) ;
and ( 
    .Z ( U630.AB ) ,
    .I0 ( masks_hold_reg_13_1 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U630.CD ) ,
    .I0 ( config1_xor_encoded_masks_148 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_148 ) ,
    .I0 ( U630.AB ) ,
    .I1 ( U630.CD ) ) ;
and ( 
    .Z ( U1049.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_26 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1049.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_26 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1049.EF ) ,
    .I0 ( xor_decoded_masks_3_26 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_26 ) ,
    .I0 ( U1049.AB ) ,
    .I1 ( U1049.CD ) ,
    .I2 ( U1049.EF ) ) ;
and ( 
    .Z ( U631.AB ) ,
    .I0 ( masks_hold_reg_13_0 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U631.CD ) ,
    .I0 ( config1_xor_encoded_masks_149 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_149 ) ,
    .I0 ( U631.AB ) ,
    .I1 ( U631.CD ) ) ;
and ( 
    .Z ( U1163.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_17 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1163.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_17 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1163.EF ) ,
    .I0 ( xor_decoded_masks_13_17 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_17 ) ,
    .I0 ( U1163.AB ) ,
    .I1 ( U1163.CD ) ,
    .I2 ( U1163.EF ) ) ;
and ( 
    .Z ( U719.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_86 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U719.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_33 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U719.EF ) ,
    .I0 ( xor_decoded_masks_6_33 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_33 ) ,
    .I0 ( U719.AB ) ,
    .I1 ( U719.CD ) ,
    .I2 ( U719.EF ) ) ;
and ( 
    .Z ( U632.AB ) ,
    .I0 ( masks_hold_reg_1_1 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U632.CD ) ,
    .I0 ( config1_xor_encoded_masks_19 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_19 ) ,
    .I0 ( U632.AB ) ,
    .I1 ( U632.CD ) ) ;
and ( 
    .Z ( U1162.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_37 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1162.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_37 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1162.EF ) ,
    .I0 ( xor_decoded_masks_13_37 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_37 ) ,
    .I0 ( U1162.AB ) ,
    .I1 ( U1162.CD ) ,
    .I2 ( U1162.EF ) ) ;
and ( 
    .Z ( U718.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_82 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U718.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_29 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U718.EF ) ,
    .I0 ( xor_decoded_masks_6_29 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_29 ) ,
    .I0 ( U718.AB ) ,
    .I1 ( U718.CD ) ,
    .I2 ( U718.EF ) ) ;
and ( 
    .Z ( U633.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_112 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U633.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_5 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U633.EF ) ,
    .I0 ( xor_decoded_masks_2_5 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_5 ) ,
    .I0 ( U633.AB ) ,
    .I1 ( U633.CD ) ,
    .I2 ( U633.EF ) ) ;
and ( 
    .Z ( U1161.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_33 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1161.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_33 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1161.EF ) ,
    .I0 ( xor_decoded_masks_13_33 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_33 ) ,
    .I0 ( U1161.AB ) ,
    .I1 ( U1161.CD ) ,
    .I2 ( U1161.EF ) ) ;
and ( 
    .Z ( U634.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_131 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U634.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_24 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U634.EF ) ,
    .I0 ( xor_decoded_masks_2_24 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_24 ) ,
    .I0 ( U634.AB ) ,
    .I1 ( U634.CD ) ,
    .I2 ( U634.EF ) ) ;
and ( 
    .Z ( U1160.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_25 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1160.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_25 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1160.EF ) ,
    .I0 ( xor_decoded_masks_13_25 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_25 ) ,
    .I0 ( U1160.AB ) ,
    .I1 ( U1160.CD ) ,
    .I2 ( U1160.EF ) ) ;
nand ( 
    .Z ( n18 ) ,
    .I0 ( n40 ) ,
    .I1 ( n52 ) ) ;
and ( 
    .Z ( U635.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_139 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U635.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_32 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U635.EF ) ,
    .I0 ( xor_decoded_masks_2_32 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_32 ) ,
    .I0 ( U635.AB ) ,
    .I1 ( U635.CD ) ,
    .I2 ( U635.EF ) ) ;
and ( 
    .Z ( U1167.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_68 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1167.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_15 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1167.EF ) ,
    .I0 ( xor_decoded_masks_14_15 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_15 ) ,
    .I0 ( U1167.AB ) ,
    .I1 ( U1167.CD ) ,
    .I2 ( U1167.EF ) ) ;
nor ( 
    .Z ( n55 ) ,
    .I0 ( n29 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U636.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_143 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U636.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_36 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U636.EF ) ,
    .I0 ( xor_decoded_masks_2_36 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_36 ) ,
    .I0 ( U636.AB ) ,
    .I1 ( U636.CD ) ,
    .I2 ( U636.EF ) ) ;
and ( 
    .Z ( U1166.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_11 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1166.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_11 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1166.EF ) ,
    .I0 ( xor_decoded_masks_13_11 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_11 ) ,
    .I0 ( U1166.AB ) ,
    .I1 ( U1166.CD ) ,
    .I2 ( U1166.EF ) ) ;
and ( 
    .Z ( U637.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_123 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U637.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_16 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U637.EF ) ,
    .I0 ( xor_decoded_masks_2_16 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_16 ) ,
    .I0 ( U637.AB ) ,
    .I1 ( U637.CD ) ,
    .I2 ( U637.EF ) ) ;
and ( 
    .Z ( U1165.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_15 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1165.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_15 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1165.EF ) ,
    .I0 ( xor_decoded_masks_13_15 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_15 ) ,
    .I0 ( U1165.AB ) ,
    .I1 ( U1165.CD ) ,
    .I2 ( U1165.EF ) ) ;
and ( 
    .Z ( U939.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_28 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U939.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_28 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U939.EF ) ,
    .I0 ( xor_decoded_masks_0_28 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_28 ) ,
    .I0 ( U939.AB ) ,
    .I1 ( U939.CD ) ,
    .I2 ( U939.EF ) ) ;
and ( 
    .Z ( U638.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_121 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U638.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_14 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U638.EF ) ,
    .I0 ( xor_decoded_masks_2_14 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_14 ) ,
    .I0 ( U638.AB ) ,
    .I1 ( U638.CD ) ,
    .I2 ( U638.EF ) ) ;
and ( 
    .Z ( U1164.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_21 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1164.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_21 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1164.EF ) ,
    .I0 ( xor_decoded_masks_13_21 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_21 ) ,
    .I0 ( U1164.AB ) ,
    .I1 ( U1164.CD ) ,
    .I2 ( U1164.EF ) ) ;
and ( 
    .Z ( U938.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_20 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U938.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_20 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U938.EF ) ,
    .I0 ( xor_decoded_masks_0_20 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_20 ) ,
    .I0 ( U938.AB ) ,
    .I1 ( U938.CD ) ,
    .I2 ( U938.EF ) ) ;
and ( 
    .Z ( U639.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_85 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U639.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_32 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U639.EF ) ,
    .I0 ( xor_decoded_masks_4_32 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_32 ) ,
    .I0 ( U639.AB ) ,
    .I1 ( U639.CD ) ,
    .I2 ( U639.EF ) ) ;
and ( 
    .Z ( U937.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_97 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U937.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_44 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U937.EF ) ,
    .I0 ( xor_decoded_masks_14_44 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_44 ) ,
    .I0 ( U937.AB ) ,
    .I1 ( U937.CD ) ,
    .I2 ( U937.EF ) ) ;
and ( 
    .Z ( U936.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_44 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U936.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_44 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U936.EF ) ,
    .I0 ( xor_decoded_masks_13_44 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_44 ) ,
    .I0 ( U936.AB ) ,
    .I1 ( U936.CD ) ,
    .I2 ( U936.EF ) ) ;
and ( 
    .Z ( U1169.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_70 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1169.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_17 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1169.EF ) ,
    .I0 ( xor_decoded_masks_14_17 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_17 ) ,
    .I0 ( U1169.AB ) ,
    .I1 ( U1169.CD ) ,
    .I2 ( U1169.EF ) ) ;
and ( 
    .Z ( U858.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_98 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U858.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_44 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U858.EF ) ,
    .I0 ( xor_decoded_masks_1_44 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_44 ) ,
    .I0 ( U858.AB ) ,
    .I1 ( U858.CD ) ,
    .I2 ( U858.EF ) ) ;
and ( 
    .Z ( U935.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_97 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U935.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_44 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U935.EF ) ,
    .I0 ( xor_decoded_masks_10_44 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_44 ) ,
    .I0 ( U935.AB ) ,
    .I1 ( U935.CD ) ,
    .I2 ( U935.EF ) ) ;
and ( 
    .Z ( U1168.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_64 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1168.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_11 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1168.EF ) ,
    .I0 ( xor_decoded_masks_14_11 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_11 ) ,
    .I0 ( U1168.AB ) ,
    .I1 ( U1168.CD ) ,
    .I2 ( U1168.EF ) ) ;
and ( 
    .Z ( U859.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_101 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U859.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_47 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U859.EF ) ,
    .I0 ( xor_decoded_masks_1_47 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_47 ) ,
    .I0 ( U859.AB ) ,
    .I1 ( U859.CD ) ,
    .I2 ( U859.EF ) ) ;
and ( 
    .Z ( U934.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_44 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U934.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_44 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U934.EF ) ,
    .I0 ( xor_decoded_masks_9_44 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_44 ) ,
    .I0 ( U934.AB ) ,
    .I1 ( U934.CD ) ,
    .I2 ( U934.EF ) ) ;
and ( 
    .Z ( U933.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_57 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U933.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_4 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U933.EF ) ,
    .I0 ( xor_decoded_masks_8_4 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_4 ) ,
    .I0 ( U933.AB ) ,
    .I1 ( U933.CD ) ,
    .I2 ( U933.EF ) ) ;
and ( 
    .Z ( U932.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_44 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U932.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_44 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U932.EF ) ,
    .I0 ( xor_decoded_masks_7_44 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_44 ) ,
    .I0 ( U932.AB ) ,
    .I1 ( U932.CD ) ,
    .I2 ( U932.EF ) ) ;
and ( 
    .Z ( U931.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_97 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U931.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_44 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U931.EF ) ,
    .I0 ( xor_decoded_masks_6_44 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_44 ) ,
    .I0 ( U931.AB ) ,
    .I1 ( U931.CD ) ,
    .I2 ( U931.EF ) ) ;
and ( 
    .Z ( U930.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_44 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U930.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_44 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U930.EF ) ,
    .I0 ( xor_decoded_masks_5_44 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_44 ) ,
    .I0 ( U930.AB ) ,
    .I1 ( U930.CD ) ,
    .I2 ( U930.EF ) ) ;
and ( 
    .Z ( U850.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_100 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U850.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_47 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U850.EF ) ,
    .I0 ( xor_decoded_masks_12_47 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_47 ) ,
    .I0 ( U850.AB ) ,
    .I1 ( U850.CD ) ,
    .I2 ( U850.EF ) ) ;
and ( 
    .Z ( U851.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_97 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U851.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_44 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U851.EF ) ,
    .I0 ( xor_decoded_masks_12_44 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_44 ) ,
    .I0 ( U851.AB ) ,
    .I1 ( U851.CD ) ,
    .I2 ( U851.EF ) ) ;
and ( 
    .Z ( U852.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_58 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U852.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_5 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U852.EF ) ,
    .I0 ( xor_decoded_masks_12_5 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_5 ) ,
    .I0 ( U852.AB ) ,
    .I1 ( U852.CD ) ,
    .I2 ( U852.EF ) ) ;
and ( 
    .Z ( U853.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_47 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U853.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_47 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U853.EF ) ,
    .I0 ( xor_decoded_masks_13_47 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_47 ) ,
    .I0 ( U853.AB ) ,
    .I1 ( U853.CD ) ,
    .I2 ( U853.EF ) ) ;
and ( 
    .Z ( U854.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_46 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U854.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_46 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U854.EF ) ,
    .I0 ( xor_decoded_masks_13_46 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_46 ) ,
    .I0 ( U854.AB ) ,
    .I1 ( U854.CD ) ,
    .I2 ( U854.EF ) ) ;
and ( 
    .Z ( U855.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_45 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U855.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_45 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U855.EF ) ,
    .I0 ( xor_decoded_masks_13_45 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_45 ) ,
    .I0 ( U855.AB ) ,
    .I1 ( U855.CD ) ,
    .I2 ( U855.EF ) ) ;
and ( 
    .Z ( U856.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_100 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U856.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_47 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U856.EF ) ,
    .I0 ( xor_decoded_masks_14_47 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_47 ) ,
    .I0 ( U856.AB ) ,
    .I1 ( U856.CD ) ,
    .I2 ( U856.EF ) ) ;
and ( 
    .Z ( U857.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_99 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U857.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_46 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U857.EF ) ,
    .I0 ( xor_decoded_masks_14_46 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_46 ) ,
    .I0 ( U857.AB ) ,
    .I1 ( U857.CD ) ,
    .I2 ( U857.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_10.DI_ ) ,
    .IN ( N135 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_10.CPI_ ) ,
    .IN ( edt_clock ) ) ;
DFF masks_shift_reg_3_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_3_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_3_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_10.DI_ ) ,
    .IN ( N212 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_1_1 ) ) ;
DFF masks_shift_reg_10_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_10_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_10_10 ) ) ;
and ( 
    .Z ( U603.AB ) ,
    .I0 ( masks_hold_reg_9_4 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U603.CD ) ,
    .I0 ( config1_xor_encoded_masks_104 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_104 ) ,
    .I0 ( U603.AB ) ,
    .I1 ( U603.CD ) ) ;
and ( 
    .Z ( U602.AB ) ,
    .I0 ( masks_hold_reg_1_6 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U602.CD ) ,
    .I0 ( config1_xor_encoded_masks_14 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_14 ) ,
    .I0 ( U602.AB ) ,
    .I1 ( U602.CD ) ) ;
and ( 
    .Z ( U1150.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_37 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1150.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_37 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1150.EF ) ,
    .I0 ( xor_decoded_masks_11_37 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_37 ) ,
    .I0 ( U1150.AB ) ,
    .I1 ( U1150.CD ) ,
    .I2 ( U1150.EF ) ) ;
and ( 
    .Z ( U601.AB ) ,
    .I0 ( masks_hold_reg_11_6 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U601.CD ) ,
    .I0 ( config1_xor_encoded_masks_124 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_124 ) ,
    .I0 ( U601.AB ) ,
    .I1 ( U601.CD ) ) ;
and ( 
    .Z ( U1151.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_17 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1151.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_17 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1151.EF ) ,
    .I0 ( xor_decoded_masks_11_17 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_17 ) ,
    .I0 ( U1151.AB ) ,
    .I1 ( U1151.CD ) ,
    .I2 ( U1151.EF ) ) ;
and ( 
    .Z ( U600.AB ) ,
    .I0 ( masks_hold_reg_2_7 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U600.CD ) ,
    .I0 ( config1_xor_encoded_masks_24 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_24 ) ,
    .I0 ( U600.AB ) ,
    .I1 ( U600.CD ) ) ;
and ( 
    .Z ( U1152.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_21 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1152.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_21 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1152.EF ) ,
    .I0 ( xor_decoded_masks_11_21 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_21 ) ,
    .I0 ( U1152.AB ) ,
    .I1 ( U1152.CD ) ,
    .I2 ( U1152.EF ) ) ;
and ( 
    .Z ( U607.AB ) ,
    .I0 ( masks_hold_reg_2_9 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U607.CD ) ,
    .I0 ( config1_xor_encoded_masks_22 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_22 ) ,
    .I0 ( U607.AB ) ,
    .I1 ( U607.CD ) ) ;
and ( 
    .Z ( U1153.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_15 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1153.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_15 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1153.EF ) ,
    .I0 ( xor_decoded_masks_11_15 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_15 ) ,
    .I0 ( U1153.AB ) ,
    .I1 ( U1153.CD ) ,
    .I2 ( U1153.EF ) ) ;
and ( 
    .Z ( U1285.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_50 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1285.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_50 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1285.EF ) ,
    .I0 ( xor_decoded_masks_9_50 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_50 ) ,
    .I0 ( U1285.AB ) ,
    .I1 ( U1285.CD ) ,
    .I2 ( U1285.EF ) ) ;
and ( 
    .Z ( U921.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_99 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U921.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_46 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U921.EF ) ,
    .I0 ( xor_decoded_masks_10_46 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_46 ) ,
    .I0 ( U921.AB ) ,
    .I1 ( U921.CD ) ,
    .I2 ( U921.EF ) ) ;
and ( 
    .Z ( U1282.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_103 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1282.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_50 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1282.EF ) ,
    .I0 ( xor_decoded_masks_6_50 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_50 ) ,
    .I0 ( U1282.AB ) ,
    .I1 ( U1282.CD ) ,
    .I2 ( U1282.EF ) ) ;
and ( 
    .Z ( U1283.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_50 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1283.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_50 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1283.EF ) ,
    .I0 ( xor_decoded_masks_7_50 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_50 ) ,
    .I0 ( U1283.AB ) ,
    .I1 ( U1283.CD ) ,
    .I2 ( U1283.EF ) ) ;
and ( 
    .Z ( U841.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_47 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U841.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_47 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U841.EF ) ,
    .I0 ( xor_decoded_masks_5_47 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_47 ) ,
    .I0 ( U841.AB ) ,
    .I1 ( U841.CD ) ,
    .I2 ( U841.EF ) ) ;
and ( 
    .Z ( U1280.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_103 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1280.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_50 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1280.EF ) ,
    .I0 ( xor_decoded_masks_4_50 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_50 ) ,
    .I0 ( U1280.AB ) ,
    .I1 ( U1280.CD ) ,
    .I2 ( U1280.EF ) ) ;
and ( 
    .Z ( U840.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_57 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U840.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_4 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U840.EF ) ,
    .I0 ( xor_decoded_masks_4_4 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_4 ) ,
    .I0 ( U840.AB ) ,
    .I1 ( U840.CD ) ,
    .I2 ( U840.EF ) ) ;
and ( 
    .Z ( U1281.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_50 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1281.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_50 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1281.EF ) ,
    .I0 ( xor_decoded_masks_5_50 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_50 ) ,
    .I0 ( U1281.AB ) ,
    .I1 ( U1281.CD ) ,
    .I2 ( U1281.EF ) ) ;
and ( 
    .Z ( U843.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_97 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U843.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_44 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U843.EF ) ,
    .I0 ( xor_decoded_masks_8_44 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_44 ) ,
    .I0 ( U843.AB ) ,
    .I1 ( U843.CD ) ,
    .I2 ( U843.EF ) ) ;
and ( 
    .Z ( U842.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_57 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U842.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_4 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U842.EF ) ,
    .I0 ( xor_decoded_masks_6_4 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_4 ) ,
    .I0 ( U842.AB ) ,
    .I1 ( U842.CD ) ,
    .I2 ( U842.EF ) ) ;
and ( 
    .Z ( U845.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_47 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U845.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_47 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U845.EF ) ,
    .I0 ( xor_decoded_masks_9_47 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_47 ) ,
    .I0 ( U845.AB ) ,
    .I1 ( U845.CD ) ,
    .I2 ( U845.EF ) ) ;
and ( 
    .Z ( U713.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_90 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U713.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_37 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U713.EF ) ,
    .I0 ( xor_decoded_masks_4_37 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_37 ) ,
    .I0 ( U713.AB ) ,
    .I1 ( U713.CD ) ,
    .I2 ( U713.EF ) ) ;
and ( 
    .Z ( U1040.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_93 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1040.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_40 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1040.EF ) ,
    .I0 ( xor_decoded_masks_8_40 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_40 ) ,
    .I0 ( U1040.AB ) ,
    .I1 ( U1040.CD ) ,
    .I2 ( U1040.EF ) ) ;
and ( 
    .Z ( U844.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_99 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U844.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_46 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U844.EF ) ,
    .I0 ( xor_decoded_masks_8_46 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_46 ) ,
    .I0 ( U844.AB ) ,
    .I1 ( U844.CD ) ,
    .I2 ( U844.EF ) ) ;
and ( 
    .Z ( U712.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_78 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U712.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_25 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U712.EF ) ,
    .I0 ( xor_decoded_masks_4_25 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_25 ) ,
    .I0 ( U712.AB ) ,
    .I1 ( U712.CD ) ,
    .I2 ( U712.EF ) ) ;
and ( 
    .Z ( U1041.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_40 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1041.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_40 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1041.EF ) ,
    .I0 ( xor_decoded_masks_9_40 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_40 ) ,
    .I0 ( U1041.AB ) ,
    .I1 ( U1041.CD ) ,
    .I2 ( U1041.EF ) ) ;
and ( 
    .Z ( U847.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_98 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U847.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_45 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U847.EF ) ,
    .I0 ( xor_decoded_masks_10_45 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_45 ) ,
    .I0 ( U847.AB ) ,
    .I1 ( U847.CD ) ,
    .I2 ( U847.EF ) ) ;
and ( 
    .Z ( U711.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_86 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U711.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_33 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U711.EF ) ,
    .I0 ( xor_decoded_masks_4_33 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_33 ) ,
    .I0 ( U711.AB ) ,
    .I1 ( U711.CD ) ,
    .I2 ( U711.EF ) ) ;
and ( 
    .Z ( U1042.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_93 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1042.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_40 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1042.EF ) ,
    .I0 ( xor_decoded_masks_10_40 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_40 ) ,
    .I0 ( U1042.AB ) ,
    .I1 ( U1042.CD ) ,
    .I2 ( U1042.EF ) ) ;
and ( 
    .Z ( U846.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_5 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U846.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_5 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U846.EF ) ,
    .I0 ( xor_decoded_masks_9_5 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_5 ) ,
    .I0 ( U846.AB ) ,
    .I1 ( U846.CD ) ,
    .I2 ( U846.EF ) ) ;
and ( 
    .Z ( U710.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_82 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U710.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_29 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U710.EF ) ,
    .I0 ( xor_decoded_masks_4_29 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_29 ) ,
    .I0 ( U710.AB ) ,
    .I1 ( U710.CD ) ,
    .I2 ( U710.EF ) ) ;
and ( 
    .Z ( U818.AB ) ,
    .I0 ( masks_hold_reg_12_5 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U818.CD ) ,
    .I0 ( config1_xor_encoded_masks_136 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_136 ) ,
    .I0 ( U818.AB ) ,
    .I1 ( U818.CD ) ) ;
and ( 
    .Z ( U819.AB ) ,
    .I0 ( masks_hold_reg_3_7 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U819.CD ) ,
    .I0 ( config1_xor_encoded_masks_35 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_35 ) ,
    .I0 ( U819.AB ) ,
    .I1 ( U819.CD ) ) ;
and ( 
    .Z ( U814.AB ) ,
    .I0 ( masks_hold_reg_3_6 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U814.CD ) ,
    .I0 ( config1_xor_encoded_masks_36 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_36 ) ,
    .I0 ( U814.AB ) ,
    .I1 ( U814.CD ) ) ;
and ( 
    .Z ( U815.AB ) ,
    .I0 ( masks_hold_reg_5_8 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U815.CD ) ,
    .I0 ( config1_xor_encoded_masks_56 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_56 ) ,
    .I0 ( U815.AB ) ,
    .I1 ( U815.CD ) ) ;
and ( 
    .Z ( U816.AB ) ,
    .I0 ( masks_hold_reg_7_10 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U816.CD ) ,
    .I0 ( config1_xor_encoded_masks_76 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_76 ) ,
    .I0 ( U816.AB ) ,
    .I1 ( U816.CD ) ) ;
and ( 
    .Z ( U481.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_56 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U481.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_3 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U481.EF ) ,
    .I0 ( xor_decoded_masks_14_3 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_3 ) ,
    .I0 ( U481.AB ) ,
    .I1 ( U481.CD ) ,
    .I2 ( U481.EF ) ) ;
and ( 
    .Z ( U817.AB ) ,
    .I0 ( masks_hold_reg_8_1 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U817.CD ) ,
    .I0 ( config1_xor_encoded_masks_96 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_96 ) ,
    .I0 ( U817.AB ) ,
    .I1 ( U817.CD ) ) ;
and ( 
    .Z ( U480.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_53 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U480.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_0 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U480.EF ) ,
    .I0 ( xor_decoded_masks_14_0 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_0 ) ,
    .I0 ( U480.AB ) ,
    .I1 ( U480.CD ) ,
    .I2 ( U480.EF ) ) ;
and ( 
    .Z ( U810.AB ) ,
    .I0 ( masks_hold_reg_4_0 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U810.CD ) ,
    .I0 ( config1_xor_encoded_masks_53 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_53 ) ,
    .I0 ( U810.AB ) ,
    .I1 ( U810.CD ) ) ;
and ( 
    .Z ( U483.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_58 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U483.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_4 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U483.EF ) ,
    .I0 ( xor_decoded_masks_1_4 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_4 ) ,
    .I0 ( U483.AB ) ,
    .I1 ( U483.CD ) ,
    .I2 ( U483.EF ) ) ;
and ( 
    .Z ( U606.AB ) ,
    .I0 ( masks_hold_reg_2_4 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U606.CD ) ,
    .I0 ( config1_xor_encoded_masks_27 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_27 ) ,
    .I0 ( U606.AB ) ,
    .I1 ( U606.CD ) ) ;
and ( 
    .Z ( U1154.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_11 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1154.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_11 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1154.EF ) ,
    .I0 ( xor_decoded_masks_11_11 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_11 ) ,
    .I0 ( U1154.AB ) ,
    .I1 ( U1154.CD ) ,
    .I2 ( U1154.EF ) ) ;
and ( 
    .Z ( U908.AB ) ,
    .I0 ( masks_hold_reg_7_9 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U908.CD ) ,
    .I0 ( config1_xor_encoded_masks_77 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_77 ) ,
    .I0 ( U908.AB ) ,
    .I1 ( U908.CD ) ) ;
and ( 
    .Z ( U605.AB ) ,
    .I0 ( masks_hold_reg_2_10 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U605.CD ) ,
    .I0 ( config1_xor_encoded_masks_21 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_21 ) ,
    .I0 ( U605.AB ) ,
    .I1 ( U605.CD ) ) ;
and ( 
    .Z ( U1155.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_74 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1155.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_21 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1155.EF ) ,
    .I0 ( xor_decoded_masks_12_21 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_21 ) ,
    .I0 ( U1155.AB ) ,
    .I1 ( U1155.CD ) ,
    .I2 ( U1155.EF ) ) ;
and ( 
    .Z ( U909.AB ) ,
    .I0 ( masks_hold_reg_12_4 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U909.CD ) ,
    .I0 ( config1_xor_encoded_masks_137 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_137 ) ,
    .I0 ( U909.AB ) ,
    .I1 ( U909.CD ) ) ;
and ( 
    .Z ( U604.AB ) ,
    .I0 ( masks_hold_reg_6_8 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U604.CD ) ,
    .I0 ( config1_xor_encoded_masks_67 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_67 ) ,
    .I0 ( U604.AB ) ,
    .I1 ( U604.CD ) ) ;
and ( 
    .Z ( U1156.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_68 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1156.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_15 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1156.EF ) ,
    .I0 ( xor_decoded_masks_12_15 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_15 ) ,
    .I0 ( U1156.AB ) ,
    .I1 ( U1156.CD ) ,
    .I2 ( U1156.EF ) ) ;
and ( 
    .Z ( U1157.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_64 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1157.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_11 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1157.EF ) ,
    .I0 ( xor_decoded_masks_12_11 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_11 ) ,
    .I0 ( U1157.AB ) ,
    .I1 ( U1157.CD ) ,
    .I2 ( U1157.EF ) ) ;
and ( 
    .Z ( U1158.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_70 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1158.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_17 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1158.EF ) ,
    .I0 ( xor_decoded_masks_12_17 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_17 ) ,
    .I0 ( U1158.AB ) ,
    .I1 ( U1158.CD ) ,
    .I2 ( U1158.EF ) ) ;
and ( 
    .Z ( U904.AB ) ,
    .I0 ( masks_hold_reg_9_7 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U904.CD ) ,
    .I0 ( config1_xor_encoded_masks_101 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_101 ) ,
    .I0 ( U904.AB ) ,
    .I1 ( U904.CD ) ) ;
and ( 
    .Z ( U609.AB ) ,
    .I0 ( masks_hold_reg_8_10 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U609.CD ) ,
    .I0 ( config1_xor_encoded_masks_87 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_87 ) ,
    .I0 ( U609.AB ) ,
    .I1 ( U609.CD ) ) ;
and ( 
    .Z ( U1159.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_29 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1159.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_29 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1159.EF ) ,
    .I0 ( xor_decoded_masks_13_29 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_29 ) ,
    .I0 ( U1159.AB ) ,
    .I1 ( U1159.CD ) ,
    .I2 ( U1159.EF ) ) ;
and ( 
    .Z ( U905.AB ) ,
    .I0 ( masks_hold_reg_1_9 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U905.CD ) ,
    .I0 ( config1_xor_encoded_masks_11 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_11 ) ,
    .I0 ( U905.AB ) ,
    .I1 ( U905.CD ) ) ;
and ( 
    .Z ( U608.AB ) ,
    .I0 ( masks_hold_reg_3_0 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U608.CD ) ,
    .I0 ( config1_xor_encoded_masks_42 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_42 ) ,
    .I0 ( U608.AB ) ,
    .I1 ( U608.CD ) ) ;
and ( 
    .Z ( U906.AB ) ,
    .I0 ( n90 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U906.CD ) ,
    .I0 ( config1_xor_encoded_masks_37 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_37 ) ,
    .I0 ( U906.AB ) ,
    .I1 ( U906.CD ) ) ;
and ( 
    .Z ( U907.AB ) ,
    .I0 ( masks_hold_reg_5_7 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U907.CD ) ,
    .I0 ( config1_xor_encoded_masks_57 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_57 ) ,
    .I0 ( U907.AB ) ,
    .I1 ( U907.CD ) ) ;
and ( 
    .Z ( U900.AB ) ,
    .I0 ( masks_hold_reg_12_0 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U900.CD ) ,
    .I0 ( config1_xor_encoded_masks_141 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_141 ) ,
    .I0 ( U900.AB ) ,
    .I1 ( U900.CD ) ) ;
and ( 
    .Z ( U901.AB ) ,
    .I0 ( masks_hold_reg_2_0 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U901.CD ) ,
    .I0 ( config1_xor_encoded_masks_31 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_31 ) ,
    .I0 ( U901.AB ) ,
    .I1 ( U901.CD ) ) ;
and ( 
    .Z ( U902.AB ) ,
    .I0 ( masks_hold_reg_4_2 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U902.CD ) ,
    .I0 ( config1_xor_encoded_masks_51 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_51 ) ,
    .I0 ( U902.AB ) ,
    .I1 ( U902.CD ) ) ;
and ( 
    .Z ( U903.AB ) ,
    .I0 ( masks_hold_reg_6_4 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U903.CD ) ,
    .I0 ( config1_xor_encoded_masks_71 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_71 ) ,
    .I0 ( U903.AB ) ,
    .I1 ( U903.CD ) ) ;
and ( 
    .Z ( U829.AB ) ,
    .I0 ( masks_hold_reg_11_9 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U829.CD ) ,
    .I0 ( config1_xor_encoded_masks_121 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_121 ) ,
    .I0 ( U829.AB ) ,
    .I1 ( U829.CD ) ) ;
and ( 
    .Z ( U828.AB ) ,
    .I0 ( masks_hold_reg_12_10 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U828.CD ) ,
    .I0 ( config1_xor_encoded_masks_131 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_131 ) ,
    .I0 ( U828.AB ) ,
    .I1 ( U828.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_7_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_0.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_0 ) ,
    .IN ( masks_hold_reg_7_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_0.QT ) ,
    .I1 ( masks_hold_reg_7_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_0.ED ) ,
    .S ( masks_hold_reg_7_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_0.ED ) ,
    .I1 ( masks_hold_reg_7_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_0.QT ) ) ;
and ( 
    .Z ( U827.AB ) ,
    .I0 ( masks_hold_reg_0_6 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U827.CD ) ,
    .I0 ( config1_xor_encoded_masks_3 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_3 ) ,
    .I0 ( U827.AB ) ,
    .I1 ( U827.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_7_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_1.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_1 ) ,
    .IN ( masks_hold_reg_7_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_1.QT ) ,
    .I1 ( masks_hold_reg_7_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_1.ED ) ,
    .S ( masks_hold_reg_7_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_1.ED ) ,
    .I1 ( masks_hold_reg_7_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_1.QT ) ) ;
and ( 
    .Z ( U826.AB ) ,
    .I0 ( masks_hold_reg_6_5 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U826.CD ) ,
    .I0 ( config1_xor_encoded_masks_70 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_70 ) ,
    .I0 ( U826.AB ) ,
    .I1 ( U826.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_7_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_2.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_2 ) ,
    .IN ( masks_hold_reg_7_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_2.QT ) ,
    .I1 ( masks_hold_reg_7_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_2.ED ) ,
    .S ( masks_hold_reg_7_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_2.ED ) ,
    .I1 ( masks_hold_reg_7_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_2.QT ) ) ;
and ( 
    .Z ( U825.AB ) ,
    .I0 ( masks_hold_reg_10_4 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U825.CD ) ,
    .I0 ( config1_xor_encoded_masks_115 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_115 ) ,
    .I0 ( U825.AB ) ,
    .I1 ( U825.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_7_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_3.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_3 ) ,
    .IN ( masks_hold_reg_7_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_3.QT ) ,
    .I1 ( masks_hold_reg_7_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_3.ED ) ,
    .S ( masks_hold_reg_7_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_3.ED ) ,
    .I1 ( masks_hold_reg_7_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_3.QT ) ) ;
and ( 
    .Z ( U824.AB ) ,
    .I0 ( masks_hold_reg_10_3 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U824.CD ) ,
    .I0 ( config1_xor_encoded_masks_116 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_116 ) ,
    .I0 ( U824.AB ) ,
    .I1 ( U824.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_7_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_4.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_4 ) ,
    .IN ( masks_hold_reg_7_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_4.QT ) ,
    .I1 ( masks_hold_reg_7_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_4.ED ) ,
    .S ( masks_hold_reg_7_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_4.ED ) ,
    .I1 ( masks_hold_reg_7_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_4.QT ) ) ;
and ( 
    .Z ( U823.AB ) ,
    .I0 ( masks_hold_reg_11_7 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U823.CD ) ,
    .I0 ( config1_xor_encoded_masks_123 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_123 ) ,
    .I0 ( U823.AB ) ,
    .I1 ( U823.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_7_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_5.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_5 ) ,
    .IN ( masks_hold_reg_7_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_5.QT ) ,
    .I1 ( masks_hold_reg_7_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_5.ED ) ,
    .S ( masks_hold_reg_7_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_5.ED ) ,
    .I1 ( masks_hold_reg_7_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_5.QT ) ) ;
and ( 
    .Z ( U822.AB ) ,
    .I0 ( masks_hold_reg_8_2 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U822.CD ) ,
    .I0 ( config1_xor_encoded_masks_95 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_95 ) ,
    .I0 ( U822.AB ) ,
    .I1 ( U822.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_7_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_6.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_6 ) ,
    .IN ( masks_hold_reg_7_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_6.QT ) ,
    .I1 ( masks_hold_reg_7_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_6.ED ) ,
    .S ( masks_hold_reg_7_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_6.ED ) ,
    .I1 ( masks_hold_reg_7_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_6.QT ) ) ;
and ( 
    .Z ( U821.AB ) ,
    .I0 ( masks_hold_reg_6_0 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U821.CD ) ,
    .I0 ( config1_xor_encoded_masks_75 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_75 ) ,
    .I0 ( U821.AB ) ,
    .I1 ( U821.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_7_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_7.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_7 ) ,
    .IN ( masks_hold_reg_7_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_7.QT ) ,
    .I1 ( masks_hold_reg_7_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_7.ED ) ,
    .S ( masks_hold_reg_7_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_7.ED ) ,
    .I1 ( masks_hold_reg_7_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_7.QT ) ) ;
and ( 
    .Z ( U820.AB ) ,
    .I0 ( masks_hold_reg_5_9 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U820.CD ) ,
    .I0 ( config1_xor_encoded_masks_55 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_55 ) ,
    .I0 ( U820.AB ) ,
    .I1 ( U820.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_7_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_8.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_8 ) ,
    .IN ( masks_hold_reg_7_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_8.QT ) ,
    .I1 ( masks_hold_reg_7_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_8.ED ) ,
    .S ( masks_hold_reg_7_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_8.ED ) ,
    .I1 ( masks_hold_reg_7_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_7_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_0_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_9.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_9 ) ,
    .IN ( masks_hold_reg_7_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_9.QT ) ,
    .I1 ( masks_hold_reg_7_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_9.ED ) ,
    .S ( masks_hold_reg_7_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_9.ED ) ,
    .I1 ( masks_hold_reg_7_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_9.QT ) ) ;
and ( 
    .Z ( U612.AB ) ,
    .I0 ( masks_hold_reg_1_3 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U612.CD ) ,
    .I0 ( config1_xor_encoded_masks_17 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_17 ) ,
    .I0 ( U612.AB ) ,
    .I1 ( U612.CD ) ) ;
and ( 
    .Z ( U613.AB ) ,
    .I0 ( masks_hold_reg_13_5 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U613.CD ) ,
    .I0 ( config1_xor_encoded_masks_144 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_144 ) ,
    .I0 ( U613.AB ) ,
    .I1 ( U613.CD ) ) ;
and ( 
    .Z ( U1141.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_17 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1141.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_17 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1141.EF ) ,
    .I0 ( xor_decoded_masks_9_17 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_17 ) ,
    .I0 ( U1141.AB ) ,
    .I1 ( U1141.CD ) ,
    .I2 ( U1141.EF ) ) ;
and ( 
    .Z ( U610.AB ) ,
    .I0 ( masks_hold_reg_13_2 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U610.CD ) ,
    .I0 ( config1_xor_encoded_masks_147 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_147 ) ,
    .I0 ( U610.AB ) ,
    .I1 ( U610.CD ) ) ;
and ( 
    .Z ( U1140.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_37 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1140.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_37 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1140.EF ) ,
    .I0 ( xor_decoded_masks_9_37 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_37 ) ,
    .I0 ( U1140.AB ) ,
    .I1 ( U1140.CD ) ,
    .I2 ( U1140.EF ) ) ;
and ( 
    .Z ( U611.AB ) ,
    .I0 ( masks_hold_reg_13_7 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U611.CD ) ,
    .I0 ( config1_xor_encoded_masks_142 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_142 ) ,
    .I0 ( U611.AB ) ,
    .I1 ( U611.CD ) ) ;
and ( 
    .Z ( U1143.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_15 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1143.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_15 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1143.EF ) ,
    .I0 ( xor_decoded_masks_9_15 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_15 ) ,
    .I0 ( U1143.AB ) ,
    .I1 ( U1143.CD ) ,
    .I2 ( U1143.EF ) ) ;
and ( 
    .Z ( U616.AB ) ,
    .I0 ( masks_hold_reg_9_6 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U616.CD ) ,
    .I0 ( config1_xor_encoded_masks_102 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_102 ) ,
    .I0 ( U616.AB ) ,
    .I1 ( U616.CD ) ) ;
and ( 
    .Z ( U1142.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_21 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1142.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_21 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1142.EF ) ,
    .I0 ( xor_decoded_masks_9_21 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_21 ) ,
    .I0 ( U1142.AB ) ,
    .I1 ( U1142.CD ) ,
    .I2 ( U1142.EF ) ) ;
and ( 
    .Z ( U588.AB ) ,
    .I0 ( masks_hold_reg_1_4 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U588.CD ) ,
    .I0 ( config1_xor_encoded_masks_16 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_16 ) ,
    .I0 ( U588.AB ) ,
    .I1 ( U588.CD ) ) ;
and ( 
    .Z ( U617.AB ) ,
    .I0 ( masks_hold_reg_9_2 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U617.CD ) ,
    .I0 ( config1_xor_encoded_masks_106 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_106 ) ,
    .I0 ( U617.AB ) ,
    .I1 ( U617.CD ) ) ;
and ( 
    .Z ( U1145.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_64 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1145.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_11 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1145.EF ) ,
    .I0 ( xor_decoded_masks_10_11 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_11 ) ,
    .I0 ( U1145.AB ) ,
    .I1 ( U1145.CD ) ,
    .I2 ( U1145.EF ) ) ;
and ( 
    .Z ( U589.AB ) ,
    .I0 ( masks_hold_reg_11_5 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U589.CD ) ,
    .I0 ( config1_xor_encoded_masks_125 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_125 ) ,
    .I0 ( U589.AB ) ,
    .I1 ( U589.CD ) ) ;
and ( 
    .Z ( U919.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_46 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U919.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_46 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U919.EF ) ,
    .I0 ( xor_decoded_masks_7_46 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_46 ) ,
    .I0 ( U919.AB ) ,
    .I1 ( U919.CD ) ,
    .I2 ( U919.EF ) ) ;
and ( 
    .Z ( U614.AB ) ,
    .I0 ( masks_hold_reg_5_2 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U614.CD ) ,
    .I0 ( config1_xor_encoded_masks_62 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_62 ) ,
    .I0 ( U614.AB ) ,
    .I1 ( U614.CD ) ) ;
and ( 
    .Z ( U1144.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_68 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1144.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_15 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1144.EF ) ,
    .I0 ( xor_decoded_masks_10_15 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_15 ) ,
    .I0 ( U1144.AB ) ,
    .I1 ( U1144.CD ) ,
    .I2 ( U1144.EF ) ) ;
and ( 
    .Z ( U918.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_99 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U918.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_46 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U918.EF ) ,
    .I0 ( xor_decoded_masks_6_46 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_46 ) ,
    .I0 ( U918.AB ) ,
    .I1 ( U918.CD ) ,
    .I2 ( U918.EF ) ) ;
and ( 
    .Z ( U615.AB ) ,
    .I0 ( masks_hold_reg_7_4 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U615.CD ) ,
    .I0 ( config1_xor_encoded_masks_82 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_82 ) ,
    .I0 ( U615.AB ) ,
    .I1 ( U615.CD ) ) ;
and ( 
    .Z ( U1147.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_29 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1147.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_29 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1147.EF ) ,
    .I0 ( xor_decoded_masks_11_29 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_29 ) ,
    .I0 ( U1147.AB ) ,
    .I1 ( U1147.CD ) ,
    .I2 ( U1147.EF ) ) ;
and ( 
    .Z ( U1146.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_70 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1146.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_17 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1146.EF ) ,
    .I0 ( xor_decoded_masks_10_17 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_17 ) ,
    .I0 ( U1146.AB ) ,
    .I1 ( U1146.CD ) ,
    .I2 ( U1146.EF ) ) ;
and ( 
    .Z ( U1149.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_33 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1149.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_33 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1149.EF ) ,
    .I0 ( xor_decoded_masks_11_33 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_33 ) ,
    .I0 ( U1149.AB ) ,
    .I1 ( U1149.CD ) ,
    .I2 ( U1149.EF ) ) ;
and ( 
    .Z ( U915.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_46 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U915.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_46 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U915.EF ) ,
    .I0 ( xor_decoded_masks_3_46 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_46 ) ,
    .I0 ( U915.AB ) ,
    .I1 ( U915.CD ) ,
    .I2 ( U915.EF ) ) ;
and ( 
    .Z ( U618.AB ) ,
    .I0 ( masks_hold_reg_7_0 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U618.CD ) ,
    .I0 ( config1_xor_encoded_masks_86 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_86 ) ,
    .I0 ( U618.AB ) ,
    .I1 ( U618.CD ) ) ;
and ( 
    .Z ( U1148.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_25 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1148.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_25 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1148.EF ) ,
    .I0 ( xor_decoded_masks_11_25 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_25 ) ,
    .I0 ( U1148.AB ) ,
    .I1 ( U1148.CD ) ,
    .I2 ( U1148.EF ) ) ;
and ( 
    .Z ( U914.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_153 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U914.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_46 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U914.EF ) ,
    .I0 ( xor_decoded_masks_2_46 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_46 ) ,
    .I0 ( U914.AB ) ,
    .I1 ( U914.CD ) ,
    .I2 ( U914.EF ) ) ;
and ( 
    .Z ( U619.AB ) ,
    .I0 ( masks_hold_reg_7_1 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U619.CD ) ,
    .I0 ( config1_xor_encoded_masks_85 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_85 ) ,
    .I0 ( U619.AB ) ,
    .I1 ( U619.CD ) ) ;
and ( 
    .Z ( U917.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_46 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U917.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_46 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U917.EF ) ,
    .I0 ( xor_decoded_masks_5_46 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_46 ) ,
    .I0 ( U917.AB ) ,
    .I1 ( U917.CD ) ,
    .I2 ( U917.EF ) ) ;
and ( 
    .Z ( U580.AB ) ,
    .I0 ( masks_hold_reg_11_2 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U580.CD ) ,
    .I0 ( config1_xor_encoded_masks_128 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_128 ) ,
    .I0 ( U580.AB ) ,
    .I1 ( U580.CD ) ) ;
and ( 
    .Z ( U916.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_99 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U916.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_46 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U916.EF ) ,
    .I0 ( xor_decoded_masks_4_46 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_46 ) ,
    .I0 ( U916.AB ) ,
    .I1 ( U916.CD ) ,
    .I2 ( U916.EF ) ) ;
and ( 
    .Z ( U581.AB ) ,
    .I0 ( masks_hold_reg_1_2 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U581.CD ) ,
    .I0 ( config1_xor_encoded_masks_18 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_18 ) ,
    .I0 ( U581.AB ) ,
    .I1 ( U581.CD ) ) ;
and ( 
    .Z ( U911.AB ) ,
    .I0 ( masks_hold_reg_0_2 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U911.CD ) ,
    .I0 ( config1_xor_encoded_masks_7 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_7 ) ,
    .I0 ( U911.AB ) ,
    .I1 ( U911.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_10.DI_ ) ,
    .IN ( N124 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_10.CPI_ ) ,
    .IN ( edt_clock ) ) ;
DFF masks_shift_reg_2_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_2_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_2_10 ) ) ;
and ( 
    .Z ( U1043.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_40 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1043.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_40 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1043.EF ) ,
    .I0 ( xor_decoded_masks_11_40 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_40 ) ,
    .I0 ( U1043.AB ) ,
    .I1 ( U1043.CD ) ,
    .I2 ( U1043.EF ) ) ;
and ( 
    .Z ( U717.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_70 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U717.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_17 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U717.EF ) ,
    .I0 ( xor_decoded_masks_4_17 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_17 ) ,
    .I0 ( U717.AB ) ,
    .I1 ( U717.CD ) ,
    .I2 ( U717.EF ) ) ;
and ( 
    .Z ( U1044.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_93 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1044.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_40 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1044.EF ) ,
    .I0 ( xor_decoded_masks_12_40 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_40 ) ,
    .I0 ( U1044.AB ) ,
    .I1 ( U1044.CD ) ,
    .I2 ( U1044.EF ) ) ;
and ( 
    .Z ( U716.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_64 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U716.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_11 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U716.EF ) ,
    .I0 ( xor_decoded_masks_4_11 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_11 ) ,
    .I0 ( U716.AB ) ,
    .I1 ( U716.CD ) ,
    .I2 ( U716.EF ) ) ;
and ( 
    .Z ( U1045.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_40 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1045.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_40 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1045.EF ) ,
    .I0 ( xor_decoded_masks_13_40 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_40 ) ,
    .I0 ( U1045.AB ) ,
    .I1 ( U1045.CD ) ,
    .I2 ( U1045.EF ) ) ;
and ( 
    .Z ( U715.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_68 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U715.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_15 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U715.EF ) ,
    .I0 ( xor_decoded_masks_4_15 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_15 ) ,
    .I0 ( U715.AB ) ,
    .I1 ( U715.CD ) ,
    .I2 ( U715.EF ) ) ;
and ( 
    .Z ( U1046.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_93 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1046.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_40 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1046.EF ) ,
    .I0 ( xor_decoded_masks_14_40 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_40 ) ,
    .I0 ( U1046.AB ) ,
    .I1 ( U1046.CD ) ,
    .I2 ( U1046.EF ) ) ;
and ( 
    .Z ( U714.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_74 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U714.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_21 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U714.EF ) ,
    .I0 ( xor_decoded_masks_4_21 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_21 ) ,
    .I0 ( U714.AB ) ,
    .I1 ( U714.CD ) ,
    .I2 ( U714.EF ) ) ;
and ( 
    .Z ( U1047.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_94 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1047.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_40 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1047.EF ) ,
    .I0 ( xor_decoded_masks_1_40 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_40 ) ,
    .I0 ( U1047.AB ) ,
    .I1 ( U1047.CD ) ,
    .I2 ( U1047.EF ) ) ;
and ( 
    .Z ( U1048.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_50 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1048.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_50 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1048.EF ) ,
    .I0 ( xor_decoded_masks_0_50 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_50 ) ,
    .I0 ( U1048.AB ) ,
    .I1 ( U1048.CD ) ,
    .I2 ( U1048.EF ) ) ;
and ( 
    .Z ( U1187.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_27 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1187.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_27 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1187.EF ) ,
    .I0 ( xor_decoded_masks_3_27 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_27 ) ,
    .I0 ( U1187.AB ) ,
    .I1 ( U1187.CD ) ,
    .I2 ( U1187.EF ) ) ;
and ( 
    .Z ( U1186.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_1 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1186.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_1 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1186.EF ) ,
    .I0 ( xor_decoded_masks_0_1 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_1 ) ,
    .I0 ( U1186.AB ) ,
    .I1 ( U1186.CD ) ,
    .I2 ( U1186.EF ) ) ;
and ( 
    .Z ( U1181.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_41 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1181.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_41 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1181.EF ) ,
    .I0 ( xor_decoded_masks_13_41 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_41 ) ,
    .I0 ( U1181.AB ) ,
    .I1 ( U1181.CD ) ,
    .I2 ( U1181.EF ) ) ;
and ( 
    .Z ( U1180.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_94 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1180.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_41 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1180.EF ) ,
    .I0 ( xor_decoded_masks_12_41 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_41 ) ,
    .I0 ( U1180.AB ) ,
    .I1 ( U1180.CD ) ,
    .I2 ( U1180.EF ) ) ;
and ( 
    .Z ( U1183.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_95 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1183.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_41 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1183.EF ) ,
    .I0 ( xor_decoded_masks_1_41 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_41 ) ,
    .I0 ( U1183.AB ) ,
    .I1 ( U1183.CD ) ,
    .I2 ( U1183.EF ) ) ;
and ( 
    .Z ( U1182.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_94 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1182.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_41 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1182.EF ) ,
    .I0 ( xor_decoded_masks_14_41 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_41 ) ,
    .I0 ( U1182.AB ) ,
    .I1 ( U1182.CD ) ,
    .I2 ( U1182.EF ) ) ;
and ( 
    .Z ( U788.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_77 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U788.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_23 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U788.EF ) ,
    .I0 ( xor_decoded_masks_1_23 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_23 ) ,
    .I0 ( U788.AB ) ,
    .I1 ( U788.CD ) ,
    .I2 ( U788.EF ) ) ;
and ( 
    .Z ( U789.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_67 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U789.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_13 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U789.EF ) ,
    .I0 ( xor_decoded_masks_1_13 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_13 ) ,
    .I0 ( U789.AB ) ,
    .I1 ( U789.CD ) ,
    .I2 ( U789.EF ) ) ;
and ( 
    .Z ( U782.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_80 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U782.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_27 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U782.EF ) ,
    .I0 ( xor_decoded_masks_14_27 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_27 ) ,
    .I0 ( U782.AB ) ,
    .I1 ( U782.CD ) ,
    .I2 ( U782.EF ) ) ;
and ( 
    .Z ( U783.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_92 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U783.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_39 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U783.EF ) ,
    .I0 ( xor_decoded_masks_14_39 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_39 ) ,
    .I0 ( U783.AB ) ,
    .I1 ( U783.CD ) ,
    .I2 ( U783.EF ) ) ;
and ( 
    .Z ( U780.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_88 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U780.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_35 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U780.EF ) ,
    .I0 ( xor_decoded_masks_12_35 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_35 ) ,
    .I0 ( U780.AB ) ,
    .I1 ( U780.CD ) ,
    .I2 ( U780.EF ) ) ;
and ( 
    .Z ( U781.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_88 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U781.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_35 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U781.EF ) ,
    .I0 ( xor_decoded_masks_14_35 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_35 ) ,
    .I0 ( U781.AB ) ,
    .I1 ( U781.CD ) ,
    .I2 ( U781.EF ) ) ;
and ( 
    .Z ( U786.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_93 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U786.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_39 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U786.EF ) ,
    .I0 ( xor_decoded_masks_1_39 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_39 ) ,
    .I0 ( U786.AB ) ,
    .I1 ( U786.CD ) ,
    .I2 ( U786.EF ) ) ;
and ( 
    .Z ( U787.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_63 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U787.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_9 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U787.EF ) ,
    .I0 ( xor_decoded_masks_1_9 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_9 ) ,
    .I0 ( U787.AB ) ,
    .I1 ( U787.CD ) ,
    .I2 ( U787.EF ) ) ;
and ( 
    .Z ( U784.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_81 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U784.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_27 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U784.EF ) ,
    .I0 ( xor_decoded_masks_1_27 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_27 ) ,
    .I0 ( U784.AB ) ,
    .I1 ( U784.CD ) ,
    .I2 ( U784.EF ) ) ;
and ( 
    .Z ( U785.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_89 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U785.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_35 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U785.EF ) ,
    .I0 ( xor_decoded_masks_1_35 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_35 ) ,
    .I0 ( U785.AB ) ,
    .I1 ( U785.CD ) ,
    .I2 ( U785.EF ) ) ;
and ( 
    .Z ( U799.AB ) ,
    .I0 ( masks_hold_reg_0_3 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U799.CD ) ,
    .I0 ( config1_xor_encoded_masks_6 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_6 ) ,
    .I0 ( U799.AB ) ,
    .I1 ( U799.CD ) ) ;
and ( 
    .Z ( U798.AB ) ,
    .I0 ( masks_hold_reg_10_0 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U798.CD ) ,
    .I0 ( config1_xor_encoded_masks_119 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_119 ) ,
    .I0 ( U798.AB ) ,
    .I1 ( U798.CD ) ) ;
and ( 
    .Z ( U793.AB ) ,
    .I0 ( masks_hold_reg_3_3 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U793.CD ) ,
    .I0 ( config1_xor_encoded_masks_39 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_39 ) ,
    .I0 ( U793.AB ) ,
    .I1 ( U793.CD ) ) ;
and ( 
    .Z ( U792.AB ) ,
    .I0 ( masks_hold_reg_0_1 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U792.CD ) ,
    .I0 ( config1_xor_encoded_masks_8 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_8 ) ,
    .I0 ( U792.AB ) ,
    .I1 ( U792.CD ) ) ;
and ( 
    .Z ( U582.AB ) ,
    .I0 ( masks_hold_reg_4_10 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U582.CD ) ,
    .I0 ( config1_xor_encoded_masks_43 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_43 ) ,
    .I0 ( U582.AB ) ,
    .I1 ( U582.CD ) ) ;
and ( 
    .Z ( U910.AB ) ,
    .I0 ( masks_hold_reg_1_8 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U910.CD ) ,
    .I0 ( config1_xor_encoded_masks_12 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_12 ) ,
    .I0 ( U910.AB ) ,
    .I1 ( U910.CD ) ) ;
and ( 
    .Z ( U583.AB ) ,
    .I0 ( masks_hold_reg_5_1 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U583.CD ) ,
    .I0 ( config1_xor_encoded_masks_63 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_63 ) ,
    .I0 ( U583.AB ) ,
    .I1 ( U583.CD ) ) ;
and ( 
    .Z ( U913.AB ) ,
    .I0 ( masks_hold_reg_3_10 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U913.CD ) ,
    .I0 ( config1_xor_encoded_masks_32 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_32 ) ,
    .I0 ( U913.AB ) ,
    .I1 ( U913.CD ) ) ;
and ( 
    .Z ( U584.AB ) ,
    .I0 ( masks_hold_reg_7_3 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U584.CD ) ,
    .I0 ( config1_xor_encoded_masks_83 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_83 ) ,
    .I0 ( U584.AB ) ,
    .I1 ( U584.CD ) ) ;
and ( 
    .Z ( U912.AB ) ,
    .I0 ( masks_hold_reg_10_2 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U912.CD ) ,
    .I0 ( config1_xor_encoded_masks_117 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_117 ) ,
    .I0 ( U912.AB ) ,
    .I1 ( U912.CD ) ) ;
and ( 
    .Z ( U838.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_100 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U838.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_47 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U838.EF ) ,
    .I0 ( xor_decoded_masks_4_47 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_47 ) ,
    .I0 ( U838.AB ) ,
    .I1 ( U838.CD ) ,
    .I2 ( U838.EF ) ) ;
and ( 
    .Z ( U585.AB ) ,
    .I0 ( masks_hold_reg_13_6 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U585.CD ) ,
    .I0 ( config1_xor_encoded_masks_143 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_143 ) ,
    .I0 ( U585.AB ) ,
    .I1 ( U585.CD ) ) ;
and ( 
    .Z ( U839.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_97 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U839.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_44 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U839.EF ) ,
    .I0 ( xor_decoded_masks_4_44 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_44 ) ,
    .I0 ( U839.AB ) ,
    .I1 ( U839.CD ) ,
    .I2 ( U839.EF ) ) ;
and ( 
    .Z ( U586.AB ) ,
    .I0 ( masks_hold_reg_11_4 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U586.CD ) ,
    .I0 ( config1_xor_encoded_masks_126 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_126 ) ,
    .I0 ( U586.AB ) ,
    .I1 ( U586.CD ) ) ;
and ( 
    .Z ( U836.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_10 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U836.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_10 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U836.EF ) ,
    .I0 ( xor_decoded_masks_13_10 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_10 ) ,
    .I0 ( U836.AB ) ,
    .I1 ( U836.CD ) ,
    .I2 ( U836.EF ) ) ;
and ( 
    .Z ( U587.AB ) ,
    .I0 ( masks_hold_reg_13_3 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U587.CD ) ,
    .I0 ( config1_xor_encoded_masks_146 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_146 ) ,
    .I0 ( U587.AB ) ,
    .I1 ( U587.CD ) ) ;
and ( 
    .Z ( U837.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_1 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U837.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_1 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U837.EF ) ,
    .I0 ( xor_decoded_masks_3_1 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_1 ) ,
    .I0 ( U837.AB ) ,
    .I1 ( U837.CD ) ,
    .I2 ( U837.EF ) ) ;
and ( 
    .Z ( U834.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_32 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U834.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_32 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U834.EF ) ,
    .I0 ( xor_decoded_masks_11_32 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_32 ) ,
    .I0 ( U834.AB ) ,
    .I1 ( U834.CD ) ,
    .I2 ( U834.EF ) ) ;
and ( 
    .Z ( U835.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_32 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U835.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_32 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U835.EF ) ,
    .I0 ( xor_decoded_masks_13_32 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_32 ) ,
    .I0 ( U835.AB ) ,
    .I1 ( U835.CD ) ,
    .I2 ( U835.EF ) ) ;
and ( 
    .Z ( U832.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_11 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U832.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_11 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U832.EF ) ,
    .I0 ( xor_decoded_masks_9_11 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_11 ) ,
    .I0 ( U832.AB ) ,
    .I1 ( U832.CD ) ,
    .I2 ( U832.EF ) ) ;
and ( 
    .Z ( U833.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_74 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U833.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_21 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U833.EF ) ,
    .I0 ( xor_decoded_masks_10_21 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_21 ) ,
    .I0 ( U833.AB ) ,
    .I1 ( U833.CD ) ,
    .I2 ( U833.EF ) ) ;
and ( 
    .Z ( U830.AB ) ,
    .I0 ( masks_hold_reg_4_3 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U830.CD ) ,
    .I0 ( config1_xor_encoded_masks_50 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_50 ) ,
    .I0 ( U830.AB ) ,
    .I1 ( U830.CD ) ) ;
and ( 
    .Z ( U831.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_14 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U831.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_14 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U831.EF ) ,
    .I0 ( xor_decoded_masks_9_14 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_14 ) ,
    .I0 ( U831.AB ) ,
    .I1 ( U831.CD ) ,
    .I2 ( U831.EF ) ) ;
and ( 
    .Z ( U1099.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_149 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1099.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_42 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1099.EF ) ,
    .I0 ( xor_decoded_masks_2_42 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_42 ) ,
    .I0 ( U1099.AB ) ,
    .I1 ( U1099.CD ) ,
    .I2 ( U1099.EF ) ) ;
and ( 
    .Z ( U1098.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_71 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1098.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_18 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1098.EF ) ,
    .I0 ( xor_decoded_masks_14_18 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_18 ) ,
    .I0 ( U1098.AB ) ,
    .I1 ( U1098.CD ) ,
    .I2 ( U1098.EF ) ) ;
and ( 
    .Z ( U1095.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_12 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1095.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_12 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1095.EF ) ,
    .I0 ( xor_decoded_masks_13_12 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_12 ) ,
    .I0 ( U1095.AB ) ,
    .I1 ( U1095.CD ) ,
    .I2 ( U1095.EF ) ) ;
and ( 
    .Z ( U1094.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_8 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1094.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_8 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1094.EF ) ,
    .I0 ( xor_decoded_masks_13_8 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_8 ) ,
    .I0 ( U1094.AB ) ,
    .I1 ( U1094.CD ) ,
    .I2 ( U1094.EF ) ) ;
and ( 
    .Z ( U1097.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_65 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1097.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_12 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1097.EF ) ,
    .I0 ( xor_decoded_masks_14_12 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_12 ) ,
    .I0 ( U1097.AB ) ,
    .I1 ( U1097.CD ) ,
    .I2 ( U1097.EF ) ) ;
and ( 
    .Z ( U1096.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_61 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1096.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_8 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1096.EF ) ,
    .I0 ( xor_decoded_masks_14_8 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_8 ) ,
    .I0 ( U1096.AB ) ,
    .I1 ( U1096.CD ) ,
    .I2 ( U1096.EF ) ) ;
and ( 
    .Z ( U1091.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_34 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1091.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_34 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1091.EF ) ,
    .I0 ( xor_decoded_masks_13_34 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_34 ) ,
    .I0 ( U1091.AB ) ,
    .I1 ( U1091.CD ) ,
    .I2 ( U1091.EF ) ) ;
and ( 
    .Z ( U1090.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_26 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1090.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_26 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1090.EF ) ,
    .I0 ( xor_decoded_masks_13_26 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_26 ) ,
    .I0 ( U1090.AB ) ,
    .I1 ( U1090.CD ) ,
    .I2 ( U1090.EF ) ) ;
and ( 
    .Z ( U599.AB ) ,
    .I0 ( masks_hold_reg_4_6 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U599.CD ) ,
    .I0 ( config1_xor_encoded_masks_47 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_47 ) ,
    .I0 ( U599.AB ) ,
    .I1 ( U599.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_8_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_10.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_10 ) ,
    .IN ( masks_hold_reg_8_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_10.QT ) ,
    .I1 ( masks_hold_reg_8_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_10.ED ) ,
    .S ( masks_hold_reg_8_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_10.ED ) ,
    .I1 ( masks_hold_reg_8_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_10.QT ) ) ;
and ( 
    .Z ( U1093.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_22 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1093.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_22 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1093.EF ) ,
    .I0 ( xor_decoded_masks_13_22 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_22 ) ,
    .I0 ( U1093.AB ) ,
    .I1 ( U1093.CD ) ,
    .I2 ( U1093.EF ) ) ;
and ( 
    .Z ( U598.AB ) ,
    .I0 ( n92 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U598.CD ) ,
    .I0 ( config1_xor_encoded_masks_44 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_44 ) ,
    .I0 ( U598.AB ) ,
    .I1 ( U598.CD ) ) ;
and ( 
    .Z ( U1092.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_38 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1092.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_38 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1092.EF ) ,
    .I0 ( xor_decoded_masks_13_38 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_38 ) ,
    .I0 ( U1092.AB ) ,
    .I1 ( U1092.CD ) ,
    .I2 ( U1092.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_5_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_9.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29283 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_9.CD ) ,
    .IN ( masks_shift_reg_5_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_24 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_25 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_24 ) ,
    .Q ( masks_shift_reg_5_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_25 ) ) ;
DFF masks_shift_reg_5_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_8.DI_ ) ,
    .IN ( n48 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay1941 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_8.CDNI_ ) ,
    .IN ( masks_shift_reg_5_9 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_8.CD ) ,
    .IN ( masks_shift_reg_5_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_8 ) ) ;
and ( 
    .Z ( U591.AB ) ,
    .I0 ( masks_hold_reg_1_5 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U591.CD ) ,
    .I0 ( config1_xor_encoded_masks_15 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_15 ) ,
    .I0 ( U591.AB ) ,
    .I1 ( U591.CD ) ) ;
and ( 
    .Z ( U590.AB ) ,
    .I0 ( masks_hold_reg_13_4 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U590.CD ) ,
    .I0 ( config1_xor_encoded_masks_145 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_145 ) ,
    .I0 ( U590.AB ) ,
    .I1 ( U590.CD ) ) ;
and ( 
    .Z ( U593.AB ) ,
    .I0 ( masks_hold_reg_0_8 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U593.CD ) ,
    .I0 ( config1_xor_encoded_masks_1 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_1 ) ,
    .I0 ( U593.AB ) ,
    .I1 ( U593.CD ) ) ;
and ( 
    .Z ( U809.AB ) ,
    .I0 ( masks_hold_reg_3_9 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U809.CD ) ,
    .I0 ( config1_xor_encoded_masks_33 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_33 ) ,
    .I0 ( U809.AB ) ,
    .I1 ( U809.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_5_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_5.CD ) ,
    .IN ( masks_shift_reg_5_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_5 ) ) ;
and ( 
    .Z ( U592.AB ) ,
    .I0 ( masks_hold_reg_9_5 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U592.CD ) ,
    .I0 ( config1_xor_encoded_masks_103 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_103 ) ,
    .I0 ( U592.AB ) ,
    .I1 ( U592.CD ) ) ;
and ( 
    .Z ( U808.AB ) ,
    .I0 ( masks_hold_reg_10_6 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U808.CD ) ,
    .I0 ( config1_xor_encoded_masks_113 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_113 ) ,
    .I0 ( U808.AB ) ,
    .I1 ( U808.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_5_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_4.CD ) ,
    .IN ( masks_shift_reg_5_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_24 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_25 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_24 ) ,
    .Q ( masks_shift_reg_5_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_25 ) ) ;
DFF masks_shift_reg_5_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_4 ) ) ;
and ( 
    .Z ( U595.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_85 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U595.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_32 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U595.EF ) ,
    .I0 ( xor_decoded_masks_8_32 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_32 ) ,
    .I0 ( U595.AB ) ,
    .I1 ( U595.CD ) ,
    .I2 ( U595.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_5_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_7.CD ) ,
    .IN ( masks_shift_reg_5_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_7 ) ) ;
and ( 
    .Z ( U594.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_117 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U594.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_10 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U594.EF ) ,
    .I0 ( xor_decoded_masks_2_10 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_10 ) ,
    .I0 ( U594.AB ) ,
    .I1 ( U594.CD ) ,
    .I2 ( U594.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_5_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_6.CD ) ,
    .IN ( masks_shift_reg_5_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_6 ) ) ;
and ( 
    .Z ( U597.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_68 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U597.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_14 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U597.EF ) ,
    .I0 ( xor_decoded_masks_1_14 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_14 ) ,
    .I0 ( U597.AB ) ,
    .I1 ( U597.CD ) ,
    .I2 ( U597.EF ) ) ;
and ( 
    .Z ( U805.AB ) ,
    .I0 ( masks_hold_reg_10_1 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U805.CD ) ,
    .I0 ( config1_xor_encoded_masks_118 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_118 ) ,
    .I0 ( U805.AB ) ,
    .I1 ( U805.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_5_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_1.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29283 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_1.CD ) ,
    .IN ( masks_shift_reg_5_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_1 ) ) ;
and ( 
    .Z ( U596.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_77 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U596.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_24 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U596.EF ) ,
    .I0 ( xor_decoded_masks_10_24 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_24 ) ,
    .I0 ( U596.AB ) ,
    .I1 ( U596.CD ) ,
    .I2 ( U596.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_5_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_0.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29283 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_0.CD ) ,
    .IN ( masks_shift_reg_5_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_0 ) ) ;
and ( 
    .Z ( U807.AB ) ,
    .I0 ( masks_hold_reg_8_7 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U807.CD ) ,
    .I0 ( config1_xor_encoded_masks_90 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_90 ) ,
    .I0 ( U807.AB ) ,
    .I1 ( U807.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_5_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_3.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29283 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_3.CD ) ,
    .IN ( masks_shift_reg_5_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_3 ) ) ;
and ( 
    .Z ( U806.AB ) ,
    .I0 ( masks_hold_reg_12_8 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U806.CD ) ,
    .I0 ( config1_xor_encoded_masks_133 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_133 ) ,
    .I0 ( U806.AB ) ,
    .I1 ( U806.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_5_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_2.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29283 ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_2.CD ) ,
    .IN ( masks_shift_reg_5_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_5_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_5_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_5_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_5_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_5_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_5_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_5_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_5_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_5_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_5_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_5_2 ) ) ;
and ( 
    .Z ( U801.AB ) ,
    .I0 ( masks_hold_reg_5_6 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U801.CD ) ,
    .I0 ( config1_xor_encoded_masks_58 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_58 ) ,
    .I0 ( U801.AB ) ,
    .I1 ( U801.CD ) ) ;
and ( 
    .Z ( U800.AB ) ,
    .I0 ( masks_hold_reg_3_4 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U800.CD ) ,
    .I0 ( config1_xor_encoded_masks_38 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_38 ) ,
    .I0 ( U800.AB ) ,
    .I1 ( U800.CD ) ) ;
and ( 
    .Z ( U803.AB ) ,
    .I0 ( masks_hold_reg_9_10 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U803.CD ) ,
    .I0 ( config1_xor_encoded_masks_98 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_98 ) ,
    .I0 ( U803.AB ) ,
    .I1 ( U803.CD ) ) ;
and ( 
    .Z ( U802.AB ) ,
    .I0 ( masks_hold_reg_7_8 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U802.CD ) ,
    .I0 ( config1_xor_encoded_masks_78 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_78 ) ,
    .I0 ( U802.AB ) ,
    .I1 ( U802.CD ) ) ;
and ( 
    .Z ( U1088.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_65 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1088.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_12 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1088.EF ) ,
    .I0 ( xor_decoded_masks_12_12 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_12 ) ,
    .I0 ( U1088.AB ) ,
    .I1 ( U1088.CD ) ,
    .I2 ( U1088.EF ) ) ;
and ( 
    .Z ( U1089.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_71 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1089.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_18 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1089.EF ) ,
    .I0 ( xor_decoded_masks_12_18 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_18 ) ,
    .I0 ( U1089.AB ) ,
    .I1 ( U1089.CD ) ,
    .I2 ( U1089.EF ) ) ;
and ( 
    .Z ( U1084.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_8 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1084.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_8 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1084.EF ) ,
    .I0 ( xor_decoded_masks_11_8 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_8 ) ,
    .I0 ( U1084.AB ) ,
    .I1 ( U1084.CD ) ,
    .I2 ( U1084.EF ) ) ;
and ( 
    .Z ( U1085.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_12 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1085.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_12 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1085.EF ) ,
    .I0 ( xor_decoded_masks_11_12 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_12 ) ,
    .I0 ( U1085.AB ) ,
    .I1 ( U1085.CD ) ,
    .I2 ( U1085.EF ) ) ;
and ( 
    .Z ( U1086.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_79 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1086.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_26 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1086.EF ) ,
    .I0 ( xor_decoded_masks_12_26 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_26 ) ,
    .I0 ( U1086.AB ) ,
    .I1 ( U1086.CD ) ,
    .I2 ( U1086.EF ) ) ;
and ( 
    .Z ( U1087.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_61 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1087.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_8 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1087.EF ) ,
    .I0 ( xor_decoded_masks_12_8 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_8 ) ,
    .I0 ( U1087.AB ) ,
    .I1 ( U1087.CD ) ,
    .I2 ( U1087.EF ) ) ;
and ( 
    .Z ( U1081.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_34 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1081.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_34 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1081.EF ) ,
    .I0 ( xor_decoded_masks_11_34 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_34 ) ,
    .I0 ( U1081.AB ) ,
    .I1 ( U1081.CD ) ,
    .I2 ( U1081.EF ) ) ;
and ( 
    .Z ( U1082.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_38 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1082.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_38 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1082.EF ) ,
    .I0 ( xor_decoded_masks_11_38 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_38 ) ,
    .I0 ( U1082.AB ) ,
    .I1 ( U1082.CD ) ,
    .I2 ( U1082.EF ) ) ;
and ( 
    .Z ( U1083.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_22 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1083.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_22 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1083.EF ) ,
    .I0 ( xor_decoded_masks_11_22 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_22 ) ,
    .I0 ( U1083.AB ) ,
    .I1 ( U1083.CD ) ,
    .I2 ( U1083.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_10.DI_ ) ,
    .IN ( N179 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_0_1 ) ) ;
DFF masks_shift_reg_7_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_7_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_7_10 ) ) ;
and ( 
    .Z ( U489.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_49 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U489.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_49 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U489.EF ) ,
    .I0 ( xor_decoded_masks_0_49 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_49 ) ,
    .I0 ( U489.AB ) ,
    .I1 ( U489.CD ) ,
    .I2 ( U489.EF ) ) ;
and ( 
    .Z ( U488.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_56 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U488.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_2 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U488.EF ) ,
    .I0 ( xor_decoded_masks_1_2 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_2 ) ,
    .I0 ( U488.AB ) ,
    .I1 ( U488.CD ) ,
    .I2 ( U488.EF ) ) ;
and ( 
    .Z ( U682.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_79 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U682.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_26 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U682.EF ) ,
    .I0 ( xor_decoded_masks_8_26 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_26 ) ,
    .I0 ( U682.AB ) ,
    .I1 ( U682.CD ) ,
    .I2 ( U682.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_1_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_5.CD ) ,
    .IN ( masks_shift_reg_1_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_5 ) ) ;
and ( 
    .Z ( U681.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_87 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U681.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_34 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U681.EF ) ,
    .I0 ( xor_decoded_masks_8_34 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_34 ) ,
    .I0 ( U681.AB ) ,
    .I1 ( U681.CD ) ,
    .I2 ( U681.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_1_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_4.CD ) ,
    .IN ( masks_shift_reg_1_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_4 ) ) ;
and ( 
    .Z ( U680.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_71 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U680.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_18 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U680.EF ) ,
    .I0 ( xor_decoded_masks_6_18 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_18 ) ,
    .I0 ( U680.AB ) ,
    .I1 ( U680.CD ) ,
    .I2 ( U680.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_1_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_7.CD ) ,
    .IN ( masks_shift_reg_1_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_7 ) ) ;
and ( 
    .Z ( U687.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_91 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U687.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_38 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U687.EF ) ,
    .I0 ( xor_decoded_masks_10_38 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_38 ) ,
    .I0 ( U687.AB ) ,
    .I1 ( U687.CD ) ,
    .I2 ( U687.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_1_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_6.CD ) ,
    .IN ( masks_shift_reg_1_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_6 ) ) ;
and ( 
    .Z ( U686.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_87 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U686.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_34 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U686.EF ) ,
    .I0 ( xor_decoded_masks_10_34 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_34 ) ,
    .I0 ( U686.AB ) ,
    .I1 ( U686.CD ) ,
    .I2 ( U686.EF ) ) ;
and ( 
    .Z ( U988.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_32 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U988.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_32 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U988.EF ) ,
    .I0 ( xor_decoded_masks_3_32 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_32 ) ,
    .I0 ( U988.AB ) ,
    .I1 ( U988.CD ) ,
    .I2 ( U988.EF ) ) ;
and ( 
    .Z ( U685.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_71 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U685.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_18 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U685.EF ) ,
    .I0 ( xor_decoded_masks_8_18 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_18 ) ,
    .I0 ( U685.AB ) ,
    .I1 ( U685.CD ) ,
    .I2 ( U685.EF ) ) ;
and ( 
    .Z ( U989.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_24 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U989.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_24 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U989.EF ) ,
    .I0 ( xor_decoded_masks_3_24 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_24 ) ,
    .I0 ( U989.AB ) ,
    .I1 ( U989.CD ) ,
    .I2 ( U989.EF ) ) ;
and ( 
    .Z ( U684.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_65 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U684.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_12 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U684.EF ) ,
    .I0 ( xor_decoded_masks_8_12 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_12 ) ,
    .I0 ( U684.AB ) ,
    .I1 ( U684.CD ) ,
    .I2 ( U684.EF ) ) ;
and ( 
    .Z ( U995.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_63 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U995.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_10 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U995.EF ) ,
    .I0 ( xor_decoded_masks_4_10 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_10 ) ,
    .I0 ( U995.AB ) ,
    .I1 ( U995.CD ) ,
    .I2 ( U995.EF ) ) ;
and ( 
    .Z ( U698.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_66 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U698.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_12 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U698.EF ) ,
    .I0 ( xor_decoded_masks_1_12 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_12 ) ,
    .I0 ( U698.AB ) ,
    .I1 ( U698.CD ) ,
    .I2 ( U698.EF ) ) ;
and ( 
    .Z ( U994.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_10 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U994.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_10 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U994.EF ) ,
    .I0 ( xor_decoded_masks_3_10 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_10 ) ,
    .I0 ( U994.AB ) ,
    .I1 ( U994.CD ) ,
    .I2 ( U994.EF ) ) ;
and ( 
    .Z ( U699.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_41 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U699.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_41 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U699.EF ) ,
    .I0 ( xor_decoded_masks_0_41 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_41 ) ,
    .I0 ( U699.AB ) ,
    .I1 ( U699.CD ) ,
    .I2 ( U699.EF ) ) ;
and ( 
    .Z ( U997.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_24 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U997.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_24 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U997.EF ) ,
    .I0 ( xor_decoded_masks_5_24 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_24 ) ,
    .I0 ( U997.AB ) ,
    .I1 ( U997.CD ) ,
    .I2 ( U997.EF ) ) ;
and ( 
    .Z ( U996.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_69 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U996.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_16 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U996.EF ) ,
    .I0 ( xor_decoded_masks_4_16 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_16 ) ,
    .I0 ( U996.AB ) ,
    .I1 ( U996.CD ) ,
    .I2 ( U996.EF ) ) ;
and ( 
    .Z ( U991.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_36 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U991.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_36 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U991.EF ) ,
    .I0 ( xor_decoded_masks_3_36 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_36 ) ,
    .I0 ( U991.AB ) ,
    .I1 ( U991.CD ) ,
    .I2 ( U991.EF ) ) ;
and ( 
    .Z ( U990.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_28 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U990.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_28 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U990.EF ) ,
    .I0 ( xor_decoded_masks_3_28 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_28 ) ,
    .I0 ( U990.AB ) ,
    .I1 ( U990.CD ) ,
    .I2 ( U990.EF ) ) ;
and ( 
    .Z ( U993.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_16 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U993.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_16 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U993.EF ) ,
    .I0 ( xor_decoded_masks_3_16 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_16 ) ,
    .I0 ( U993.AB ) ,
    .I1 ( U993.CD ) ,
    .I2 ( U993.EF ) ) ;
and ( 
    .Z ( U692.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_91 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U692.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_38 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U692.EF ) ,
    .I0 ( xor_decoded_masks_14_38 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_38 ) ,
    .I0 ( U692.AB ) ,
    .I1 ( U692.CD ) ,
    .I2 ( U692.EF ) ) ;
and ( 
    .Z ( U992.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_14 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U992.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_14 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U992.EF ) ,
    .I0 ( xor_decoded_masks_3_14 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_14 ) ,
    .I0 ( U992.AB ) ,
    .I1 ( U992.CD ) ,
    .I2 ( U992.EF ) ) ;
and ( 
    .Z ( U693.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_80 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U693.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_26 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U693.EF ) ,
    .I0 ( xor_decoded_masks_1_26 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_26 ) ,
    .I0 ( U693.AB ) ,
    .I1 ( U693.CD ) ,
    .I2 ( U693.EF ) ) ;
and ( 
    .Z ( U690.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_87 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U690.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_34 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U690.EF ) ,
    .I0 ( xor_decoded_masks_14_34 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_34 ) ,
    .I0 ( U690.AB ) ,
    .I1 ( U690.CD ) ,
    .I2 ( U690.EF ) ) ;
and ( 
    .Z ( U691.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_79 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U691.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_26 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U691.EF ) ,
    .I0 ( xor_decoded_masks_14_26 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_26 ) ,
    .I0 ( U691.AB ) ,
    .I1 ( U691.CD ) ,
    .I2 ( U691.EF ) ) ;
and ( 
    .Z ( U696.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_62 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U696.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_8 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U696.EF ) ,
    .I0 ( xor_decoded_masks_1_8 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_8 ) ,
    .I0 ( U696.AB ) ,
    .I1 ( U696.CD ) ,
    .I2 ( U696.EF ) ) ;
and ( 
    .Z ( U697.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_76 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U697.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_22 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U697.EF ) ,
    .I0 ( xor_decoded_masks_1_22 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_22 ) ,
    .I0 ( U697.AB ) ,
    .I1 ( U697.CD ) ,
    .I2 ( U697.EF ) ) ;
and ( 
    .Z ( U999.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_36 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U999.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_36 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U999.EF ) ,
    .I0 ( xor_decoded_masks_5_36 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_36 ) ,
    .I0 ( U999.AB ) ,
    .I1 ( U999.CD ) ,
    .I2 ( U999.EF ) ) ;
and ( 
    .Z ( U694.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_88 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U694.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_34 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U694.EF ) ,
    .I0 ( xor_decoded_masks_1_34 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_34 ) ,
    .I0 ( U694.AB ) ,
    .I1 ( U694.CD ) ,
    .I2 ( U694.EF ) ) ;
and ( 
    .Z ( U998.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_32 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U998.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_32 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U998.EF ) ,
    .I0 ( xor_decoded_masks_5_32 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_32 ) ,
    .I0 ( U998.AB ) ,
    .I1 ( U998.CD ) ,
    .I2 ( U998.EF ) ) ;
and ( 
    .Z ( U695.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_92 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U695.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_38 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U695.EF ) ,
    .I0 ( xor_decoded_masks_1_38 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_38 ) ,
    .I0 ( U695.AB ) ,
    .I1 ( U695.CD ) ,
    .I2 ( U695.EF ) ) ;
and ( 
    .Z ( U885.AB ) ,
    .I0 ( masks_hold_reg_12_9 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U885.CD ) ,
    .I0 ( config1_xor_encoded_masks_132 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_132 ) ,
    .I0 ( U885.AB ) ,
    .I1 ( U885.CD ) ) ;
and ( 
    .Z ( U887.AB ) ,
    .I0 ( masks_hold_reg_3_8 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U887.CD ) ,
    .I0 ( config1_xor_encoded_masks_34 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_34 ) ,
    .I0 ( U887.AB ) ,
    .I1 ( U887.CD ) ) ;
and ( 
    .Z ( U886.AB ) ,
    .I0 ( masks_hold_reg_0_9 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U886.CD ) ,
    .I0 ( config1_xor_encoded_masks_0 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_0 ) ,
    .I0 ( U886.AB ) ,
    .I1 ( U886.CD ) ) ;
and ( 
    .Z ( U881.AB ) ,
    .I0 ( masks_hold_reg_11_0 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U881.CD ) ,
    .I0 ( config1_xor_encoded_masks_130 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_130 ) ,
    .I0 ( U881.AB ) ,
    .I1 ( U881.CD ) ) ;
and ( 
    .Z ( U880.AB ) ,
    .I0 ( masks_hold_reg_2_1 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U880.CD ) ,
    .I0 ( config1_xor_encoded_masks_30 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_30 ) ,
    .I0 ( U880.AB ) ,
    .I1 ( U880.CD ) ) ;
and ( 
    .Z ( U883.AB ) ,
    .I0 ( masks_hold_reg_11_10 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U883.CD ) ,
    .I0 ( config1_xor_encoded_masks_120 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_120 ) ,
    .I0 ( U883.AB ) ,
    .I1 ( U883.CD ) ) ;
and ( 
    .Z ( U811.AB ) ,
    .I0 ( masks_hold_reg_6_2 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U811.CD ) ,
    .I0 ( config1_xor_encoded_masks_73 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_73 ) ,
    .I0 ( U811.AB ) ,
    .I1 ( U811.CD ) ) ;
and ( 
    .Z ( U482.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_55 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U482.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_2 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U482.EF ) ,
    .I0 ( xor_decoded_masks_14_2 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_2 ) ,
    .I0 ( U482.AB ) ,
    .I1 ( U482.CD ) ,
    .I2 ( U482.EF ) ) ;
and ( 
    .Z ( U812.AB ) ,
    .I0 ( masks_hold_reg_8_4 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U812.CD ) ,
    .I0 ( config1_xor_encoded_masks_93 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_93 ) ,
    .I0 ( U812.AB ) ,
    .I1 ( U812.CD ) ) ;
and ( 
    .Z ( U485.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_60 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U485.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_6 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U485.EF ) ,
    .I0 ( xor_decoded_masks_1_6 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_6 ) ,
    .I0 ( U485.AB ) ,
    .I1 ( U485.CD ) ,
    .I2 ( U485.EF ) ) ;
and ( 
    .Z ( U813.AB ) ,
    .I0 ( masks_hold_reg_1_7 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U813.CD ) ,
    .I0 ( config1_xor_encoded_masks_13 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_13 ) ,
    .I0 ( U813.AB ) ,
    .I1 ( U813.CD ) ) ;
and ( 
    .Z ( U484.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_61 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U484.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_7 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U484.EF ) ,
    .I0 ( xor_decoded_masks_1_7 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_7 ) ,
    .I0 ( U484.AB ) ,
    .I1 ( U484.CD ) ,
    .I2 ( U484.EF ) ) ;
and ( 
    .Z ( U487.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_57 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U487.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_3 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U487.EF ) ,
    .I0 ( xor_decoded_masks_1_3 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_3 ) ,
    .I0 ( U487.AB ) ,
    .I1 ( U487.CD ) ,
    .I2 ( U487.EF ) ) ;
and ( 
    .Z ( U486.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_54 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U486.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_0 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U486.EF ) ,
    .I0 ( xor_decoded_masks_1_0 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_0 ) ,
    .I0 ( U486.AB ) ,
    .I1 ( U486.CD ) ,
    .I2 ( U486.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_12_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_4 ) ,
    .IN ( masks_hold_reg_12_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_4.QT ) ,
    .I1 ( masks_hold_reg_12_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_4.ED ) ,
    .S ( masks_hold_reg_12_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_4.ED ) ,
    .I1 ( masks_hold_reg_12_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_4.QT ) ) ;
and ( 
    .Z ( U1198.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_9 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1198.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_9 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1198.EF ) ,
    .I0 ( xor_decoded_masks_5_9 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_9 ) ,
    .I0 ( U1198.AB ) ,
    .I1 ( U1198.CD ) ,
    .I2 ( U1198.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_12_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_5 ) ,
    .IN ( masks_hold_reg_12_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_5.QT ) ,
    .I1 ( masks_hold_reg_12_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_5.ED ) ,
    .S ( masks_hold_reg_12_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_5.ED ) ,
    .I1 ( masks_hold_reg_12_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_5.QT ) ) ;
and ( 
    .Z ( U1199.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_13 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1199.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_13 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1199.EF ) ,
    .I0 ( xor_decoded_masks_5_13 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_13 ) ,
    .I0 ( U1199.AB ) ,
    .I1 ( U1199.CD ) ,
    .I2 ( U1199.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_12_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_6 ) ,
    .IN ( masks_hold_reg_12_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_6.QT ) ,
    .I1 ( masks_hold_reg_12_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_6.ED ) ,
    .S ( masks_hold_reg_12_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_6.ED ) ,
    .I1 ( masks_hold_reg_12_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_12_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_7 ) ,
    .IN ( masks_hold_reg_12_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_7.QT ) ,
    .I1 ( masks_hold_reg_12_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_7.ED ) ,
    .S ( masks_hold_reg_12_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_7.ED ) ,
    .I1 ( masks_hold_reg_12_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_12_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_9.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_9.CD ) ,
    .IN ( masks_shift_reg_12_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_12_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_0 ) ,
    .IN ( masks_hold_reg_12_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_0.QT ) ,
    .I1 ( masks_hold_reg_12_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_0.ED ) ,
    .S ( masks_hold_reg_12_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_0.ED ) ,
    .I1 ( masks_hold_reg_12_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_0.QT ) ) ;
and ( 
    .Z ( U1194.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_27 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1194.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_27 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1194.EF ) ,
    .I0 ( xor_decoded_masks_5_27 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_27 ) ,
    .I0 ( U1194.AB ) ,
    .I1 ( U1194.CD ) ,
    .I2 ( U1194.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_8.DI_ ) ,
    .IN ( n67 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_8.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_8.CD ) ,
    .IN ( masks_shift_reg_12_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_12_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_1 ) ,
    .IN ( masks_hold_reg_12_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_1.QT ) ,
    .I1 ( masks_hold_reg_12_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_1.ED ) ,
    .S ( masks_hold_reg_12_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_1.ED ) ,
    .I1 ( masks_hold_reg_12_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_1.QT ) ) ;
and ( 
    .Z ( U1195.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_35 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1195.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_35 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1195.EF ) ,
    .I0 ( xor_decoded_masks_5_35 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_35 ) ,
    .I0 ( U1195.AB ) ,
    .I1 ( U1195.CD ) ,
    .I2 ( U1195.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_12_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_2 ) ,
    .IN ( masks_hold_reg_12_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_2.QT ) ,
    .I1 ( masks_hold_reg_12_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_2.ED ) ,
    .S ( masks_hold_reg_12_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_2.ED ) ,
    .I1 ( masks_hold_reg_12_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_2.QT ) ) ;
and ( 
    .Z ( U1196.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_39 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1196.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_39 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1196.EF ) ,
    .I0 ( xor_decoded_masks_5_39 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_39 ) ,
    .I0 ( U1196.AB ) ,
    .I1 ( U1196.CD ) ,
    .I2 ( U1196.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_12_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_3 ) ,
    .IN ( masks_hold_reg_12_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_3.QT ) ,
    .I1 ( masks_hold_reg_12_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_3.ED ) ,
    .S ( masks_hold_reg_12_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_3.ED ) ,
    .I1 ( masks_hold_reg_12_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_3.QT ) ) ;
and ( 
    .Z ( U1197.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_23 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1197.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_23 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1197.EF ) ,
    .I0 ( xor_decoded_masks_5_23 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_23 ) ,
    .I0 ( U1197.AB ) ,
    .I1 ( U1197.CD ) ,
    .I2 ( U1197.EF ) ) ;
and ( 
    .Z ( U1190.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_9 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1190.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_9 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1190.EF ) ,
    .I0 ( xor_decoded_masks_3_9 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_9 ) ,
    .I0 ( U1190.AB ) ,
    .I1 ( U1190.CD ) ,
    .I2 ( U1190.EF ) ) ;
and ( 
    .Z ( U1191.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_19 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1191.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_19 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1191.EF ) ,
    .I0 ( xor_decoded_masks_3_19 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_19 ) ,
    .I0 ( U1191.AB ) ,
    .I1 ( U1191.CD ) ,
    .I2 ( U1191.EF ) ) ;
and ( 
    .Z ( U498.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_15 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U498.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_15 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U498.EF ) ,
    .I0 ( xor_decoded_masks_0_15 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_15 ) ,
    .I0 ( U498.AB ) ,
    .I1 ( U498.CD ) ,
    .I2 ( U498.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_12_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_3.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_3.CD ) ,
    .IN ( masks_shift_reg_12_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_3 ) ) ;
and ( 
    .Z ( U1192.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_13 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1192.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_13 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1192.EF ) ,
    .I0 ( xor_decoded_masks_3_13 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_13 ) ,
    .I0 ( U1192.AB ) ,
    .I1 ( U1192.CD ) ,
    .I2 ( U1192.EF ) ) ;
and ( 
    .Z ( U499.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_14 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U499.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_14 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U499.EF ) ,
    .I0 ( xor_decoded_masks_0_14 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_14 ) ,
    .I0 ( U499.AB ) ,
    .I1 ( U499.CD ) ,
    .I2 ( U499.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_12_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_2.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_2.CD ) ,
    .IN ( masks_shift_reg_12_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_2 ) ) ;
and ( 
    .Z ( U1193.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_72 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1193.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_19 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1193.EF ) ,
    .I0 ( xor_decoded_masks_4_19 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_19 ) ,
    .I0 ( U1193.AB ) ,
    .I1 ( U1193.CD ) ,
    .I2 ( U1193.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_12_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_1.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_1.CD ) ,
    .IN ( masks_shift_reg_12_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_12_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_8.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_8 ) ,
    .IN ( masks_hold_reg_12_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_8.QT ) ,
    .I1 ( masks_hold_reg_12_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_8.ED ) ,
    .S ( masks_hold_reg_12_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_8.ED ) ,
    .I1 ( masks_hold_reg_12_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_12_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_0.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_0.CD ) ,
    .IN ( masks_shift_reg_12_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_12_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_9.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_9 ) ,
    .IN ( masks_hold_reg_12_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_9.QT ) ,
    .I1 ( masks_hold_reg_12_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_9.ED ) ,
    .S ( masks_hold_reg_12_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_9.ED ) ,
    .I1 ( masks_hold_reg_12_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_9.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_7.DI_ ) ,
    .IN ( n42 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_7.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_7.CD ) ,
    .IN ( masks_shift_reg_12_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_6.DI_ ) ,
    .IN ( n46 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_6.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_6.CD ) ,
    .IN ( masks_shift_reg_12_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_12_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_5.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_5.CD ) ,
    .IN ( masks_shift_reg_12_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_12_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_4.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_4.CD ) ,
    .IN ( masks_shift_reg_12_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_12_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_12_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_12_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_12_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_12_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_12_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_12_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_12_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_12_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_12_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_12_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_12_4 ) ) ;
and ( 
    .Z ( U490.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_48 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U490.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_48 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U490.EF ) ,
    .I0 ( xor_decoded_masks_0_48 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_48 ) ,
    .I0 ( U490.AB ) ,
    .I1 ( U490.CD ) ,
    .I2 ( U490.EF ) ) ;
and ( 
    .Z ( U491.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_10 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U491.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_10 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U491.EF ) ,
    .I0 ( xor_decoded_masks_0_10 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_10 ) ,
    .I0 ( U491.AB ) ,
    .I1 ( U491.CD ) ,
    .I2 ( U491.EF ) ) ;
and ( 
    .Z ( U492.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_12 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U492.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_12 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U492.EF ) ,
    .I0 ( xor_decoded_masks_0_12 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_12 ) ,
    .I0 ( U492.AB ) ,
    .I1 ( U492.CD ) ,
    .I2 ( U492.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_10.DI_ ) ,
    .IN ( N168 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2881 ) ) ;
DFF masks_shift_reg_6_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_6_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_6_10 ) ) ;
and ( 
    .Z ( U493.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_13 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U493.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_13 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U493.EF ) ,
    .I0 ( xor_decoded_masks_0_13 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_13 ) ,
    .I0 ( U493.AB ) ,
    .I1 ( U493.CD ) ,
    .I2 ( U493.EF ) ) ;
and ( 
    .Z ( U494.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_3 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U494.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_3 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U494.EF ) ,
    .I0 ( xor_decoded_masks_0_3 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_3 ) ,
    .I0 ( U494.AB ) ,
    .I1 ( U494.CD ) ,
    .I2 ( U494.EF ) ) ;
and ( 
    .Z ( U495.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_0 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U495.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_0 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U495.EF ) ,
    .I0 ( xor_decoded_masks_0_0 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_0 ) ,
    .I0 ( U495.AB ) ,
    .I1 ( U495.CD ) ,
    .I2 ( U495.EF ) ) ;
and ( 
    .Z ( U496.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_2 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U496.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_2 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U496.EF ) ,
    .I0 ( xor_decoded_masks_0_2 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_2 ) ,
    .I0 ( U496.AB ) ,
    .I1 ( U496.CD ) ,
    .I2 ( U496.EF ) ) ;
and ( 
    .Z ( U497.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_8 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U497.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_8 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U497.EF ) ,
    .I0 ( xor_decoded_masks_0_8 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_8 ) ,
    .I0 ( U497.AB ) ,
    .I1 ( U497.CD ) ,
    .I2 ( U497.EF ) ) ;
and ( 
    .Z ( U1189.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_39 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1189.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_39 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1189.EF ) ,
    .I0 ( xor_decoded_masks_3_39 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_39 ) ,
    .I0 ( U1189.AB ) ,
    .I1 ( U1189.CD ) ,
    .I2 ( U1189.EF ) ) ;
and ( 
    .Z ( U1188.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_31 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1188.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_31 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1188.EF ) ,
    .I0 ( xor_decoded_masks_3_31 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_31 ) ,
    .I0 ( U1188.AB ) ,
    .I1 ( U1188.CD ) ,
    .I2 ( U1188.EF ) ) ;
and ( 
    .Z ( U1185.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_11 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1185.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_11 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1185.EF ) ,
    .I0 ( xor_decoded_masks_0_11 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_11 ) ,
    .I0 ( U1185.AB ) ,
    .I1 ( U1185.CD ) ,
    .I2 ( U1185.EF ) ) ;
and ( 
    .Z ( U1184.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_51 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1184.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_51 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1184.EF ) ,
    .I0 ( xor_decoded_masks_0_51 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_51 ) ,
    .I0 ( U1184.AB ) ,
    .I1 ( U1184.CD ) ,
    .I2 ( U1184.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_9_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_6.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_6 ) ,
    .IN ( masks_hold_reg_9_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_6.QT ) ,
    .I1 ( masks_hold_reg_9_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_6.ED ) ,
    .S ( masks_hold_reg_9_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_6.ED ) ,
    .I1 ( masks_hold_reg_9_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_6.QT ) ) ;
and ( 
    .Z ( U895.AB ) ,
    .I0 ( masks_hold_reg_8_6 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U895.CD ) ,
    .I0 ( config1_xor_encoded_masks_91 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_91 ) ,
    .I0 ( U895.AB ) ,
    .I1 ( U895.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_9_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_7.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_7 ) ,
    .IN ( masks_hold_reg_9_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_7.QT ) ,
    .I1 ( masks_hold_reg_9_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_7.ED ) ,
    .S ( masks_hold_reg_9_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_7.ED ) ,
    .I1 ( masks_hold_reg_9_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_7.QT ) ) ;
and ( 
    .Z ( U896.AB ) ,
    .I0 ( masks_hold_reg_10_8 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U896.CD ) ,
    .I0 ( config1_xor_encoded_masks_111 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_111 ) ,
    .I0 ( U896.AB ) ,
    .I1 ( U896.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_9_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_4.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_4 ) ,
    .IN ( masks_hold_reg_9_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_4.QT ) ,
    .I1 ( masks_hold_reg_9_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_4.ED ) ,
    .S ( masks_hold_reg_9_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_4.ED ) ,
    .I1 ( masks_hold_reg_9_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_4.QT ) ) ;
and ( 
    .Z ( U897.AB ) ,
    .I0 ( masks_hold_reg_3_1 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U897.CD ) ,
    .I0 ( config1_xor_encoded_masks_41 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_41 ) ,
    .I0 ( U897.AB ) ,
    .I1 ( U897.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_9_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_5.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_5 ) ,
    .IN ( masks_hold_reg_9_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_5.QT ) ,
    .I1 ( masks_hold_reg_9_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_5.ED ) ,
    .S ( masks_hold_reg_9_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_5.ED ) ,
    .I1 ( masks_hold_reg_9_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_5.QT ) ) ;
and ( 
    .Z ( U890.AB ) ,
    .I0 ( masks_hold_reg_8_3 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U890.CD ) ,
    .I0 ( config1_xor_encoded_masks_94 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_94 ) ,
    .I0 ( U890.AB ) ,
    .I1 ( U890.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_9_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_2.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_2 ) ,
    .IN ( masks_hold_reg_9_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_2.QT ) ,
    .I1 ( masks_hold_reg_9_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_2.ED ) ,
    .S ( masks_hold_reg_9_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_2.ED ) ,
    .I1 ( masks_hold_reg_9_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_2.QT ) ) ;
and ( 
    .Z ( U891.AB ) ,
    .I0 ( masks_hold_reg_12_7 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U891.CD ) ,
    .I0 ( config1_xor_encoded_masks_134 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_134 ) ,
    .I0 ( U891.AB ) ,
    .I1 ( U891.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_9_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_3.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_3 ) ,
    .IN ( masks_hold_reg_9_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_3.QT ) ,
    .I1 ( masks_hold_reg_9_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_3.ED ) ,
    .S ( masks_hold_reg_9_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_3.ED ) ,
    .I1 ( masks_hold_reg_9_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_3.QT ) ) ;
and ( 
    .Z ( U892.AB ) ,
    .I0 ( masks_hold_reg_10_5 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U892.CD ) ,
    .I0 ( config1_xor_encoded_masks_114 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_114 ) ,
    .I0 ( U892.AB ) ,
    .I1 ( U892.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_9_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_0.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_0 ) ,
    .IN ( masks_hold_reg_9_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_0.QT ) ,
    .I1 ( masks_hold_reg_9_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_0.ED ) ,
    .S ( masks_hold_reg_9_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_0.ED ) ,
    .I1 ( masks_hold_reg_9_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_0.QT ) ) ;
and ( 
    .Z ( U893.AB ) ,
    .I0 ( masks_hold_reg_0_7 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U893.CD ) ,
    .I0 ( config1_xor_encoded_masks_2 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_2 ) ,
    .I0 ( U893.AB ) ,
    .I1 ( U893.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_9_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_1.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_1 ) ,
    .IN ( masks_hold_reg_9_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_1.QT ) ,
    .I1 ( masks_hold_reg_9_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_1.ED ) ,
    .S ( masks_hold_reg_9_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_1.ED ) ,
    .I1 ( masks_hold_reg_9_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_1.QT ) ) ;
and ( 
    .Z ( U898.AB ) ,
    .I0 ( masks_hold_reg_5_3 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U898.CD ) ,
    .I0 ( config1_xor_encoded_masks_61 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_61 ) ,
    .I0 ( U898.AB ) ,
    .I1 ( U898.CD ) ) ;
and ( 
    .Z ( U899.AB ) ,
    .I0 ( masks_hold_reg_7_5 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U899.CD ) ,
    .I0 ( config1_xor_encoded_masks_81 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_81 ) ,
    .I0 ( U899.AB ) ,
    .I1 ( U899.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_7_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_0_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_reg_10.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_7_10 ) ,
    .IN ( masks_hold_reg_7_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_7_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_7_reg_10.QT ) ,
    .I1 ( masks_hold_reg_7_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_7_reg_10.ED ) ,
    .S ( masks_hold_reg_7_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_7_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_7_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_7_reg_10.ED ) ,
    .I1 ( masks_hold_reg_7_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_7_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_7_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_7_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_7_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_7_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_7_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_7_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_7_reg_10.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_3_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_10.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_10 ) ,
    .IN ( masks_hold_reg_3_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_10.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_3_reg_10.QT ) ,
    .I1 ( masks_hold_reg_3_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_10.ED ) ,
    .S ( masks_hold_reg_3_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_10.ED ) ,
    .I1 ( masks_hold_reg_3_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_3_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_3_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_10.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_8_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_0.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_0.CD ) ,
    .IN ( masks_shift_reg_8_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_8_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_1.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_1.CD ) ,
    .IN ( masks_shift_reg_8_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_8_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_2.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_2.CD ) ,
    .IN ( masks_shift_reg_8_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_8_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_3.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_3.CD ) ,
    .IN ( masks_shift_reg_8_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_8_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_4.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_4.CD ) ,
    .IN ( masks_shift_reg_8_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_8_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_5.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_5.CD ) ,
    .IN ( masks_shift_reg_8_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_8_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_6.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_6.CD ) ,
    .IN ( masks_shift_reg_8_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_7.DI_ ) ,
    .IN ( n93 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_7.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_7.CD ) ,
    .IN ( masks_shift_reg_8_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_8_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_8.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_8.CD ) ,
    .IN ( masks_shift_reg_8_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_2_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_8.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_8.CD ) ,
    .IN ( masks_shift_reg_2_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_8_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_9.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_9.CD ) ,
    .IN ( masks_shift_reg_8_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_8_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_8_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_8_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_8_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_8_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_8_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_8_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_8_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_8_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_8_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_8_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_2_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_9.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_9.CD ) ,
    .IN ( masks_shift_reg_2_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_2_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_2.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_2.CD ) ,
    .IN ( masks_shift_reg_2_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_2_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_3.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_3.CD ) ,
    .IN ( masks_shift_reg_2_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_2_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_0.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_0.CD ) ,
    .IN ( masks_shift_reg_2_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_2_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_1.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_1.CD ) ,
    .IN ( masks_shift_reg_2_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_2_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_6.CD ) ,
    .IN ( masks_shift_reg_2_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_2_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_7.CD ) ,
    .IN ( masks_shift_reg_2_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_2_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_4.CD ) ,
    .IN ( masks_shift_reg_2_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_2_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_2_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_5.CD ) ,
    .IN ( masks_shift_reg_2_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_2_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_2_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_2_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_2_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_2_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_2_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_2_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_2_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_2_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_2_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_2_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_2_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_10.DI_ ) ,
    .IN ( N113 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_10.CPI_ ) ,
    .IN ( edt_clock ) ) ;
DFF masks_shift_reg_1_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_1_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_1_10 ) ) ;
and ( 
    .Z ( U791.AB ) ,
    .I0 ( masks_hold_reg_0_0 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U791.CD ) ,
    .I0 ( n37 ) ,
    .I1 ( config1_xor_encoded_masks_9 ) ) ;
or ( 
    .Z ( xor_encoded_masks_9 ) ,
    .I0 ( U791.AB ) ,
    .I1 ( U791.CD ) ) ;
and ( 
    .Z ( U790.AB ) ,
    .I0 ( masks_hold_reg_10_9 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U790.CD ) ,
    .I0 ( config1_xor_encoded_masks_110 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_110 ) ,
    .I0 ( U790.AB ) ,
    .I1 ( U790.CD ) ) ;
and ( 
    .Z ( U797.AB ) ,
    .I0 ( masks_hold_reg_12_2 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U797.CD ) ,
    .I0 ( config1_xor_encoded_masks_139 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_139 ) ,
    .I0 ( U797.AB ) ,
    .I1 ( U797.CD ) ) ;
and ( 
    .Z ( U796.AB ) ,
    .I0 ( masks_hold_reg_9_9 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U796.CD ) ,
    .I0 ( config1_xor_encoded_masks_99 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_99 ) ,
    .I0 ( U796.AB ) ,
    .I1 ( U796.CD ) ) ;
and ( 
    .Z ( U795.AB ) ,
    .I0 ( masks_hold_reg_7_7 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U795.CD ) ,
    .I0 ( config1_xor_encoded_masks_79 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_79 ) ,
    .I0 ( U795.AB ) ,
    .I1 ( U795.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_10_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_9.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_9.CD ) ,
    .IN ( masks_shift_reg_10_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_9 ) ) ;
and ( 
    .Z ( U794.AB ) ,
    .I0 ( masks_hold_reg_5_5 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U794.CD ) ,
    .I0 ( config1_xor_encoded_masks_59 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_59 ) ,
    .I0 ( U794.AB ) ,
    .I1 ( U794.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_10_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_8.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_8.CD ) ,
    .IN ( masks_shift_reg_10_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_10_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_1.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_1.CD ) ,
    .IN ( masks_shift_reg_10_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_3.DI_ ) ,
    .IN ( n83 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_3.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_3 ) ,
    .IN ( masks_hold_reg_4_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_3.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_4_reg_3.QT ) ,
    .I1 ( masks_hold_reg_4_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_3.ED ) ,
    .S ( masks_hold_reg_4_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_3.ED ) ,
    .I1 ( masks_hold_reg_4_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_4_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_4_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_10_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_0.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_0.CD ) ,
    .IN ( masks_shift_reg_10_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_2.DI_ ) ,
    .IN ( n82 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_2.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_2 ) ,
    .IN ( masks_hold_reg_4_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_2.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_2.QT ) ,
    .I1 ( masks_hold_reg_4_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_2.ED ) ,
    .S ( masks_hold_reg_4_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_2.ED ) ,
    .I1 ( masks_hold_reg_4_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_2.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_10_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_3.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_3.CD ) ,
    .IN ( masks_shift_reg_10_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_1.DI_ ) ,
    .IN ( n81 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_1.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_1 ) ,
    .IN ( masks_hold_reg_4_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_1.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_1.QT ) ,
    .I1 ( masks_hold_reg_4_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_1.ED ) ,
    .S ( masks_hold_reg_4_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_1.ED ) ,
    .I1 ( masks_hold_reg_4_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_1.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_10_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_2.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_2.CD ) ,
    .IN ( masks_shift_reg_10_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_4_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_0.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_0 ) ,
    .IN ( masks_hold_reg_4_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_0.QT ) ,
    .I1 ( masks_hold_reg_4_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_0.ED ) ,
    .S ( masks_hold_reg_4_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_0.ED ) ,
    .I1 ( masks_hold_reg_4_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_0.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_10_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_5.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_5.CD ) ,
    .IN ( masks_shift_reg_10_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_7.DI_ ) ,
    .IN ( n89 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_7.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_7 ) ,
    .IN ( masks_hold_reg_4_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_7.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_7.QT ) ,
    .I1 ( masks_hold_reg_4_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_7.ED ) ,
    .S ( masks_hold_reg_4_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_7.ED ) ,
    .I1 ( masks_hold_reg_4_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_10_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_4.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_4.CD ) ,
    .IN ( masks_shift_reg_10_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_6.DI_ ) ,
    .IN ( n88 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_6.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_6 ) ,
    .IN ( masks_hold_reg_4_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_6.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_6.QT ) ,
    .I1 ( masks_hold_reg_4_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_6.ED ) ,
    .S ( masks_hold_reg_4_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_6.ED ) ,
    .I1 ( masks_hold_reg_4_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_10_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_7.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_7.CD ) ,
    .IN ( masks_shift_reg_10_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_5.DI_ ) ,
    .IN ( n80 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_5.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_5 ) ,
    .IN ( masks_hold_reg_4_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_5.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_5.QT ) ,
    .I1 ( masks_hold_reg_4_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_5.ED ) ,
    .S ( masks_hold_reg_4_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_5.ED ) ,
    .I1 ( masks_hold_reg_4_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_5.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_10_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_10_reg_6.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_6.CD ) ,
    .IN ( masks_shift_reg_10_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_10_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_10_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_10_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_10_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_10_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_10_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_10_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_10_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_10_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_10_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_10_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_10_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_4.DI_ ) ,
    .IN ( n35 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_4.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_4 ) ,
    .IN ( masks_hold_reg_4_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_4_reg_4.QT ) ,
    .I1 ( masks_hold_reg_4_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_4.ED ) ,
    .S ( masks_hold_reg_4_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_4.ED ) ,
    .I1 ( masks_hold_reg_4_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_4_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_4_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_4.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_6_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_8.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_8.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_8.CD ) ,
    .IN ( masks_shift_reg_6_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_9.DI_ ) ,
    .IN ( n94 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_9.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_9 ) ,
    .IN ( masks_hold_reg_4_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_9.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_9.QT ) ,
    .I1 ( masks_hold_reg_4_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_9.ED ) ,
    .S ( masks_hold_reg_4_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_9.ED ) ,
    .I1 ( masks_hold_reg_4_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_9.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_6_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_9.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_9.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_9.CD ) ,
    .IN ( masks_shift_reg_6_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_4_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_8.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_8 ) ,
    .IN ( masks_hold_reg_4_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_8.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_4_reg_8.QT ) ,
    .I1 ( masks_hold_reg_4_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_8.ED ) ,
    .S ( masks_hold_reg_4_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_8.ED ) ,
    .I1 ( masks_hold_reg_4_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_4_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_4_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_6_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_6.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_6.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_6.CD ) ,
    .IN ( masks_shift_reg_6_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_6_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_7.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_7.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29287 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_7.CD ) ,
    .IN ( masks_shift_reg_6_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_6_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_4.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_4.CD ) ,
    .IN ( masks_shift_reg_6_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_5.DI_ ) ,
    .IN ( n95 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_5.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_5.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_5.CD ) ,
    .IN ( masks_shift_reg_6_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_6_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_2.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_2.CD ) ,
    .IN ( masks_shift_reg_6_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_1_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_9.CPI_ ) ,
    .IN ( edt_clock ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_9.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_9.CD ) ,
    .IN ( masks_shift_reg_1_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_6_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_3.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_3.CD ) ,
    .IN ( masks_shift_reg_6_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_1_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_8.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_8.CD ) ,
    .IN ( masks_shift_reg_1_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_6_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_0.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_0.CD ) ,
    .IN ( masks_shift_reg_6_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_6_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_6_reg_1.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_1.CD ) ,
    .IN ( masks_shift_reg_6_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_6_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_6_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_6_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_6_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_6_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_6_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_6_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_6_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_6_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_6_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_6_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_6_1 ) ) ;
and ( 
    .Z ( U984.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_100 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U984.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_47 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U984.EF ) ,
    .I0 ( xor_decoded_masks_8_47 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_47 ) ,
    .I0 ( U984.AB ) ,
    .I1 ( U984.CD ) ,
    .I2 ( U984.EF ) ) ;
and ( 
    .Z ( U689.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_91 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U689.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_38 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U689.EF ) ,
    .I0 ( xor_decoded_masks_12_38 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_38 ) ,
    .I0 ( U689.AB ) ,
    .I1 ( U689.CD ) ,
    .I2 ( U689.EF ) ) ;
and ( 
    .Z ( U985.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_100 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U985.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_47 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U985.EF ) ,
    .I0 ( xor_decoded_masks_10_47 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_47 ) ,
    .I0 ( U985.AB ) ,
    .I1 ( U985.CD ) ,
    .I2 ( U985.EF ) ) ;
and ( 
    .Z ( U688.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_87 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U688.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_34 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U688.EF ) ,
    .I0 ( xor_decoded_masks_12_34 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_34 ) ,
    .I0 ( U688.AB ) ,
    .I1 ( U688.CD ) ,
    .I2 ( U688.EF ) ) ;
and ( 
    .Z ( U986.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_9 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U986.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_9 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U986.EF ) ,
    .I0 ( xor_decoded_masks_0_9 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_9 ) ,
    .I0 ( U986.AB ) ,
    .I1 ( U986.CD ) ,
    .I2 ( U986.EF ) ) ;
and ( 
    .Z ( U987.AB ) ,
    .I0 ( masks_hold_reg_12_6 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U987.CD ) ,
    .I0 ( config1_xor_encoded_masks_135 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_135 ) ,
    .I0 ( U987.AB ) ,
    .I1 ( U987.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_1_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_1.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_1.CD ) ,
    .IN ( masks_shift_reg_1_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_1 ) ) ;
and ( 
    .Z ( U980.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_154 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U980.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_47 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U980.EF ) ,
    .I0 ( xor_decoded_masks_2_47 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_47 ) ,
    .I0 ( U980.AB ) ,
    .I1 ( U980.CD ) ,
    .I2 ( U980.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_1_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_0.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_0.CD ) ,
    .IN ( masks_shift_reg_1_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_0 ) ) ;
and ( 
    .Z ( U981.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_47 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U981.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_47 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U981.EF ) ,
    .I0 ( xor_decoded_masks_3_47 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_47 ) ,
    .I0 ( U981.AB ) ,
    .I1 ( U981.CD ) ,
    .I2 ( U981.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_1_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_3.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_3.CD ) ,
    .IN ( masks_shift_reg_1_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_3 ) ) ;
and ( 
    .Z ( U982.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_100 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U982.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_47 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U982.EF ) ,
    .I0 ( xor_decoded_masks_6_47 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_47 ) ,
    .I0 ( U982.AB ) ,
    .I1 ( U982.CD ) ,
    .I2 ( U982.EF ) ) ;
and ( 
    .Z ( U683.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_91 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U683.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_38 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U683.EF ) ,
    .I0 ( xor_decoded_masks_8_38 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_38 ) ,
    .I0 ( U683.AB ) ,
    .I1 ( U683.CD ) ,
    .I2 ( U683.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_1_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_1_reg_2.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_2.CD ) ,
    .IN ( masks_shift_reg_1_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_1_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_1_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_1_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_1_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_1_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_1_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_1_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_1_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_1_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_1_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_1_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_1_2 ) ) ;
and ( 
    .Z ( U983.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_47 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U983.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_47 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U983.EF ) ,
    .I0 ( xor_decoded_masks_7_47 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_47 ) ,
    .I0 ( U983.AB ) ,
    .I1 ( U983.CD ) ,
    .I2 ( U983.EF ) ) ;
and ( 
    .Z ( U327.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_39 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U327.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_39 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U327.EF ) ,
    .I0 ( xor_decoded_masks_0_39 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_39 ) ,
    .I0 ( U327.AB ) ,
    .I1 ( U327.CD ) ,
    .I2 ( U327.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_6_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_6.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_6.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_6 ) ,
    .IN ( masks_hold_reg_6_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_6.QT ) ,
    .I1 ( masks_hold_reg_6_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_6.ED ) ,
    .S ( masks_hold_reg_6_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_6.ED ) ,
    .I1 ( masks_hold_reg_6_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_4_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_8.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_8.CD ) ,
    .IN ( masks_shift_reg_4_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_6_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_9.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_9.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_9 ) ,
    .IN ( masks_hold_reg_6_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_9.QT ) ,
    .I1 ( masks_hold_reg_6_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_9.ED ) ,
    .S ( masks_hold_reg_6_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_9.ED ) ,
    .I1 ( masks_hold_reg_6_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_9.QT ) ) ;
and ( 
    .Z ( U321.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_40 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U321.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_40 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U321.EF ) ,
    .I0 ( xor_decoded_masks_0_40 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_40 ) ,
    .I0 ( U321.AB ) ,
    .I1 ( U321.CD ) ,
    .I2 ( U321.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_4_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_9.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_9.CD ) ,
    .IN ( masks_shift_reg_4_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_6_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_8.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_8.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_8 ) ,
    .IN ( masks_hold_reg_6_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_8.QT ) ,
    .I1 ( masks_hold_reg_6_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_8.ED ) ,
    .S ( masks_hold_reg_6_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_8.ED ) ,
    .I1 ( masks_hold_reg_6_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_8.QT ) ) ;
and ( 
    .Z ( U322.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_42 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U322.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_42 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U322.EF ) ,
    .I0 ( xor_decoded_masks_0_42 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_42 ) ,
    .I0 ( U322.AB ) ,
    .I1 ( U322.CD ) ,
    .I2 ( U322.EF ) ) ;
and ( 
    .Z ( U323.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_43 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U323.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_43 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U323.EF ) ,
    .I0 ( xor_decoded_masks_0_43 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_43 ) ,
    .I0 ( U323.AB ) ,
    .I1 ( U323.CD ) ,
    .I2 ( U323.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_4_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_4.CD ) ,
    .IN ( masks_shift_reg_4_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_4_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_5.CD ) ,
    .IN ( masks_shift_reg_4_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_4_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_6.CD ) ,
    .IN ( masks_shift_reg_4_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_4_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_7.CD ) ,
    .IN ( masks_shift_reg_4_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_7 ) ) ;
nor ( 
    .Z ( n66 ) ,
    .I0 ( n26 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
and ( 
    .Z ( U328.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_36 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U328.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_36 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U328.EF ) ,
    .I0 ( xor_decoded_masks_0_36 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_36 ) ,
    .I0 ( U328.AB ) ,
    .I1 ( U328.CD ) ,
    .I2 ( U328.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_4_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_0.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_0.CD ) ,
    .IN ( masks_shift_reg_4_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_0 ) ) ;
and ( 
    .Z ( U329.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_38 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U329.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_38 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U329.EF ) ,
    .I0 ( xor_decoded_masks_0_38 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_38 ) ,
    .I0 ( U329.AB ) ,
    .I1 ( U329.CD ) ,
    .I2 ( U329.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_4_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_1.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_1.CD ) ,
    .IN ( masks_shift_reg_4_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_4_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_2.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_2.CD ) ,
    .IN ( masks_shift_reg_4_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_4_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2781 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_3.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_3.CD ) ,
    .IN ( masks_shift_reg_4_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_4_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_4_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_4_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_4_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_4_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_4_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_4_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_4_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_4_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_4_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_4_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_4_3 ) ) ;
nor ( 
    .Z ( n20 ) ,
    .I0 ( n40 ) ,
    .I1 ( edt_update_hfs_netlink_29281 ) ) ;
and ( 
    .Z ( U566.AB ) ,
    .I0 ( masks_hold_reg_8_8 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U566.CD ) ,
    .I0 ( config1_xor_encoded_masks_89 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_89 ) ,
    .I0 ( U566.AB ) ,
    .I1 ( U566.CD ) ) ;
and ( 
    .Z ( U567.AB ) ,
    .I0 ( masks_hold_reg_0_5 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U567.CD ) ,
    .I0 ( config1_xor_encoded_masks_4 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_4 ) ,
    .I0 ( U567.AB ) ,
    .I1 ( U567.CD ) ) ;
and ( 
    .Z ( U1235.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_66 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1235.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_13 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1235.EF ) ,
    .I0 ( xor_decoded_masks_14_13 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_13 ) ,
    .I0 ( U1235.AB ) ,
    .I1 ( U1235.CD ) ,
    .I2 ( U1235.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_5_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_2 ) ,
    .IN ( masks_hold_reg_5_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_2.QT ) ,
    .I1 ( masks_hold_reg_5_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_2.ED ) ,
    .S ( masks_hold_reg_5_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_2.ED ) ,
    .I1 ( masks_hold_reg_5_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_2.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_10_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_6 ) ,
    .IN ( masks_hold_reg_10_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_6.QT ) ,
    .I1 ( masks_hold_reg_10_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_6.ED ) ,
    .S ( masks_hold_reg_10_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_6.ED ) ,
    .I1 ( masks_hold_reg_10_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_10_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_7 ) ,
    .IN ( masks_hold_reg_10_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_7.QT ) ,
    .I1 ( masks_hold_reg_10_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_7.ED ) ,
    .S ( masks_hold_reg_10_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_7.ED ) ,
    .I1 ( masks_hold_reg_10_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_10_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_4 ) ,
    .IN ( masks_hold_reg_10_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_4.QT ) ,
    .I1 ( masks_hold_reg_10_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_4.ED ) ,
    .S ( masks_hold_reg_10_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_4.ED ) ,
    .I1 ( masks_hold_reg_10_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_4.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_10_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_5 ) ,
    .IN ( masks_hold_reg_10_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_5.QT ) ,
    .I1 ( masks_hold_reg_10_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_5.ED ) ,
    .S ( masks_hold_reg_10_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_5.ED ) ,
    .I1 ( masks_hold_reg_10_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_5.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_10_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_2 ) ,
    .IN ( masks_hold_reg_10_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_2.QT ) ,
    .I1 ( masks_hold_reg_10_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_2.ED ) ,
    .S ( masks_hold_reg_10_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_2.ED ) ,
    .I1 ( masks_hold_reg_10_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_2.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_10_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_3 ) ,
    .IN ( masks_hold_reg_10_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_3.QT ) ,
    .I1 ( masks_hold_reg_10_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_3.ED ) ,
    .S ( masks_hold_reg_10_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_3.ED ) ,
    .I1 ( masks_hold_reg_10_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_10_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_0 ) ,
    .IN ( masks_hold_reg_10_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_10_reg_0.QT ) ,
    .I1 ( masks_hold_reg_10_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_0.ED ) ,
    .S ( masks_hold_reg_10_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_0.ED ) ,
    .I1 ( masks_hold_reg_10_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_10_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_10_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_0.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_10_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_1 ) ,
    .IN ( masks_hold_reg_10_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_1.QT ) ,
    .I1 ( masks_hold_reg_10_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_1.ED ) ,
    .S ( masks_hold_reg_10_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_1.ED ) ,
    .I1 ( masks_hold_reg_10_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_1.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_10_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_8.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_8 ) ,
    .IN ( masks_hold_reg_10_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_8.QT ) ,
    .I1 ( masks_hold_reg_10_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_8.ED ) ,
    .S ( masks_hold_reg_10_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_8.ED ) ,
    .I1 ( masks_hold_reg_10_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_10_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_9.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_9 ) ,
    .IN ( masks_hold_reg_10_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_9.QT ) ,
    .I1 ( masks_hold_reg_10_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_9.ED ) ,
    .S ( masks_hold_reg_10_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_9.ED ) ,
    .I1 ( masks_hold_reg_10_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_9.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_10.DI_ ) ,
    .IN ( edt_channels_out_from_constant_shift_control_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_2_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_10.CDNI_ ) ,
    .IN ( n54 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_10.CD ) ,
    .IN ( masks_shift_reg_0_reg_10.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_24 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_25 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_10.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_10.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_10.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_10.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_10.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_10.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_10.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_24 ) ,
    .Q ( masks_shift_reg_0_reg_10.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_25 ) ) ;
DFF masks_shift_reg_0_reg_10.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_10.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_10 ) ) ;
and ( 
    .Z ( U360.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_70 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U360.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_16 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U360.EF ) ,
    .I0 ( xor_decoded_masks_1_16 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_16 ) ,
    .I0 ( U360.AB ) ,
    .I1 ( U360.CD ) ,
    .I2 ( U360.EF ) ) ;
and ( 
    .Z ( U361.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_72 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U361.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_18 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U361.EF ) ,
    .I0 ( xor_decoded_masks_1_18 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_18 ) ,
    .I0 ( U361.AB ) ,
    .I1 ( U361.CD ) ,
    .I2 ( U361.EF ) ) ;
and ( 
    .Z ( U362.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_73 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U362.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_19 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U362.EF ) ,
    .I0 ( xor_decoded_masks_1_19 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_19 ) ,
    .I0 ( U362.AB ) ,
    .I1 ( U362.CD ) ,
    .I2 ( U362.EF ) ) ;
and ( 
    .Z ( U363.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_111 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U363.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_4 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U363.EF ) ,
    .I0 ( xor_decoded_masks_2_4 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_4 ) ,
    .I0 ( U363.AB ) ,
    .I1 ( U363.CD ) ,
    .I2 ( U363.EF ) ) ;
and ( 
    .Z ( U364.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_127 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U364.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_20 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U364.EF ) ,
    .I0 ( xor_decoded_masks_2_20 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_20 ) ,
    .I0 ( U364.AB ) ,
    .I1 ( U364.CD ) ,
    .I2 ( U364.EF ) ) ;
and ( 
    .Z ( U365.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_81 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U365.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_28 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U365.EF ) ,
    .I0 ( xor_decoded_masks_12_28 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_28 ) ,
    .I0 ( U365.AB ) ,
    .I1 ( U365.CD ) ,
    .I2 ( U365.EF ) ) ;
and ( 
    .Z ( U366.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_81 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U366.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_28 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U366.EF ) ,
    .I0 ( xor_decoded_masks_14_28 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_28 ) ,
    .I0 ( U366.AB ) ,
    .I1 ( U366.CD ) ,
    .I2 ( U366.EF ) ) ;
and ( 
    .Z ( U368.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_0 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U368.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_0 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U368.EF ) ,
    .I0 ( xor_decoded_masks_13_0 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_0 ) ,
    .I0 ( U368.AB ) ,
    .I1 ( U368.CD ) ,
    .I2 ( U368.EF ) ) ;
and ( 
    .Z ( U369.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_16 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U369.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_16 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U369.EF ) ,
    .I0 ( xor_decoded_masks_13_16 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_16 ) ,
    .I0 ( U369.AB ) ,
    .I1 ( U369.CD ) ,
    .I2 ( U369.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_0_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_7.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_7 ) ,
    .IN ( masks_hold_reg_0_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_7.QT ) ,
    .I1 ( masks_hold_reg_0_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_7.ED ) ,
    .S ( masks_hold_reg_0_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_7.ED ) ,
    .I1 ( masks_hold_reg_0_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_0_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_6.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_6 ) ,
    .IN ( masks_hold_reg_0_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_6.QT ) ,
    .I1 ( masks_hold_reg_0_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_6.ED ) ,
    .S ( masks_hold_reg_0_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_6.ED ) ,
    .I1 ( masks_hold_reg_0_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_0_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_5.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_5 ) ,
    .IN ( masks_hold_reg_0_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_5.QT ) ,
    .I1 ( masks_hold_reg_0_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_5.ED ) ,
    .S ( masks_hold_reg_0_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_5.ED ) ,
    .I1 ( masks_hold_reg_0_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_5.QT ) ) ;
and ( 
    .Z ( U371.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_31 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U371.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_31 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U371.EF ) ,
    .I0 ( xor_decoded_masks_11_31 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_31 ) ,
    .I0 ( U371.AB ) ,
    .I1 ( U371.CD ) ,
    .I2 ( U371.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_0_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_4.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_4 ) ,
    .IN ( masks_hold_reg_0_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_4.QT ) ,
    .I1 ( masks_hold_reg_0_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_4.ED ) ,
    .S ( masks_hold_reg_0_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_4.ED ) ,
    .I1 ( masks_hold_reg_0_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_4.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_0_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_3.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_3 ) ,
    .IN ( masks_hold_reg_0_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_3.QT ) ,
    .I1 ( masks_hold_reg_0_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_3.ED ) ,
    .S ( masks_hold_reg_0_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_3.ED ) ,
    .I1 ( masks_hold_reg_0_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_3.QT ) ) ;
and ( 
    .Z ( U373.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_34 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U373.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_34 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U373.EF ) ,
    .I0 ( xor_decoded_masks_3_34 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_34 ) ,
    .I0 ( U373.AB ) ,
    .I1 ( U373.CD ) ,
    .I2 ( U373.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_0_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_2.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_2 ) ,
    .IN ( masks_hold_reg_0_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_2.QT ) ,
    .I1 ( masks_hold_reg_0_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_2.ED ) ,
    .S ( masks_hold_reg_0_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_2.ED ) ,
    .I1 ( masks_hold_reg_0_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_2.QT ) ) ;
and ( 
    .Z ( U372.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_48 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U372.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_48 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U372.EF ) ,
    .I0 ( xor_decoded_masks_11_48 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_48 ) ,
    .I0 ( U372.AB ) ,
    .I1 ( U372.CD ) ,
    .I2 ( U372.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_0_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_1.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_1 ) ,
    .IN ( masks_hold_reg_0_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_1.QT ) ,
    .I1 ( masks_hold_reg_0_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_1.ED ) ,
    .S ( masks_hold_reg_0_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_1.ED ) ,
    .I1 ( masks_hold_reg_0_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_1.QT ) ) ;
and ( 
    .Z ( U375.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_35 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U375.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_35 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U375.EF ) ,
    .I0 ( xor_decoded_masks_3_35 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_35 ) ,
    .I0 ( U375.AB ) ,
    .I1 ( U375.CD ) ,
    .I2 ( U375.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_0_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_0.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_0 ) ,
    .IN ( masks_hold_reg_0_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_0.QT ) ,
    .I1 ( masks_hold_reg_0_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_0.ED ) ,
    .S ( masks_hold_reg_0_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_0.ED ) ,
    .I1 ( masks_hold_reg_0_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_0.QT ) ) ;
and ( 
    .Z ( U374.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_33 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U374.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_33 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U374.EF ) ,
    .I0 ( xor_decoded_masks_3_33 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_33 ) ,
    .I0 ( U374.AB ) ,
    .I1 ( U374.CD ) ,
    .I2 ( U374.EF ) ) ;
and ( 
    .Z ( U377.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_23 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U377.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_23 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U377.EF ) ,
    .I0 ( xor_decoded_masks_3_23 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_23 ) ,
    .I0 ( U377.AB ) ,
    .I1 ( U377.CD ) ,
    .I2 ( U377.EF ) ) ;
and ( 
    .Z ( U376.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_22 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U376.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_22 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U376.EF ) ,
    .I0 ( xor_decoded_masks_3_22 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_22 ) ,
    .I0 ( U376.AB ) ,
    .I1 ( U376.CD ) ,
    .I2 ( U376.EF ) ) ;
and ( 
    .Z ( U379.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_28 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U379.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_28 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U379.EF ) ,
    .I0 ( xor_decoded_masks_5_28 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_28 ) ,
    .I0 ( U379.AB ) ,
    .I1 ( U379.CD ) ,
    .I2 ( U379.EF ) ) ;
and ( 
    .Z ( U378.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_76 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U378.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_23 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U378.EF ) ,
    .I0 ( xor_decoded_masks_4_23 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_23 ) ,
    .I0 ( U378.AB ) ,
    .I1 ( U378.CD ) ,
    .I2 ( U378.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_13_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_5 ) ,
    .IN ( masks_hold_reg_13_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_5.QT ) ,
    .I1 ( masks_hold_reg_13_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_5.ED ) ,
    .S ( masks_hold_reg_13_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_5.ED ) ,
    .I1 ( masks_hold_reg_13_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_5.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_0_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_9.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_9 ) ,
    .IN ( masks_hold_reg_0_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_9.QT ) ,
    .I1 ( masks_hold_reg_0_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_9.ED ) ,
    .S ( masks_hold_reg_0_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_9.ED ) ,
    .I1 ( masks_hold_reg_0_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_9.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_13_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_4 ) ,
    .IN ( masks_hold_reg_13_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_4.QT ) ,
    .I1 ( masks_hold_reg_13_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_4.ED ) ,
    .S ( masks_hold_reg_13_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_4.ED ) ,
    .I1 ( masks_hold_reg_13_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_4.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_0_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_8.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_8 ) ,
    .IN ( masks_hold_reg_0_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_0_reg_8.QT ) ,
    .I1 ( masks_hold_reg_0_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_8.ED ) ,
    .S ( masks_hold_reg_0_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_8.ED ) ,
    .I1 ( masks_hold_reg_0_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_0_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_0_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_13_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_7 ) ,
    .IN ( masks_hold_reg_13_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_7.QT ) ,
    .I1 ( masks_hold_reg_13_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_7.ED ) ,
    .S ( masks_hold_reg_13_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_7.ED ) ,
    .I1 ( masks_hold_reg_13_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_13_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_6 ) ,
    .IN ( masks_hold_reg_13_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_6.QT ) ,
    .I1 ( masks_hold_reg_13_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_6.ED ) ,
    .S ( masks_hold_reg_13_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_6.ED ) ,
    .I1 ( masks_hold_reg_13_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_13_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_1 ) ,
    .IN ( masks_hold_reg_13_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_1.QT ) ,
    .I1 ( masks_hold_reg_13_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_1.ED ) ,
    .S ( masks_hold_reg_13_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_1.ED ) ,
    .I1 ( masks_hold_reg_13_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_1.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_13_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_0 ) ,
    .IN ( masks_hold_reg_13_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_0.QT ) ,
    .I1 ( masks_hold_reg_13_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_0.ED ) ,
    .S ( masks_hold_reg_13_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_0.ED ) ,
    .I1 ( masks_hold_reg_13_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_0.QT ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_10.DI_ ) ,
    .IN ( N157 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_5_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_5 ) ) ;
DFF masks_shift_reg_5_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_5_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_5_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_5_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_13_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_3 ) ,
    .IN ( masks_hold_reg_13_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_3.QT ) ,
    .I1 ( masks_hold_reg_13_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_3.ED ) ,
    .S ( masks_hold_reg_13_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_3.ED ) ,
    .I1 ( masks_hold_reg_13_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_13_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_13_2 ) ,
    .IN ( masks_hold_reg_13_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_13_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_13_reg_2.QT ) ,
    .I1 ( masks_hold_reg_13_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_13_reg_2.ED ) ,
    .S ( masks_hold_reg_13_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_13_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_13_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_13_reg_2.ED ) ,
    .I1 ( masks_hold_reg_13_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_13_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_13_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_13_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_13_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_13_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_13_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_13_reg_2.QT ) ) ;
and ( 
    .Z ( U342.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_81 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U342.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_28 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U342.EF ) ,
    .I0 ( xor_decoded_masks_6_28 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_28 ) ,
    .I0 ( U342.AB ) ,
    .I1 ( U342.CD ) ,
    .I2 ( U342.EF ) ) ;
and ( 
    .Z ( U882.AB ) ,
    .I0 ( masks_hold_reg_9_8 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U882.CD ) ,
    .I0 ( config1_xor_encoded_masks_100 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_100 ) ,
    .I0 ( U882.AB ) ,
    .I1 ( U882.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_4_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_reg_10.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_4_10 ) ,
    .IN ( masks_hold_reg_4_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_4_reg_10.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_4_reg_10.QT ) ,
    .I1 ( masks_hold_reg_4_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_4_reg_10.ED ) ,
    .S ( masks_hold_reg_4_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_4_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_4_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_4_reg_10.ED ) ,
    .I1 ( masks_hold_reg_4_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_4_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_4_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_4_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_4_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_4_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_4_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_4_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_4_reg_10.QT ) ) ;
and ( 
    .Z ( U889.AB ) ,
    .I0 ( masks_hold_reg_6_1 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U889.CD ) ,
    .I0 ( config1_xor_encoded_masks_74 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_74 ) ,
    .I0 ( U889.AB ) ,
    .I1 ( U889.CD ) ) ;
and ( 
    .Z ( U888.AB ) ,
    .I0 ( masks_hold_reg_5_10 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U888.CD ) ,
    .I0 ( config1_xor_encoded_masks_54 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_54 ) ,
    .I0 ( U888.AB ) ,
    .I1 ( U888.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_0_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_0_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( n3 ) ,
    .IN ( masks_hold_reg_0_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_27 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_28 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_29 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_0_reg_10.SYNTEST_VL_LSI_MUX21_26786.I0 ( 
    .I0 ( masks_hold_reg_0_reg_10.QT ) ,
    .I1 ( masks_hold_reg_0_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_0_reg_10.ED ) ,
    .S ( masks_hold_reg_0_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_0_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_29 ) ) ;
and ( 
    .Z ( masks_hold_reg_0_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_0_reg_10.ED ) ,
    .I1 ( masks_hold_reg_0_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_0_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_0_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_27 ) ,
    .Q ( masks_hold_reg_0_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_0_reg_10.SYNTEST_EXP_ADDED_NET_28 ) ) ;
DFF masks_hold_reg_0_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_0_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_0_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_0_reg_10.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_3_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_4.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_4 ) ,
    .IN ( masks_hold_reg_3_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_4.QT ) ,
    .I1 ( masks_hold_reg_3_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_4.ED ) ,
    .S ( masks_hold_reg_3_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_4.ED ) ,
    .I1 ( masks_hold_reg_3_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_4.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_3_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_5.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_5 ) ,
    .IN ( masks_hold_reg_3_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_5.QT ) ,
    .I1 ( masks_hold_reg_3_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_5.ED ) ,
    .S ( masks_hold_reg_3_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_5.ED ) ,
    .I1 ( masks_hold_reg_3_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_5.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_3_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_6.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_6 ) ,
    .IN ( masks_hold_reg_3_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_6.QT ) ,
    .I1 ( masks_hold_reg_3_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_6.ED ) ,
    .S ( masks_hold_reg_3_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_6.ED ) ,
    .I1 ( masks_hold_reg_3_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_6.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_3_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_7.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_7 ) ,
    .IN ( masks_hold_reg_3_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_7.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_3_reg_7.QT ) ,
    .I1 ( masks_hold_reg_3_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_7.ED ) ,
    .S ( masks_hold_reg_3_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_7.ED ) ,
    .I1 ( masks_hold_reg_3_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_3_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_3_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_7.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_3_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_0.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_0 ) ,
    .IN ( masks_hold_reg_3_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_3_reg_0.QT ) ,
    .I1 ( masks_hold_reg_3_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_0.ED ) ,
    .S ( masks_hold_reg_3_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_0.ED ) ,
    .I1 ( masks_hold_reg_3_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_3_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_3_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_0.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_3_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_1.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_1 ) ,
    .IN ( masks_hold_reg_3_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_1.QT ) ,
    .I1 ( masks_hold_reg_3_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_1.ED ) ,
    .S ( masks_hold_reg_3_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_1.ED ) ,
    .I1 ( masks_hold_reg_3_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_1.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_3_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_2.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_2 ) ,
    .IN ( masks_hold_reg_3_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_2.QT ) ,
    .I1 ( masks_hold_reg_3_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_2.ED ) ,
    .S ( masks_hold_reg_3_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_2.ED ) ,
    .I1 ( masks_hold_reg_3_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_2.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_3_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_3.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_3 ) ,
    .IN ( masks_hold_reg_3_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_3_reg_3.QT ) ,
    .I1 ( masks_hold_reg_3_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_3.ED ) ,
    .S ( masks_hold_reg_3_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_3.ED ) ,
    .I1 ( masks_hold_reg_3_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_3_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_3_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_9_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_8.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_8 ) ,
    .IN ( masks_hold_reg_9_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_8.QT ) ,
    .I1 ( masks_hold_reg_9_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_8.ED ) ,
    .S ( masks_hold_reg_9_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_8.ED ) ,
    .I1 ( masks_hold_reg_9_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_8.DI_ ) ,
    .IN ( n87 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_8.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_8 ) ,
    .IN ( masks_hold_reg_3_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_8.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_3_reg_8.QT ) ,
    .I1 ( masks_hold_reg_3_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_8.ED ) ,
    .S ( masks_hold_reg_3_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_8.ED ) ,
    .I1 ( masks_hold_reg_3_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_3_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_3_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_9_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_9.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_9 ) ,
    .IN ( masks_hold_reg_9_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_9.QT ) ,
    .I1 ( masks_hold_reg_9_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_9.ED ) ,
    .S ( masks_hold_reg_9_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_9.ED ) ,
    .I1 ( masks_hold_reg_9_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_9.QT ) ) ;
and ( 
    .Z ( U894.AB ) ,
    .I0 ( masks_hold_reg_10_7 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U894.CD ) ,
    .I0 ( config1_xor_encoded_masks_112 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_112 ) ,
    .I0 ( U894.AB ) ,
    .I1 ( U894.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_3_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_reg_9.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_3_9 ) ,
    .IN ( masks_hold_reg_3_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_3_reg_9.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_3_reg_9.QT ) ,
    .I1 ( masks_hold_reg_3_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_3_reg_9.ED ) ,
    .S ( masks_hold_reg_3_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_3_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_3_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_3_reg_9.ED ) ,
    .I1 ( masks_hold_reg_3_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_3_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_3_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_3_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_3_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_3_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_3_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_3_reg_9.QT ) ) ;
and ( 
    .Z ( U478.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_60 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U478.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_7 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U478.EF ) ,
    .I0 ( xor_decoded_masks_14_7 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_7 ) ,
    .I0 ( U478.AB ) ,
    .I1 ( U478.CD ) ,
    .I2 ( U478.EF ) ) ;
and ( 
    .Z ( U564.AB ) ,
    .I0 ( masks_hold_reg_0_4 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U564.CD ) ,
    .I0 ( config1_xor_encoded_masks_5 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_5 ) ,
    .I0 ( U564.AB ) ,
    .I1 ( U564.CD ) ) ;
and ( 
    .Z ( U1234.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_62 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1234.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_9 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1234.EF ) ,
    .I0 ( xor_decoded_masks_14_9 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_9 ) ,
    .I0 ( U1234.AB ) ,
    .I1 ( U1234.CD ) ,
    .I2 ( U1234.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_5_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_3 ) ,
    .IN ( masks_hold_reg_5_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_3.QT ) ,
    .I1 ( masks_hold_reg_5_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_3.ED ) ,
    .S ( masks_hold_reg_5_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_3.ED ) ,
    .I1 ( masks_hold_reg_5_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_3.QT ) ) ;
and ( 
    .Z ( U565.AB ) ,
    .I0 ( n86 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U565.CD ) ,
    .I0 ( config1_xor_encoded_masks_25 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_25 ) ,
    .I0 ( U565.AB ) ,
    .I1 ( U565.CD ) ) ;
and ( 
    .Z ( U1237.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_150 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1237.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_43 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1237.EF ) ,
    .I0 ( xor_decoded_masks_2_43 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_43 ) ,
    .I0 ( U1237.AB ) ,
    .I1 ( U1237.CD ) ,
    .I2 ( U1237.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_9_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_reg_10.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_9_10 ) ,
    .IN ( masks_hold_reg_9_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_9_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_9_reg_10.QT ) ,
    .I1 ( masks_hold_reg_9_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_9_reg_10.ED ) ,
    .S ( masks_hold_reg_9_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_9_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_9_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_9_reg_10.ED ) ,
    .I1 ( masks_hold_reg_9_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_9_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_9_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_9_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_9_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_9_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_9_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_9_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_9_reg_10.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_5_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_0 ) ,
    .IN ( masks_hold_reg_5_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_0.QT ) ,
    .I1 ( masks_hold_reg_5_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_0.ED ) ,
    .S ( masks_hold_reg_5_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_0.ED ) ,
    .I1 ( masks_hold_reg_5_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_0.QT ) ) ;
and ( 
    .Z ( U1236.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_72 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1236.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_19 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1236.EF ) ,
    .I0 ( xor_decoded_masks_14_19 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_19 ) ,
    .I0 ( U1236.AB ) ,
    .I1 ( U1236.CD ) ,
    .I2 ( U1236.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_5_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_1 ) ,
    .IN ( masks_hold_reg_5_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_1.QT ) ,
    .I1 ( masks_hold_reg_5_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_1.ED ) ,
    .S ( masks_hold_reg_5_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_1.ED ) ,
    .I1 ( masks_hold_reg_5_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_1.QT ) ) ;
and ( 
    .Z ( U1231.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_23 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1231.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_23 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1231.EF ) ,
    .I0 ( xor_decoded_masks_13_23 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_23 ) ,
    .I0 ( U1231.AB ) ,
    .I1 ( U1231.CD ) ,
    .I2 ( U1231.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_5_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_6.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_6 ) ,
    .IN ( masks_hold_reg_5_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_6.QT ) ,
    .I1 ( masks_hold_reg_5_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_6.ED ) ,
    .S ( masks_hold_reg_5_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_6.ED ) ,
    .I1 ( masks_hold_reg_5_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_6.QT ) ) ;
and ( 
    .Z ( U1230.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_39 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1230.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_39 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1230.EF ) ,
    .I0 ( xor_decoded_masks_13_39 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_39 ) ,
    .I0 ( U1230.AB ) ,
    .I1 ( U1230.CD ) ,
    .I2 ( U1230.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_5_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_7.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_7 ) ,
    .IN ( masks_hold_reg_5_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_7.QT ) ,
    .I1 ( masks_hold_reg_5_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_7.ED ) ,
    .S ( masks_hold_reg_5_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_7.ED ) ,
    .I1 ( masks_hold_reg_5_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_7.QT ) ) ;
and ( 
    .Z ( U1233.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_13 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1233.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_13 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1233.EF ) ,
    .I0 ( xor_decoded_masks_13_13 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_13 ) ,
    .I0 ( U1233.AB ) ,
    .I1 ( U1233.CD ) ,
    .I2 ( U1233.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_5_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_4 ) ,
    .IN ( masks_hold_reg_5_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_4.QT ) ,
    .I1 ( masks_hold_reg_5_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_4.ED ) ,
    .S ( masks_hold_reg_5_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_4.ED ) ,
    .I1 ( masks_hold_reg_5_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_4.QT ) ) ;
and ( 
    .Z ( U1232.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_9 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1232.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_9 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1232.EF ) ,
    .I0 ( xor_decoded_masks_13_9 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_9 ) ,
    .I0 ( U1232.AB ) ,
    .I1 ( U1232.CD ) ,
    .I2 ( U1232.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_5_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_5.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_5 ) ,
    .IN ( masks_hold_reg_5_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_5.QT ) ,
    .I1 ( masks_hold_reg_5_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_5.ED ) ,
    .S ( masks_hold_reg_5_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_5.ED ) ,
    .I1 ( masks_hold_reg_5_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_5.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_5_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_8.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_8 ) ,
    .IN ( masks_hold_reg_5_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_5_reg_8.QT ) ,
    .I1 ( masks_hold_reg_5_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_8.ED ) ,
    .S ( masks_hold_reg_5_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_8.ED ) ,
    .I1 ( masks_hold_reg_5_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_5_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_5_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_5_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay1941 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_9.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_9 ) ,
    .IN ( masks_hold_reg_5_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_9.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_5_reg_9.QT ) ,
    .I1 ( masks_hold_reg_5_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_9.ED ) ,
    .S ( masks_hold_reg_5_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_9.ED ) ,
    .I1 ( masks_hold_reg_5_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_5_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_9.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_5_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_9.QT ) ) ;
and ( 
    .Z ( U1239.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_96 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1239.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_43 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1239.EF ) ,
    .I0 ( xor_decoded_masks_4_43 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_43 ) ,
    .I0 ( U1239.AB ) ,
    .I1 ( U1239.CD ) ,
    .I2 ( U1239.EF ) ) ;
and ( 
    .Z ( U568.AB ) ,
    .I0 ( masks_hold_reg_10_10 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U568.CD ) ,
    .I0 ( config1_xor_encoded_masks_109 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_109 ) ,
    .I0 ( U568.AB ) ,
    .I1 ( U568.CD ) ) ;
and ( 
    .Z ( U1238.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_43 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1238.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_43 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1238.EF ) ,
    .I0 ( xor_decoded_masks_3_43 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_43 ) ,
    .I0 ( U1238.AB ) ,
    .I1 ( U1238.CD ) ,
    .I2 ( U1238.EF ) ) ;
and ( 
    .Z ( U335.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_138 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U335.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_31 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U335.EF ) ,
    .I0 ( xor_decoded_masks_2_31 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_31 ) ,
    .I0 ( U335.AB ) ,
    .I1 ( U335.CD ) ,
    .I2 ( U335.EF ) ) ;
and ( 
    .Z ( U569.AB ) ,
    .I0 ( masks_hold_reg_2_5 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U569.CD ) ,
    .I0 ( config1_xor_encoded_masks_26 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_26 ) ,
    .I0 ( U569.AB ) ,
    .I1 ( U569.CD ) ) ;
and ( 
    .Z ( U334.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_137 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U334.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_30 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U334.EF ) ,
    .I0 ( xor_decoded_masks_2_30 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_30 ) ,
    .I0 ( U334.AB ) ,
    .I1 ( U334.CD ) ,
    .I2 ( U334.EF ) ) ;
and ( 
    .Z ( U337.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_130 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U337.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_23 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U337.EF ) ,
    .I0 ( xor_decoded_masks_2_23 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_23 ) ,
    .I0 ( U337.AB ) ,
    .I1 ( U337.CD ) ,
    .I2 ( U337.EF ) ) ;
and ( 
    .Z ( U336.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_129 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U336.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_22 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U336.EF ) ,
    .I0 ( xor_decoded_masks_2_22 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_22 ) ,
    .I0 ( U336.AB ) ,
    .I1 ( U336.CD ) ,
    .I2 ( U336.EF ) ) ;
and ( 
    .Z ( U331.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_32 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U331.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_32 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U331.EF ) ,
    .I0 ( xor_decoded_masks_0_32 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_32 ) ,
    .I0 ( U331.AB ) ,
    .I1 ( U331.CD ) ,
    .I2 ( U331.EF ) ) ;
and ( 
    .Z ( U330.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_33 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U330.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_33 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U330.EF ) ,
    .I0 ( xor_decoded_masks_0_33 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_33 ) ,
    .I0 ( U330.AB ) ,
    .I1 ( U330.CD ) ,
    .I2 ( U330.EF ) ) ;
and ( 
    .Z ( U333.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_135 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U333.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_28 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U333.EF ) ,
    .I0 ( xor_decoded_masks_2_28 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_28 ) ,
    .I0 ( U333.AB ) ,
    .I1 ( U333.CD ) ,
    .I2 ( U333.EF ) ) ;
and ( 
    .Z ( U332.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_34 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U332.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_34 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U332.EF ) ,
    .I0 ( xor_decoded_masks_0_34 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_34 ) ,
    .I0 ( U332.AB ) ,
    .I1 ( U332.CD ) ,
    .I2 ( U332.EF ) ) ;
and ( 
    .Z ( U339.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_84 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U339.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_31 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U339.EF ) ,
    .I0 ( xor_decoded_masks_4_31 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_31 ) ,
    .I0 ( U339.AB ) ,
    .I1 ( U339.CD ) ,
    .I2 ( U339.EF ) ) ;
and ( 
    .Z ( U338.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_81 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U338.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_28 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U338.EF ) ,
    .I0 ( xor_decoded_masks_4_28 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_28 ) ,
    .I0 ( U338.AB ) ,
    .I1 ( U338.CD ) ,
    .I2 ( U338.EF ) ) ;
and ( 
    .Z ( U577.AB ) ,
    .I0 ( masks_hold_reg_4_8 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U577.CD ) ,
    .I0 ( config1_xor_encoded_masks_45 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_45 ) ,
    .I0 ( U577.AB ) ,
    .I1 ( U577.CD ) ) ;
and ( 
    .Z ( U576.AB ) ,
    .I0 ( masks_hold_reg_2_8 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U576.CD ) ,
    .I0 ( config1_xor_encoded_masks_23 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_23 ) ,
    .I0 ( U576.AB ) ,
    .I1 ( U576.CD ) ) ;
and ( 
    .Z ( U1224.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_92 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1224.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_39 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1224.EF ) ,
    .I0 ( xor_decoded_masks_12_39 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_39 ) ,
    .I0 ( U1224.AB ) ,
    .I1 ( U1224.CD ) ,
    .I2 ( U1224.EF ) ) ;
and ( 
    .Z ( U575.AB ) ,
    .I0 ( masks_hold_reg_4_7 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U575.CD ) ,
    .I0 ( config1_xor_encoded_masks_46 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_46 ) ,
    .I0 ( U575.AB ) ,
    .I1 ( U575.CD ) ) ;
and ( 
    .Z ( U1225.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_62 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1225.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_9 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1225.EF ) ,
    .I0 ( xor_decoded_masks_12_9 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_9 ) ,
    .I0 ( U1225.AB ) ,
    .I1 ( U1225.CD ) ,
    .I2 ( U1225.EF ) ) ;
and ( 
    .Z ( U574.AB ) ,
    .I0 ( masks_hold_reg_6_10 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U574.CD ) ,
    .I0 ( config1_xor_encoded_masks_65 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_65 ) ,
    .I0 ( U574.AB ) ,
    .I1 ( U574.CD ) ) ;
and ( 
    .Z ( U1226.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_66 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1226.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_13 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1226.EF ) ,
    .I0 ( xor_decoded_masks_12_13 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_13 ) ,
    .I0 ( U1226.AB ) ,
    .I1 ( U1226.CD ) ,
    .I2 ( U1226.EF ) ) ;
and ( 
    .Z ( U573.AB ) ,
    .I0 ( masks_hold_reg_4_4 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U573.CD ) ,
    .I0 ( config1_xor_encoded_masks_49 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_49 ) ,
    .I0 ( U573.AB ) ,
    .I1 ( U573.CD ) ) ;
and ( 
    .Z ( U1227.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_72 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1227.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_19 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1227.EF ) ,
    .I0 ( xor_decoded_masks_12_19 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_19 ) ,
    .I0 ( U1227.AB ) ,
    .I1 ( U1227.CD ) ,
    .I2 ( U1227.EF ) ) ;
and ( 
    .Z ( U572.AB ) ,
    .I0 ( masks_hold_reg_2_2 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U572.CD ) ,
    .I0 ( config1_xor_encoded_masks_29 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_29 ) ,
    .I0 ( U572.AB ) ,
    .I1 ( U572.CD ) ) ;
and ( 
    .Z ( U1220.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_23 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1220.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_23 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1220.EF ) ,
    .I0 ( xor_decoded_masks_11_23 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_23 ) ,
    .I0 ( U1220.AB ) ,
    .I1 ( U1220.CD ) ,
    .I2 ( U1220.EF ) ) ;
and ( 
    .Z ( U571.AB ) ,
    .I0 ( masks_hold_reg_6_6 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U571.CD ) ,
    .I0 ( config1_xor_encoded_masks_69 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_69 ) ,
    .I0 ( U571.AB ) ,
    .I1 ( U571.CD ) ) ;
and ( 
    .Z ( U1221.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_9 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1221.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_9 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1221.EF ) ,
    .I0 ( xor_decoded_masks_11_9 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_9 ) ,
    .I0 ( U1221.AB ) ,
    .I1 ( U1221.CD ) ,
    .I2 ( U1221.EF ) ) ;
and ( 
    .Z ( U570.AB ) ,
    .I0 ( masks_hold_reg_8_9 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U570.CD ) ,
    .I0 ( config1_xor_encoded_masks_88 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_88 ) ,
    .I0 ( U570.AB ) ,
    .I1 ( U570.CD ) ) ;
and ( 
    .Z ( U1222.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_13 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1222.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_13 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1222.EF ) ,
    .I0 ( xor_decoded_masks_11_13 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_13 ) ,
    .I0 ( U1222.AB ) ,
    .I1 ( U1222.CD ) ,
    .I2 ( U1222.EF ) ) ;
and ( 
    .Z ( U1223.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_80 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1223.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_27 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1223.EF ) ,
    .I0 ( xor_decoded_masks_12_27 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_27 ) ,
    .I0 ( U1223.AB ) ,
    .I1 ( U1223.CD ) ,
    .I2 ( U1223.EF ) ) ;
and ( 
    .Z ( U1228.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_27 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1228.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_27 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1228.EF ) ,
    .I0 ( xor_decoded_masks_13_27 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_27 ) ,
    .I0 ( U1228.AB ) ,
    .I1 ( U1228.CD ) ,
    .I2 ( U1228.EF ) ) ;
and ( 
    .Z ( U579.AB ) ,
    .I0 ( masks_hold_reg_2_3 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U579.CD ) ,
    .I0 ( config1_xor_encoded_masks_28 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_28 ) ,
    .I0 ( U579.AB ) ,
    .I1 ( U579.CD ) ) ;
and ( 
    .Z ( U1229.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_35 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1229.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_35 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1229.EF ) ,
    .I0 ( xor_decoded_masks_13_35 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_35 ) ,
    .I0 ( U1229.AB ) ,
    .I1 ( U1229.CD ) ,
    .I2 ( U1229.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_10_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_10_10 ) ,
    .IN ( masks_hold_reg_10_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_10_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_10_reg_10.QT ) ,
    .I1 ( masks_hold_reg_10_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_10_reg_10.ED ) ,
    .S ( masks_hold_reg_10_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_10_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_10_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_10_reg_10.ED ) ,
    .I1 ( masks_hold_reg_10_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_10_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_10_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_10_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_10_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_10_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_10_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_10_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_10_reg_10.QT ) ) ;
and ( 
    .Z ( U578.AB ) ,
    .I0 ( masks_hold_reg_4_5 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U578.CD ) ,
    .I0 ( config1_xor_encoded_masks_48 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_48 ) ,
    .I0 ( U578.AB ) ,
    .I1 ( U578.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_13_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_2.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_2.CD ) ,
    .IN ( masks_shift_reg_13_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_13_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_3.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_3.CD ) ,
    .IN ( masks_shift_reg_13_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_13_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_0.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_0.CD ) ,
    .IN ( masks_shift_reg_13_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_13_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_1.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_1.CD ) ,
    .IN ( masks_shift_reg_13_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_13_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_6.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_6.CD ) ,
    .IN ( masks_shift_reg_13_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_7.DI_ ) ,
    .IN ( edt_channels_out_from_constant_shift_control_13 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_7.CDNI_ ) ,
    .IN ( n54 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_7.CD ) ,
    .IN ( masks_shift_reg_13_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_13_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_4.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_4.CD ) ,
    .IN ( masks_shift_reg_13_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_13_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_13_reg_5.CDNI_ ) ,
    .IN ( n53 ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_5.CD ) ,
    .IN ( masks_shift_reg_13_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_13_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_13_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_13_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_13_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_13_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_13_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_13_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_13_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_13_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_13_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_13_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_13_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_13_5 ) ) ;
and ( 
    .Z ( U343.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_84 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U343.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_31 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U343.EF ) ,
    .I0 ( xor_decoded_masks_6_31 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_31 ) ,
    .I0 ( U343.AB ) ,
    .I1 ( U343.CD ) ,
    .I2 ( U343.EF ) ) ;
and ( 
    .Z ( U340.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_83 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U340.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_30 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U340.EF ) ,
    .I0 ( xor_decoded_masks_4_30 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_30 ) ,
    .I0 ( U340.AB ) ,
    .I1 ( U340.CD ) ,
    .I2 ( U340.EF ) ) ;
and ( 
    .Z ( U341.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_75 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U341.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_22 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U341.EF ) ,
    .I0 ( xor_decoded_masks_4_22 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_22 ) ,
    .I0 ( U341.AB ) ,
    .I1 ( U341.CD ) ,
    .I2 ( U341.EF ) ) ;
and ( 
    .Z ( U346.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_76 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U346.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_23 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U346.EF ) ,
    .I0 ( xor_decoded_masks_6_23 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_23 ) ,
    .I0 ( U346.AB ) ,
    .I1 ( U346.CD ) ,
    .I2 ( U346.EF ) ) ;
and ( 
    .Z ( U347.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_81 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U347.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_28 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U347.EF ) ,
    .I0 ( xor_decoded_masks_8_28 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_28 ) ,
    .I0 ( U347.AB ) ,
    .I1 ( U347.CD ) ,
    .I2 ( U347.EF ) ) ;
and ( 
    .Z ( U344.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_83 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U344.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_30 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U344.EF ) ,
    .I0 ( xor_decoded_masks_6_30 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_30 ) ,
    .I0 ( U344.AB ) ,
    .I1 ( U344.CD ) ,
    .I2 ( U344.EF ) ) ;
and ( 
    .Z ( U345.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_75 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U345.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_22 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U345.EF ) ,
    .I0 ( xor_decoded_masks_6_22 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_22 ) ,
    .I0 ( U345.AB ) ,
    .I1 ( U345.CD ) ,
    .I2 ( U345.EF ) ) ;
and ( 
    .Z ( U348.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_84 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U348.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_31 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U348.EF ) ,
    .I0 ( xor_decoded_masks_8_31 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_31 ) ,
    .I0 ( U348.AB ) ,
    .I1 ( U348.CD ) ,
    .I2 ( U348.EF ) ) ;
and ( 
    .Z ( U349.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_83 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U349.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_30 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U349.EF ) ,
    .I0 ( xor_decoded_masks_8_30 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_30 ) ,
    .I0 ( U349.AB ) ,
    .I1 ( U349.CD ) ,
    .I2 ( U349.EF ) ) ;
and ( 
    .Z ( U353.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_83 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U353.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_30 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U353.EF ) ,
    .I0 ( xor_decoded_masks_10_30 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_30 ) ,
    .I0 ( U353.AB ) ,
    .I1 ( U353.CD ) ,
    .I2 ( U353.EF ) ) ;
and ( 
    .Z ( U352.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_84 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U352.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_31 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U352.EF ) ,
    .I0 ( xor_decoded_masks_10_31 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_31 ) ,
    .I0 ( U352.AB ) ,
    .I1 ( U352.CD ) ,
    .I2 ( U352.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_10.DI_ ) ,
    .IN ( N146 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_4_reg_10.CPI_ ) ,
    .IN ( edt_clock ) ) ;
DFF masks_shift_reg_4_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_4_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_4_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_4_10 ) ) ;
and ( 
    .Z ( U351.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_81 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U351.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_28 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U351.EF ) ,
    .I0 ( xor_decoded_masks_10_28 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_28 ) ,
    .I0 ( U351.AB ) ,
    .I1 ( U351.CD ) ,
    .I2 ( U351.EF ) ) ;
and ( 
    .Z ( U350.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_75 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U350.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_22 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U350.EF ) ,
    .I0 ( xor_decoded_masks_8_22 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_22 ) ,
    .I0 ( U350.AB ) ,
    .I1 ( U350.CD ) ,
    .I2 ( U350.EF ) ) ;
and ( 
    .Z ( U357.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_82 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U357.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_28 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U357.EF ) ,
    .I0 ( xor_decoded_masks_1_28 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_28 ) ,
    .I0 ( U357.AB ) ,
    .I1 ( U357.CD ) ,
    .I2 ( U357.EF ) ) ;
and ( 
    .Z ( U356.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_83 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U356.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_30 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U356.EF ) ,
    .I0 ( xor_decoded_masks_14_30 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_30 ) ,
    .I0 ( U356.AB ) ,
    .I1 ( U356.CD ) ,
    .I2 ( U356.EF ) ) ;
and ( 
    .Z ( U355.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_84 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U355.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_31 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U355.EF ) ,
    .I0 ( xor_decoded_masks_14_31 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_31 ) ,
    .I0 ( U355.AB ) ,
    .I1 ( U355.CD ) ,
    .I2 ( U355.EF ) ) ;
and ( 
    .Z ( U354.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_84 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U354.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_31 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U354.EF ) ,
    .I0 ( xor_decoded_masks_12_31 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_31 ) ,
    .I0 ( U354.AB ) ,
    .I1 ( U354.CD ) ,
    .I2 ( U354.EF ) ) ;
and ( 
    .Z ( U359.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_85 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U359.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_31 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U359.EF ) ,
    .I0 ( xor_decoded_masks_1_31 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_31 ) ,
    .I0 ( U359.AB ) ,
    .I1 ( U359.CD ) ,
    .I2 ( U359.EF ) ) ;
and ( 
    .Z ( U358.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_84 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U358.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_30 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U358.EF ) ,
    .I0 ( xor_decoded_masks_1_30 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_30 ) ,
    .I0 ( U358.AB ) ,
    .I1 ( U358.CD ) ,
    .I2 ( U358.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_6_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_1.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_1 ) ,
    .IN ( masks_hold_reg_6_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_1.QT ) ,
    .I1 ( masks_hold_reg_6_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_1.ED ) ,
    .S ( masks_hold_reg_6_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_1.ED ) ,
    .I1 ( masks_hold_reg_6_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_1.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_6_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_0.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_0.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_0 ) ,
    .IN ( masks_hold_reg_6_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_0.QT ) ,
    .I1 ( masks_hold_reg_6_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_0.ED ) ,
    .S ( masks_hold_reg_6_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_0.ED ) ,
    .I1 ( masks_hold_reg_6_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_0.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_6_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_3.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_3 ) ,
    .IN ( masks_hold_reg_6_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_3.QT ) ,
    .I1 ( masks_hold_reg_6_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_3.ED ) ,
    .S ( masks_hold_reg_6_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_3.ED ) ,
    .I1 ( masks_hold_reg_6_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_6_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_2.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_2 ) ,
    .IN ( masks_hold_reg_6_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_2.QT ) ,
    .I1 ( masks_hold_reg_6_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_2.ED ) ,
    .S ( masks_hold_reg_6_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_2.ED ) ,
    .I1 ( masks_hold_reg_6_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_2.QT ) ) ;
and ( 
    .Z ( U324.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_44 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U324.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_44 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U324.EF ) ,
    .I0 ( xor_decoded_masks_0_44 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_44 ) ,
    .I0 ( U324.AB ) ,
    .I1 ( U324.CD ) ,
    .I2 ( U324.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_6_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_5.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_5 ) ,
    .IN ( masks_hold_reg_6_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_5.QT ) ,
    .I1 ( masks_hold_reg_6_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_5.ED ) ,
    .S ( masks_hold_reg_6_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_5.ED ) ,
    .I1 ( masks_hold_reg_6_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_5.QT ) ) ;
and ( 
    .Z ( U325.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_46 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U325.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_46 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U325.EF ) ,
    .I0 ( xor_decoded_masks_0_46 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_46 ) ,
    .I0 ( U325.AB ) ,
    .I1 ( U325.CD ) ,
    .I2 ( U325.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_6_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_4.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_4 ) ,
    .IN ( masks_hold_reg_6_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_4.QT ) ,
    .I1 ( masks_hold_reg_6_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_4.ED ) ,
    .S ( masks_hold_reg_6_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_4.ED ) ,
    .I1 ( masks_hold_reg_6_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_4.QT ) ) ;
and ( 
    .Z ( U326.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_47 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U326.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_47 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U326.EF ) ,
    .I0 ( xor_decoded_masks_0_47 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_47 ) ,
    .I0 ( U326.AB ) ,
    .I1 ( U326.CD ) ,
    .I2 ( U326.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_6_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_7.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_7 ) ,
    .IN ( masks_hold_reg_6_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_6_reg_7.QT ) ,
    .I1 ( masks_hold_reg_6_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_7.ED ) ,
    .S ( masks_hold_reg_6_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_7.ED ) ,
    .I1 ( masks_hold_reg_6_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_6_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_6_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_7.QT ) ) ;
and ( 
    .Z ( U1037.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_40 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1037.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_40 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1037.EF ) ,
    .I0 ( xor_decoded_masks_5_40 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_40 ) ,
    .I0 ( U1037.AB ) ,
    .I1 ( U1037.CD ) ,
    .I2 ( U1037.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_11_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_0.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_0.CD ) ,
    .IN ( masks_shift_reg_11_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_0 ) ) ;
and ( 
    .Z ( U766.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_66 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U766.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_13 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U766.EF ) ,
    .I0 ( xor_decoded_masks_4_13 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_13 ) ,
    .I0 ( U766.AB ) ,
    .I1 ( U766.CD ) ,
    .I2 ( U766.EF ) ) ;
and ( 
    .Z ( U1036.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_93 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1036.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_40 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1036.EF ) ,
    .I0 ( xor_decoded_masks_4_40 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_40 ) ,
    .I0 ( U1036.AB ) ,
    .I1 ( U1036.CD ) ,
    .I2 ( U1036.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_11_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_1.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_1.CD ) ,
    .IN ( masks_shift_reg_11_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_1 ) ) ;
and ( 
    .Z ( U767.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_88 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U767.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_35 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U767.EF ) ,
    .I0 ( xor_decoded_masks_6_35 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_35 ) ,
    .I0 ( U767.AB ) ,
    .I1 ( U767.CD ) ,
    .I2 ( U767.EF ) ) ;
and ( 
    .Z ( U1035.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_40 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1035.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_40 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1035.EF ) ,
    .I0 ( xor_decoded_masks_3_40 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_40 ) ,
    .I0 ( U1035.AB ) ,
    .I1 ( U1035.CD ) ,
    .I2 ( U1035.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_11_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_2.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_2.CD ) ,
    .IN ( masks_shift_reg_11_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_2 ) ) ;
and ( 
    .Z ( U449.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_55 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U449.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_2 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U449.EF ) ,
    .I0 ( xor_decoded_masks_8_2 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_2 ) ,
    .I0 ( U449.AB ) ,
    .I1 ( U449.CD ) ,
    .I2 ( U449.EF ) ) ;
and ( 
    .Z ( U760.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_116 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U760.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_9 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U760.EF ) ,
    .I0 ( xor_decoded_masks_2_9 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_9 ) ,
    .I0 ( U760.AB ) ,
    .I1 ( U760.CD ) ,
    .I2 ( U760.EF ) ) ;
and ( 
    .Z ( U1034.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_147 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1034.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_40 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1034.EF ) ,
    .I0 ( xor_decoded_masks_2_40 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_40 ) ,
    .I0 ( U1034.AB ) ,
    .I1 ( U1034.CD ) ,
    .I2 ( U1034.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_11_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_3.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_3.CD ) ,
    .IN ( masks_shift_reg_11_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_3 ) ) ;
and ( 
    .Z ( U448.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_56 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U448.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_3 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U448.EF ) ,
    .I0 ( xor_decoded_masks_8_3 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_3 ) ,
    .I0 ( U448.AB ) ,
    .I1 ( U448.CD ) ,
    .I2 ( U448.EF ) ) ;
and ( 
    .Z ( U761.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_120 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U761.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_13 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U761.EF ) ,
    .I0 ( xor_decoded_masks_2_13 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_13 ) ,
    .I0 ( U761.AB ) ,
    .I1 ( U761.CD ) ,
    .I2 ( U761.EF ) ) ;
and ( 
    .Z ( U1033.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_69 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1033.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_16 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1033.EF ) ,
    .I0 ( xor_decoded_masks_14_16 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_16 ) ,
    .I0 ( U1033.AB ) ,
    .I1 ( U1033.CD ) ,
    .I2 ( U1033.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_11_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_4.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_4.CD ) ,
    .IN ( masks_shift_reg_11_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_4 ) ) ;
and ( 
    .Z ( U762.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_88 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U762.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_35 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U762.EF ) ,
    .I0 ( xor_decoded_masks_4_35 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_35 ) ,
    .I0 ( U762.AB ) ,
    .I1 ( U762.CD ) ,
    .I2 ( U762.EF ) ) ;
and ( 
    .Z ( U1032.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_63 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1032.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_10 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1032.EF ) ,
    .I0 ( xor_decoded_masks_14_10 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_10 ) ,
    .I0 ( U1032.AB ) ,
    .I1 ( U1032.CD ) ,
    .I2 ( U1032.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_11_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_5.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_5.CD ) ,
    .IN ( masks_shift_reg_11_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_5 ) ) ;
and ( 
    .Z ( U763.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_80 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U763.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_27 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U763.EF ) ,
    .I0 ( xor_decoded_masks_4_27 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_27 ) ,
    .I0 ( U763.AB ) ,
    .I1 ( U763.CD ) ,
    .I2 ( U763.EF ) ) ;
and ( 
    .Z ( U1031.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_67 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1031.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_14 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1031.EF ) ,
    .I0 ( xor_decoded_masks_14_14 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_14 ) ,
    .I0 ( U1031.AB ) ,
    .I1 ( U1031.CD ) ,
    .I2 ( U1031.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_11_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_6.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_6.CD ) ,
    .IN ( masks_shift_reg_11_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_6 ) ) ;
and ( 
    .Z ( U1030.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_14 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1030.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_14 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1030.EF ) ,
    .I0 ( xor_decoded_masks_13_14 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_14 ) ,
    .I0 ( U1030.AB ) ,
    .I1 ( U1030.CD ) ,
    .I2 ( U1030.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_11_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_7.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_7.CD ) ,
    .IN ( masks_shift_reg_11_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_7 ) ) ;
and ( 
    .Z ( U768.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_80 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U768.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_27 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U768.EF ) ,
    .I0 ( xor_decoded_masks_6_27 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_27 ) ,
    .I0 ( U768.AB ) ,
    .I1 ( U768.CD ) ,
    .I2 ( U768.EF ) ) ;
and ( 
    .Z ( U769.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_92 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U769.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_39 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U769.EF ) ,
    .I0 ( xor_decoded_masks_6_39 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_39 ) ,
    .I0 ( U769.AB ) ,
    .I1 ( U769.CD ) ,
    .I2 ( U769.EF ) ) ;
and ( 
    .Z ( U533.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_73 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U533.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_20 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U533.EF ) ,
    .I0 ( xor_decoded_masks_12_20 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_20 ) ,
    .I0 ( U533.AB ) ,
    .I1 ( U533.CD ) ,
    .I2 ( U533.EF ) ) ;
and ( 
    .Z ( U1039.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_40 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1039.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_40 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1039.EF ) ,
    .I0 ( xor_decoded_masks_7_40 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_40 ) ,
    .I0 ( U1039.AB ) ,
    .I1 ( U1039.CD ) ,
    .I2 ( U1039.EF ) ) ;
and ( 
    .Z ( U532.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_73 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U532.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_20 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U532.EF ) ,
    .I0 ( xor_decoded_masks_10_20 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_20 ) ,
    .I0 ( U532.AB ) ,
    .I1 ( U532.CD ) ,
    .I2 ( U532.EF ) ) ;
and ( 
    .Z ( U1260.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_51 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1260.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_51 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1260.EF ) ,
    .I0 ( xor_decoded_masks_7_51 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_51 ) ,
    .I0 ( U1260.AB ) ,
    .I1 ( U1260.CD ) ,
    .I2 ( U1260.EF ) ) ;
and ( 
    .Z ( U1038.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_93 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1038.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_40 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1038.EF ) ,
    .I0 ( xor_decoded_masks_6_40 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_40 ) ,
    .I0 ( U1038.AB ) ,
    .I1 ( U1038.CD ) ,
    .I2 ( U1038.EF ) ) ;
and ( 
    .Z ( U531.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_73 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U531.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_20 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U531.EF ) ,
    .I0 ( xor_decoded_masks_8_20 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_20 ) ,
    .I0 ( U531.AB ) ,
    .I1 ( U531.CD ) ,
    .I2 ( U531.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_7_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_0_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_9.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_9.CD ) ,
    .IN ( masks_shift_reg_7_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_8.DI_ ) ,
    .IN ( n51 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_8.CDNI_ ) ,
    .IN ( masks_shift_reg_7_9 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_8.CD ) ,
    .IN ( masks_shift_reg_7_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_7_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_7.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_7.CD ) ,
    .IN ( masks_shift_reg_7_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_7_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_6.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_6.CD ) ,
    .IN ( masks_shift_reg_7_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_6 ) ) ;
and ( 
    .Z ( U1217.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_27 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1217.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_27 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1217.EF ) ,
    .I0 ( xor_decoded_masks_11_27 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_27 ) ,
    .I0 ( U1217.AB ) ,
    .I1 ( U1217.CD ) ,
    .I2 ( U1217.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_7_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_5.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_5.CD ) ,
    .IN ( masks_shift_reg_7_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_5 ) ) ;
and ( 
    .Z ( U1216.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_72 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1216.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_19 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1216.EF ) ,
    .I0 ( xor_decoded_masks_10_19 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_19 ) ,
    .I0 ( U1216.AB ) ,
    .I1 ( U1216.CD ) ,
    .I2 ( U1216.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_4.DI_ ) ,
    .IN ( n36 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_4.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_4.CD ) ,
    .IN ( masks_shift_reg_7_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_4 ) ) ;
and ( 
    .Z ( U1215.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_66 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1215.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_13 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1215.EF ) ,
    .I0 ( xor_decoded_masks_10_13 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_13 ) ,
    .I0 ( U1215.AB ) ,
    .I1 ( U1215.CD ) ,
    .I2 ( U1215.EF ) ) ;
and ( 
    .Z ( U540.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_3 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U540.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_3 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U540.EF ) ,
    .I0 ( xor_decoded_masks_7_3 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_3 ) ,
    .I0 ( U540.AB ) ,
    .I1 ( U540.CD ) ,
    .I2 ( U540.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_7_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_3.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_3.CD ) ,
    .IN ( masks_shift_reg_7_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_3 ) ) ;
and ( 
    .Z ( U1214.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_62 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1214.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_9 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1214.EF ) ,
    .I0 ( xor_decoded_masks_10_9 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_9 ) ,
    .I0 ( U1214.AB ) ,
    .I1 ( U1214.CD ) ,
    .I2 ( U1214.EF ) ) ;
and ( 
    .Z ( U541.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_60 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U541.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_7 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U541.EF ) ,
    .I0 ( xor_decoded_masks_12_7 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_7 ) ,
    .I0 ( U541.AB ) ,
    .I1 ( U541.CD ) ,
    .I2 ( U541.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_7_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_2.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_2.CD ) ,
    .IN ( masks_shift_reg_7_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_2 ) ) ;
and ( 
    .Z ( U1213.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_92 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1213.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_39 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1213.EF ) ,
    .I0 ( xor_decoded_masks_10_39 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_39 ) ,
    .I0 ( U1213.AB ) ,
    .I1 ( U1213.CD ) ,
    .I2 ( U1213.EF ) ) ;
and ( 
    .Z ( U542.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_101 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U542.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_48 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U542.EF ) ,
    .I0 ( xor_decoded_masks_12_48 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_48 ) ,
    .I0 ( U542.AB ) ,
    .I1 ( U542.CD ) ,
    .I2 ( U542.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_7_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_1.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_1.CD ) ,
    .IN ( masks_shift_reg_7_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_1 ) ) ;
and ( 
    .Z ( U1212.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_13 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1212.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_13 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1212.EF ) ,
    .I0 ( xor_decoded_masks_9_13 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_13 ) ,
    .I0 ( U1212.AB ) ,
    .I1 ( U1212.CD ) ,
    .I2 ( U1212.EF ) ) ;
and ( 
    .Z ( U543.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_49 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U543.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_49 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U543.EF ) ,
    .I0 ( xor_decoded_masks_3_49 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_49 ) ,
    .I0 ( U543.AB ) ,
    .I1 ( U543.CD ) ,
    .I2 ( U543.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_7_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2801 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_7_reg_0.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_0.CD ) ,
    .IN ( masks_shift_reg_7_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_7_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_7_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_7_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_7_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_7_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_7_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_7_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_7_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_7_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_7_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_7_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_7_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_7_0 ) ) ;
and ( 
    .Z ( U1211.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_9 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1211.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_9 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1211.EF ) ,
    .I0 ( xor_decoded_masks_9_9 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_9 ) ,
    .I0 ( U1211.AB ) ,
    .I1 ( U1211.CD ) ,
    .I2 ( U1211.EF ) ) ;
and ( 
    .Z ( U1210.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_23 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1210.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_23 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1210.EF ) ,
    .I0 ( xor_decoded_masks_9_23 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_23 ) ,
    .I0 ( U1210.AB ) ,
    .I1 ( U1210.CD ) ,
    .I2 ( U1210.EF ) ) ;
and ( 
    .Z ( U467.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_57 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U467.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_4 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U467.EF ) ,
    .I0 ( xor_decoded_masks_12_4 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_4 ) ,
    .I0 ( U467.AB ) ,
    .I1 ( U467.CD ) ,
    .I2 ( U467.EF ) ) ;
and ( 
    .Z ( U466.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_3 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U466.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_3 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U466.EF ) ,
    .I0 ( xor_decoded_masks_11_3 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_3 ) ,
    .I0 ( U466.AB ) ,
    .I1 ( U466.CD ) ,
    .I2 ( U466.EF ) ) ;
and ( 
    .Z ( U465.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_0 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U465.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_0 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U465.EF ) ,
    .I0 ( xor_decoded_masks_11_0 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_0 ) ,
    .I0 ( U465.AB ) ,
    .I1 ( U465.CD ) ,
    .I2 ( U465.EF ) ) ;
and ( 
    .Z ( U464.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_6 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U464.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_6 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U464.EF ) ,
    .I0 ( xor_decoded_masks_11_6 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_6 ) ,
    .I0 ( U464.AB ) ,
    .I1 ( U464.CD ) ,
    .I2 ( U464.EF ) ) ;
and ( 
    .Z ( U463.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_7 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U463.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_7 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U463.EF ) ,
    .I0 ( xor_decoded_masks_11_7 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_7 ) ,
    .I0 ( U463.AB ) ,
    .I1 ( U463.CD ) ,
    .I2 ( U463.EF ) ) ;
and ( 
    .Z ( U462.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_4 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U462.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_4 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U462.EF ) ,
    .I0 ( xor_decoded_masks_11_4 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_4 ) ,
    .I0 ( U462.AB ) ,
    .I1 ( U462.CD ) ,
    .I2 ( U462.EF ) ) ;
and ( 
    .Z ( U1219.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_39 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1219.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_39 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1219.EF ) ,
    .I0 ( xor_decoded_masks_11_39 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_39 ) ,
    .I0 ( U1219.AB ) ,
    .I1 ( U1219.CD ) ,
    .I2 ( U1219.EF ) ) ;
and ( 
    .Z ( U461.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_55 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U461.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_2 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U461.EF ) ,
    .I0 ( xor_decoded_masks_10_2 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_2 ) ,
    .I0 ( U461.AB ) ,
    .I1 ( U461.CD ) ,
    .I2 ( U461.EF ) ) ;
and ( 
    .Z ( U1218.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_35 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1218.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_35 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1218.EF ) ,
    .I0 ( xor_decoded_masks_11_35 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_35 ) ,
    .I0 ( U1218.AB ) ,
    .I1 ( U1218.CD ) ,
    .I2 ( U1218.EF ) ) ;
or ( 
    .Z ( U315.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_3 ) ) ;
or ( 
    .Z ( U315.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_6 ) ) ;
and ( 
    .Z ( U315.ZN ) ,
    .I0 ( U315.AB ) ,
    .I1 ( U315.CD ) ) ;
not ( 
    .O1 ( N168 ) ,
    .IN ( U315.ZN ) ) ;
and ( 
    .Z ( U460.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_56 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U460.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_3 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U460.EF ) ,
    .I0 ( xor_decoded_masks_10_3 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_3 ) ,
    .I0 ( U460.AB ) ,
    .I1 ( U460.CD ) ,
    .I2 ( U460.EF ) ) ;
or ( 
    .Z ( U314.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_2 ) ) ;
or ( 
    .Z ( U314.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_4 ) ) ;
and ( 
    .Z ( U314.ZN ) ,
    .I0 ( U314.AB ) ,
    .I1 ( U314.CD ) ) ;
not ( 
    .O1 ( N146 ) ,
    .IN ( U314.ZN ) ) ;
or ( 
    .Z ( U313.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_1 ) ) ;
or ( 
    .Z ( U313.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_2 ) ) ;
and ( 
    .Z ( U313.ZN ) ,
    .I0 ( U313.AB ) ,
    .I1 ( U313.CD ) ) ;
not ( 
    .O1 ( N124 ) ,
    .IN ( U313.ZN ) ) ;
and ( 
    .Z ( U469.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_53 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U469.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_0 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U469.EF ) ,
    .I0 ( xor_decoded_masks_12_0 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_0 ) ,
    .I0 ( U469.AB ) ,
    .I1 ( U469.CD ) ,
    .I2 ( U469.EF ) ) ;
and ( 
    .Z ( U468.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_59 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U468.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_6 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U468.EF ) ,
    .I0 ( xor_decoded_masks_12_6 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_6 ) ,
    .I0 ( U468.AB ) ,
    .I1 ( U468.CD ) ,
    .I2 ( U468.EF ) ) ;
or ( 
    .Z ( U555.AB ) ,
    .I0 ( n11 ) ,
    .I1 ( n18 ) ) ;
or ( 
    .Z ( U555.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_5 ) ) ;
and ( 
    .Z ( U555.ZN ) ,
    .I0 ( U555.AB ) ,
    .I1 ( U555.CD ) ) ;
not ( 
    .O1 ( N157 ) ,
    .IN ( U555.ZN ) ) ;
or ( 
    .Z ( U554.AB ) ,
    .I0 ( n12 ) ,
    .I1 ( n18 ) ) ;
or ( 
    .Z ( U554.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_3 ) ) ;
and ( 
    .Z ( U554.ZN ) ,
    .I0 ( U554.AB ) ,
    .I1 ( U554.CD ) ) ;
not ( 
    .O1 ( N135 ) ,
    .IN ( U554.ZN ) ) ;
and ( 
    .Z ( U1206.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_72 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1206.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_19 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1206.EF ) ,
    .I0 ( xor_decoded_masks_8_19 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_19 ) ,
    .I0 ( U1206.AB ) ,
    .I1 ( U1206.CD ) ,
    .I2 ( U1206.EF ) ) ;
and ( 
    .Z ( U1207.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_27 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1207.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_27 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1207.EF ) ,
    .I0 ( xor_decoded_masks_9_27 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_27 ) ,
    .I0 ( U1207.AB ) ,
    .I1 ( U1207.CD ) ,
    .I2 ( U1207.EF ) ) ;
and ( 
    .Z ( U1204.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_9 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1204.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_9 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1204.EF ) ,
    .I0 ( xor_decoded_masks_7_9 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_9 ) ,
    .I0 ( U1204.AB ) ,
    .I1 ( U1204.CD ) ,
    .I2 ( U1204.EF ) ) ;
or ( 
    .Z ( U551.AB ) ,
    .I0 ( n41 ) ,
    .I1 ( n16 ) ) ;
and ( 
    .Z ( U551.ZN ) ,
    .I0 ( U551.AB ) ,
    .I1 ( n13 ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_0 ) ,
    .IN ( U551.ZN ) ) ;
and ( 
    .Z ( U1205.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_13 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1205.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_13 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1205.EF ) ,
    .I0 ( xor_decoded_masks_7_13 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_13 ) ,
    .I0 ( U1205.AB ) ,
    .I1 ( U1205.CD ) ,
    .I2 ( U1205.EF ) ) ;
not ( 
    .O1 ( n24 ) ,
    .IN ( n20 ) ) ;
and ( 
    .Z ( U1202.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_39 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1202.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_39 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1202.EF ) ,
    .I0 ( xor_decoded_masks_7_39 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_39 ) ,
    .I0 ( U1202.AB ) ,
    .I1 ( U1202.CD ) ,
    .I2 ( U1202.EF ) ) ;
or ( 
    .Z ( U553.AB ) ,
    .I0 ( n16 ) ,
    .I1 ( n18 ) ) ;
or ( 
    .Z ( U553.CD ) ,
    .I0 ( n24 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_1 ) ) ;
and ( 
    .Z ( U553.ZN ) ,
    .I0 ( U553.AB ) ,
    .I1 ( U553.CD ) ) ;
not ( 
    .O1 ( N113 ) ,
    .IN ( U553.ZN ) ) ;
and ( 
    .Z ( U1203.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_23 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1203.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_23 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1203.EF ) ,
    .I0 ( xor_decoded_masks_7_23 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_23 ) ,
    .I0 ( U1203.AB ) ,
    .I1 ( U1203.CD ) ,
    .I2 ( U1203.EF ) ) ;
or ( 
    .Z ( U552.AB ) ,
    .I0 ( n41 ) ,
    .I1 ( n12 ) ) ;
and ( 
    .Z ( U552.ZN ) ,
    .I0 ( U552.AB ) ,
    .I1 ( n13 ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_2 ) ,
    .IN ( U552.ZN ) ) ;
and ( 
    .Z ( U1200.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_27 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1200.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_27 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1200.EF ) ,
    .I0 ( xor_decoded_masks_7_27 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_27 ) ,
    .I0 ( U1200.AB ) ,
    .I1 ( U1200.CD ) ,
    .I2 ( U1200.EF ) ) ;
and ( 
    .Z ( U1201.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_35 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1201.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_35 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1201.EF ) ,
    .I0 ( xor_decoded_masks_7_35 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_35 ) ,
    .I0 ( U1201.AB ) ,
    .I1 ( U1201.CD ) ,
    .I2 ( U1201.EF ) ) ;
and ( 
    .Z ( U476.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_2 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U476.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_2 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U476.EF ) ,
    .I0 ( xor_decoded_masks_13_2 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_2 ) ,
    .I0 ( U476.AB ) ,
    .I1 ( U476.CD ) ,
    .I2 ( U476.EF ) ) ;
and ( 
    .Z ( U477.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_57 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U477.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_4 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U477.EF ) ,
    .I0 ( xor_decoded_masks_14_4 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_4 ) ,
    .I0 ( U477.AB ) ,
    .I1 ( U477.CD ) ,
    .I2 ( U477.EF ) ) ;
and ( 
    .Z ( U474.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_6 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U474.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_6 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U474.EF ) ,
    .I0 ( xor_decoded_masks_13_6 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_6 ) ,
    .I0 ( U474.AB ) ,
    .I1 ( U474.CD ) ,
    .I2 ( U474.EF ) ) ;
and ( 
    .Z ( U475.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_3 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U475.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_3 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U475.EF ) ,
    .I0 ( xor_decoded_masks_13_3 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_3 ) ,
    .I0 ( U475.AB ) ,
    .I1 ( U475.CD ) ,
    .I2 ( U475.EF ) ) ;
and ( 
    .Z ( U472.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_4 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U472.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_4 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U472.EF ) ,
    .I0 ( xor_decoded_masks_13_4 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_4 ) ,
    .I0 ( U472.AB ) ,
    .I1 ( U472.CD ) ,
    .I2 ( U472.EF ) ) ;
and ( 
    .Z ( U473.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_7 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U473.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_7 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U473.EF ) ,
    .I0 ( xor_decoded_masks_13_7 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_7 ) ,
    .I0 ( U473.AB ) ,
    .I1 ( U473.CD ) ,
    .I2 ( U473.EF ) ) ;
and ( 
    .Z ( U1208.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_35 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1208.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_35 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1208.EF ) ,
    .I0 ( xor_decoded_masks_9_35 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_35 ) ,
    .I0 ( U1208.AB ) ,
    .I1 ( U1208.CD ) ,
    .I2 ( U1208.EF ) ) ;
and ( 
    .Z ( U470.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_56 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U470.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_3 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U470.EF ) ,
    .I0 ( xor_decoded_masks_12_3 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_3 ) ,
    .I0 ( U470.AB ) ,
    .I1 ( U470.CD ) ,
    .I2 ( U470.EF ) ) ;
and ( 
    .Z ( U1209.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_39 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1209.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_39 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1209.EF ) ,
    .I0 ( xor_decoded_masks_9_39 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_39 ) ,
    .I0 ( U1209.AB ) ,
    .I1 ( U1209.CD ) ,
    .I2 ( U1209.EF ) ) ;
and ( 
    .Z ( U471.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_55 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U471.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_2 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U471.EF ) ,
    .I0 ( xor_decoded_masks_12_2 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_2 ) ,
    .I0 ( U471.AB ) ,
    .I1 ( U471.CD ) ,
    .I2 ( U471.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_0_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_2.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_2.CD ) ,
    .IN ( masks_shift_reg_0_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_2 ) ) ;
and ( 
    .Z ( U450.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_4 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U450.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_4 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U450.EF ) ,
    .I0 ( xor_decoded_masks_9_4 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_4 ) ,
    .I0 ( U450.AB ) ,
    .I1 ( U450.CD ) ,
    .I2 ( U450.EF ) ) ;
and ( 
    .Z ( U1304.AB ) ,
    .I0 ( edt_configuration_hfs_netlink_29291 ) ,
    .I1 ( masks_shift_reg_12_2 ) ) ;
and ( 
    .Z ( U1304.CD ) ,
    .I0 ( masks_shift_reg_13_0 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_13 ) ,
    .I0 ( U1304.AB ) ,
    .I1 ( U1304.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_0_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_3.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_3.CD ) ,
    .IN ( masks_shift_reg_0_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_3 ) ) ;
and ( 
    .Z ( U451.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_7 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U451.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_7 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U451.EF ) ,
    .I0 ( xor_decoded_masks_9_7 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_7 ) ,
    .I0 ( U451.AB ) ,
    .I1 ( U451.CD ) ,
    .I2 ( U451.EF ) ) ;
and ( 
    .Z ( U1303.AB ) ,
    .I0 ( edt_configuration_hfs_netlink_29290 ) ,
    .I1 ( masks_shift_reg_12_2 ) ) ;
and ( 
    .Z ( U1303.CD ) ,
    .I0 ( edt_channels_out_from_constant_shift_control_14 ) ,
    .I1 ( n45 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_14 ) ,
    .I0 ( U1303.AB ) ,
    .I1 ( U1303.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_0_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_4.CD ) ,
    .IN ( masks_shift_reg_0_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_4 ) ) ;
and ( 
    .Z ( U452.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_6 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U452.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_6 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U452.EF ) ,
    .I0 ( xor_decoded_masks_9_6 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_6 ) ,
    .I0 ( U452.AB ) ,
    .I1 ( U452.CD ) ,
    .I2 ( U452.EF ) ) ;
nand ( 
    .Z ( n13 ) ,
    .I0 ( masks_shift_reg_1_9 ) ,
    .I1 ( n37 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_0_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_5.CD ) ,
    .IN ( masks_shift_reg_0_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_5 ) ) ;
and ( 
    .Z ( U453.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_0 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U453.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_0 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U453.EF ) ,
    .I0 ( xor_decoded_masks_9_0 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_0 ) ,
    .I0 ( U453.AB ) ,
    .I1 ( U453.CD ) ,
    .I2 ( U453.EF ) ) ;
not ( 
    .O1 ( n8 ) ,
    .IN ( masks_shift_reg_5_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_0_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_6.CD ) ,
    .IN ( masks_shift_reg_0_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_6 ) ) ;
or ( 
    .Z ( U1300.AB ) ,
    .I0 ( n44 ) ,
    .I1 ( n8 ) ) ;
or ( 
    .Z ( U1300.CD ) ,
    .I0 ( n41 ) ,
    .I1 ( n9 ) ) ;
and ( 
    .Z ( U1300.ZN ) ,
    .I0 ( U1300.AB ) ,
    .I1 ( U1300.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_6 ) ,
    .IN ( U1300.ZN ) ) ;
and ( 
    .Z ( U775.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_92 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U775.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_39 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U775.EF ) ,
    .I0 ( xor_decoded_masks_8_39 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_39 ) ,
    .I0 ( U775.AB ) ,
    .I1 ( U775.CD ) ,
    .I2 ( U775.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_0_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_7.CD ) ,
    .IN ( masks_shift_reg_0_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_7 ) ) ;
and ( 
    .Z ( U774.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_80 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U774.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_27 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U774.EF ) ,
    .I0 ( xor_decoded_masks_8_27 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_27 ) ,
    .I0 ( U774.AB ) ,
    .I1 ( U774.CD ) ,
    .I2 ( U774.EF ) ) ;
and ( 
    .Z ( U1026.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_69 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1026.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_16 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1026.EF ) ,
    .I0 ( xor_decoded_masks_12_16 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_16 ) ,
    .I0 ( U1026.AB ) ,
    .I1 ( U1026.CD ) ,
    .I2 ( U1026.EF ) ) ;
and ( 
    .Z ( U777.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_66 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U777.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_13 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U777.EF ) ,
    .I0 ( xor_decoded_masks_8_13 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_13 ) ,
    .I0 ( U777.AB ) ,
    .I1 ( U777.CD ) ,
    .I2 ( U777.EF ) ) ;
and ( 
    .Z ( U1027.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_24 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1027.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_24 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1027.EF ) ,
    .I0 ( xor_decoded_masks_13_24 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_24 ) ,
    .I0 ( U1027.AB ) ,
    .I1 ( U1027.CD ) ,
    .I2 ( U1027.EF ) ) ;
and ( 
    .Z ( U776.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_62 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U776.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_9 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U776.EF ) ,
    .I0 ( xor_decoded_masks_8_9 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_9 ) ,
    .I0 ( U776.AB ) ,
    .I1 ( U776.CD ) ,
    .I2 ( U776.EF ) ) ;
and ( 
    .Z ( U1024.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_67 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1024.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_14 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1024.EF ) ,
    .I0 ( xor_decoded_masks_12_14 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_14 ) ,
    .I0 ( U1024.AB ) ,
    .I1 ( U1024.CD ) ,
    .I2 ( U1024.EF ) ) ;
and ( 
    .Z ( U458.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_59 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U458.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_6 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U458.EF ) ,
    .I0 ( xor_decoded_masks_10_6 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_6 ) ,
    .I0 ( U458.AB ) ,
    .I1 ( U458.CD ) ,
    .I2 ( U458.EF ) ) ;
and ( 
    .Z ( U771.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_66 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U771.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_13 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U771.EF ) ,
    .I0 ( xor_decoded_masks_6_13 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_13 ) ,
    .I0 ( U771.AB ) ,
    .I1 ( U771.CD ) ,
    .I2 ( U771.EF ) ) ;
and ( 
    .Z ( U1025.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_63 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1025.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_10 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1025.EF ) ,
    .I0 ( xor_decoded_masks_12_10 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_10 ) ,
    .I0 ( U1025.AB ) ,
    .I1 ( U1025.CD ) ,
    .I2 ( U1025.EF ) ) ;
and ( 
    .Z ( U459.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_53 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U459.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_0 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U459.EF ) ,
    .I0 ( xor_decoded_masks_10_0 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_0 ) ,
    .I0 ( U459.AB ) ,
    .I1 ( U459.CD ) ,
    .I2 ( U459.EF ) ) ;
and ( 
    .Z ( U770.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_62 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U770.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_9 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U770.EF ) ,
    .I0 ( xor_decoded_masks_6_9 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_9 ) ,
    .I0 ( U770.AB ) ,
    .I1 ( U770.CD ) ,
    .I2 ( U770.EF ) ) ;
and ( 
    .Z ( U773.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_88 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U773.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_35 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U773.EF ) ,
    .I0 ( xor_decoded_masks_8_35 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_35 ) ,
    .I0 ( U773.AB ) ,
    .I1 ( U773.CD ) ,
    .I2 ( U773.EF ) ) ;
and ( 
    .Z ( U1023.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_89 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1023.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_36 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1023.EF ) ,
    .I0 ( xor_decoded_masks_12_36 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_36 ) ,
    .I0 ( U1023.AB ) ,
    .I1 ( U1023.CD ) ,
    .I2 ( U1023.EF ) ) ;
and ( 
    .Z ( U1309.AB ) ,
    .I0 ( n37 ) ,
    .I1 ( masks_shift_reg_3_9 ) ) ;
and ( 
    .Z ( U1309.CD ) ,
    .I0 ( masks_shift_reg_3_0 ) ,
    .I1 ( n39 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_3 ) ,
    .I0 ( U1309.AB ) ,
    .I1 ( U1309.CD ) ) ;
and ( 
    .Z ( U772.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_72 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U772.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_19 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U772.EF ) ,
    .I0 ( xor_decoded_masks_6_19 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_19 ) ,
    .I0 ( U772.AB ) ,
    .I1 ( U772.CD ) ,
    .I2 ( U772.EF ) ) ;
and ( 
    .Z ( U1020.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_20 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1020.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_20 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1020.EF ) ,
    .I0 ( xor_decoded_masks_11_20 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_20 ) ,
    .I0 ( U1020.AB ) ,
    .I1 ( U1020.CD ) ,
    .I2 ( U1020.EF ) ) ;
and ( 
    .Z ( U1308.AB ) ,
    .I0 ( n40 ) ,
    .I1 ( masks_shift_reg_7_9 ) ) ;
and ( 
    .Z ( U1308.CD ) ,
    .I0 ( masks_shift_reg_7_0 ) ,
    .I1 ( n43 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_7 ) ,
    .I0 ( U1308.AB ) ,
    .I1 ( U1308.CD ) ) ;
and ( 
    .Z ( U1021.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_14 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1021.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_14 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1021.EF ) ,
    .I0 ( xor_decoded_masks_11_14 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_14 ) ,
    .I0 ( U1021.AB ) ,
    .I1 ( U1021.CD ) ,
    .I2 ( U1021.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_12_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_12_10 ) ,
    .IN ( masks_hold_reg_12_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_12_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_12_reg_10.QT ) ,
    .I1 ( masks_hold_reg_12_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_12_reg_10.ED ) ,
    .S ( masks_hold_reg_12_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_12_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_12_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_12_reg_10.ED ) ,
    .I1 ( masks_hold_reg_12_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_12_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_12_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_12_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_12_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_12_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_12_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_12_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_12_reg_10.QT ) ) ;
and ( 
    .Z ( U779.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_80 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U779.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_27 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U779.EF ) ,
    .I0 ( xor_decoded_masks_10_27 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_27 ) ,
    .I0 ( U779.AB ) ,
    .I1 ( U779.CD ) ,
    .I2 ( U779.EF ) ) ;
and ( 
    .Z ( U778.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_88 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U778.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_35 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U778.EF ) ,
    .I0 ( xor_decoded_masks_10_35 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_35 ) ,
    .I0 ( U778.AB ) ,
    .I1 ( U778.CD ) ,
    .I2 ( U778.EF ) ) ;
and ( 
    .Z ( U500.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_5 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U500.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_5 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U500.EF ) ,
    .I0 ( xor_decoded_masks_0_5 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_5 ) ,
    .I0 ( U500.AB ) ,
    .I1 ( U500.CD ) ,
    .I2 ( U500.EF ) ) ;
and ( 
    .Z ( U1028.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_36 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1028.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_36 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1028.EF ) ,
    .I0 ( xor_decoded_masks_13_36 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_36 ) ,
    .I0 ( U1028.AB ) ,
    .I1 ( U1028.CD ) ,
    .I2 ( U1028.EF ) ) ;
and ( 
    .Z ( U501.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_4 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U501.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_4 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U501.EF ) ,
    .I0 ( xor_decoded_masks_0_4 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_4 ) ,
    .I0 ( U501.AB ) ,
    .I1 ( U501.CD ) ,
    .I2 ( U501.EF ) ) ;
and ( 
    .Z ( U1253.AB ) ,
    .I0 ( masks_hold_reg_4_1 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U1253.CD ) ,
    .I0 ( config1_xor_encoded_masks_52 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_52 ) ,
    .I0 ( U1253.AB ) ,
    .I1 ( U1253.CD ) ) ;
and ( 
    .Z ( U1029.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_20 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1029.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_20 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1029.EF ) ,
    .I0 ( xor_decoded_masks_13_20 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_20 ) ,
    .I0 ( U1029.AB ) ,
    .I1 ( U1029.CD ) ,
    .I2 ( U1029.EF ) ) ;
and ( 
    .Z ( U502.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_6 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U502.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_6 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U502.EF ) ,
    .I0 ( xor_decoded_masks_0_6 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_6 ) ,
    .I0 ( U502.AB ) ,
    .I1 ( U502.CD ) ,
    .I2 ( U502.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_6_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_10.CPI_ ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29286 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_6_10 ) ,
    .IN ( masks_hold_reg_6_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_6_reg_10.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_6_reg_10.QT ) ,
    .I1 ( masks_hold_reg_6_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_6_reg_10.ED ) ,
    .S ( masks_hold_reg_6_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_6_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_6_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_6_reg_10.ED ) ,
    .I1 ( masks_hold_reg_6_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_6_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_6_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_6_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_6_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_6_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_6_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_6_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_6_reg_10.QT ) ) ;
and ( 
    .Z ( U1252.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_7 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1252.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_7 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1252.EF ) ,
    .I0 ( xor_decoded_masks_0_7 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_7 ) ,
    .I0 ( U1252.AB ) ,
    .I1 ( U1252.CD ) ,
    .I2 ( U1252.EF ) ) ;
and ( 
    .Z ( U503.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_155 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U503.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_48 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U503.EF ) ,
    .I0 ( xor_decoded_masks_2_48 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_48 ) ,
    .I0 ( U503.AB ) ,
    .I1 ( U503.CD ) ,
    .I2 ( U503.EF ) ) ;
and ( 
    .Z ( U1251.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_53 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1251.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_53 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1251.EF ) ,
    .I0 ( xor_decoded_masks_0_53 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_53 ) ,
    .I0 ( U1251.AB ) ,
    .I1 ( U1251.CD ) ,
    .I2 ( U1251.EF ) ) ;
and ( 
    .Z ( U504.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_48 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U504.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_48 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U504.EF ) ,
    .I0 ( xor_decoded_masks_3_48 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_48 ) ,
    .I0 ( U504.AB ) ,
    .I1 ( U504.CD ) ,
    .I2 ( U504.EF ) ) ;
and ( 
    .Z ( U1250.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_97 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1250.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_43 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1250.EF ) ,
    .I0 ( xor_decoded_masks_1_43 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_43 ) ,
    .I0 ( U1250.AB ) ,
    .I1 ( U1250.CD ) ,
    .I2 ( U1250.EF ) ) ;
and ( 
    .Z ( U505.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_101 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U505.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_48 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U505.EF ) ,
    .I0 ( xor_decoded_masks_4_48 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_48 ) ,
    .I0 ( U505.AB ) ,
    .I1 ( U505.CD ) ,
    .I2 ( U505.EF ) ) ;
and ( 
    .Z ( U1257.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_51 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1257.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_51 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1257.EF ) ,
    .I0 ( xor_decoded_masks_3_51 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_51 ) ,
    .I0 ( U1257.AB ) ,
    .I1 ( U1257.CD ) ,
    .I2 ( U1257.EF ) ) ;
and ( 
    .Z ( U479.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_59 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U479.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_6 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U479.EF ) ,
    .I0 ( xor_decoded_masks_14_6 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_6 ) ,
    .I0 ( U479.AB ) ,
    .I1 ( U479.CD ) ,
    .I2 ( U479.EF ) ) ;
and ( 
    .Z ( U522.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_102 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U522.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_49 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U522.EF ) ,
    .I0 ( xor_decoded_masks_10_49 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_49 ) ,
    .I0 ( U522.AB ) ,
    .I1 ( U522.CD ) ,
    .I2 ( U522.EF ) ) ;
and ( 
    .Z ( U523.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_49 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U523.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_49 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U523.EF ) ,
    .I0 ( xor_decoded_masks_11_49 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_49 ) ,
    .I0 ( U523.AB ) ,
    .I1 ( U523.CD ) ,
    .I2 ( U523.EF ) ) ;
and ( 
    .Z ( U1271.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_52 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1271.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_52 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1271.EF ) ,
    .I0 ( xor_decoded_masks_9_52 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_52 ) ,
    .I0 ( U1271.AB ) ,
    .I1 ( U1271.CD ) ,
    .I2 ( U1271.EF ) ) ;
and ( 
    .Z ( U520.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_102 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U520.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_49 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U520.EF ) ,
    .I0 ( xor_decoded_masks_8_49 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_49 ) ,
    .I0 ( U520.AB ) ,
    .I1 ( U520.CD ) ,
    .I2 ( U520.EF ) ) ;
and ( 
    .Z ( U1270.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_105 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1270.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_52 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1270.EF ) ,
    .I0 ( xor_decoded_masks_8_52 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_52 ) ,
    .I0 ( U1270.AB ) ,
    .I1 ( U1270.CD ) ,
    .I2 ( U1270.EF ) ) ;
and ( 
    .Z ( U521.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_49 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U521.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_49 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U521.EF ) ,
    .I0 ( xor_decoded_masks_9_49 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_49 ) ,
    .I0 ( U521.AB ) ,
    .I1 ( U521.CD ) ,
    .I2 ( U521.EF ) ) ;
and ( 
    .Z ( U1273.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_52 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1273.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_52 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1273.EF ) ,
    .I0 ( xor_decoded_masks_11_52 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_52 ) ,
    .I0 ( U1273.AB ) ,
    .I1 ( U1273.CD ) ,
    .I2 ( U1273.EF ) ) ;
and ( 
    .Z ( U526.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_102 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U526.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_49 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U526.EF ) ,
    .I0 ( xor_decoded_masks_14_49 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_49 ) ,
    .I0 ( U526.AB ) ,
    .I1 ( U526.CD ) ,
    .I2 ( U526.EF ) ) ;
and ( 
    .Z ( U1272.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_105 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1272.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_52 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1272.EF ) ,
    .I0 ( xor_decoded_masks_10_52 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_52 ) ,
    .I0 ( U1272.AB ) ,
    .I1 ( U1272.CD ) ,
    .I2 ( U1272.EF ) ) ;
and ( 
    .Z ( U527.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_103 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U527.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_49 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U527.EF ) ,
    .I0 ( xor_decoded_masks_1_49 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_49 ) ,
    .I0 ( U527.AB ) ,
    .I1 ( U527.CD ) ,
    .I2 ( U527.EF ) ) ;
and ( 
    .Z ( U1275.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_52 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1275.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_52 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1275.EF ) ,
    .I0 ( xor_decoded_masks_13_52 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_52 ) ,
    .I0 ( U1275.AB ) ,
    .I1 ( U1275.CD ) ,
    .I2 ( U1275.EF ) ) ;
and ( 
    .Z ( U524.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_102 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U524.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_49 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U524.EF ) ,
    .I0 ( xor_decoded_masks_12_49 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_49 ) ,
    .I0 ( U524.AB ) ,
    .I1 ( U524.CD ) ,
    .I2 ( U524.EF ) ) ;
and ( 
    .Z ( U1274.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_105 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1274.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_52 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1274.EF ) ,
    .I0 ( xor_decoded_masks_12_52 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_52 ) ,
    .I0 ( U1274.AB ) ,
    .I1 ( U1274.CD ) ,
    .I2 ( U1274.EF ) ) ;
and ( 
    .Z ( U525.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_49 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U525.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_49 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U525.EF ) ,
    .I0 ( xor_decoded_masks_13_49 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_49 ) ,
    .I0 ( U525.AB ) ,
    .I1 ( U525.CD ) ,
    .I2 ( U525.EF ) ) ;
and ( 
    .Z ( U1277.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_106 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1277.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_52 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1277.EF ) ,
    .I0 ( xor_decoded_masks_1_52 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_52 ) ,
    .I0 ( U1277.AB ) ,
    .I1 ( U1277.CD ) ,
    .I2 ( U1277.EF ) ) ;
and ( 
    .Z ( U1276.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_105 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1276.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_52 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1276.EF ) ,
    .I0 ( xor_decoded_masks_14_52 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_52 ) ,
    .I0 ( U1276.AB ) ,
    .I1 ( U1276.CD ) ,
    .I2 ( U1276.EF ) ) ;
and ( 
    .Z ( U1279.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_50 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1279.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_50 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1279.EF ) ,
    .I0 ( xor_decoded_masks_3_50 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_50 ) ,
    .I0 ( U1279.AB ) ,
    .I1 ( U1279.CD ) ,
    .I2 ( U1279.EF ) ) ;
and ( 
    .Z ( U445.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_60 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U445.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_7 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U445.EF ) ,
    .I0 ( xor_decoded_masks_8_7 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_7 ) ,
    .I0 ( U445.AB ) ,
    .I1 ( U445.CD ) ,
    .I2 ( U445.EF ) ) ;
and ( 
    .Z ( U528.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_20 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U528.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_20 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U528.EF ) ,
    .I0 ( xor_decoded_masks_3_20 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_20 ) ,
    .I0 ( U528.AB ) ,
    .I1 ( U528.CD ) ,
    .I2 ( U528.EF ) ) ;
and ( 
    .Z ( U1278.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_157 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1278.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_50 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1278.EF ) ,
    .I0 ( xor_decoded_masks_2_50 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_50 ) ,
    .I0 ( U1278.AB ) ,
    .I1 ( U1278.CD ) ,
    .I2 ( U1278.EF ) ) ;
and ( 
    .Z ( U444.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_58 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U444.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_5 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U444.EF ) ,
    .I0 ( xor_decoded_masks_8_5 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_5 ) ,
    .I0 ( U444.AB ) ,
    .I1 ( U444.CD ) ,
    .I2 ( U444.EF ) ) ;
not ( 
    .O1 ( n7 ) ,
    .IN ( masks_shift_reg_8_0 ) ) ;
and ( 
    .Z ( U529.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_73 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U529.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_20 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U529.EF ) ,
    .I0 ( xor_decoded_masks_4_20 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_20 ) ,
    .I0 ( U529.AB ) ,
    .I1 ( U529.CD ) ,
    .I2 ( U529.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_11_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_8.CDNI_ ) ,
    .IN ( n52 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_8.CD ) ,
    .IN ( masks_shift_reg_11_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_8 ) ) ;
and ( 
    .Z ( U447.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_53 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U447.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_0 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U447.EF ) ,
    .I0 ( xor_decoded_masks_8_0 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_0 ) ,
    .I0 ( U447.AB ) ,
    .I1 ( U447.CD ) ,
    .I2 ( U447.EF ) ) ;
not ( 
    .O1 ( n9 ) ,
    .IN ( masks_shift_reg_6_0 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_11_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_1_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_9.CDNI_ ) ,
    .IN ( edt_update_hfs_netlink_29289 ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_9.CD ) ,
    .IN ( masks_shift_reg_11_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_11_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_11_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_11_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_11_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_11_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_11_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_11_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_11_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_11_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_11_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_11_9 ) ) ;
and ( 
    .Z ( U446.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_59 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U446.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_6 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U446.EF ) ,
    .I0 ( xor_decoded_masks_8_6 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_6 ) ,
    .I0 ( U446.AB ) ,
    .I1 ( U446.CD ) ,
    .I2 ( U446.EF ) ) ;
not ( 
    .O1 ( n12 ) ,
    .IN ( masks_shift_reg_2_0 ) ) ;
and ( 
    .Z ( U441.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_7 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U441.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_7 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U441.EF ) ,
    .I0 ( xor_decoded_masks_7_7 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_7 ) ,
    .I0 ( U441.AB ) ,
    .I1 ( U441.CD ) ,
    .I2 ( U441.EF ) ) ;
not ( 
    .O1 ( n15 ) ,
    .IN ( masks_shift_reg_10_0 ) ) ;
and ( 
    .Z ( U440.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_4 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U440.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_4 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U440.EF ) ,
    .I0 ( xor_decoded_masks_7_4 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_4 ) ,
    .I0 ( U440.AB ) ,
    .I1 ( U440.CD ) ,
    .I2 ( U440.EF ) ) ;
not ( 
    .O1 ( n11 ) ,
    .IN ( masks_shift_reg_4_0 ) ) ;
and ( 
    .Z ( U443.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_2 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U443.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_2 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U443.EF ) ,
    .I0 ( xor_decoded_masks_7_2 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_2 ) ,
    .I0 ( U443.AB ) ,
    .I1 ( U443.CD ) ,
    .I2 ( U443.EF ) ) ;
not ( 
    .O1 ( n16 ) ,
    .IN ( masks_shift_reg_0_0 ) ) ;
and ( 
    .Z ( U442.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_0 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U442.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_0 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U442.EF ) ,
    .I0 ( xor_decoded_masks_7_0 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_0 ) ,
    .I0 ( U442.AB ) ,
    .I1 ( U442.CD ) ,
    .I2 ( U442.EF ) ) ;
and ( 
    .Z ( U1310.AB ) ,
    .I0 ( n41 ) ,
    .I1 ( masks_shift_reg_5_9 ) ) ;
and ( 
    .Z ( U1310.CD ) ,
    .I0 ( masks_shift_reg_5_0 ) ,
    .I1 ( n44 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_5 ) ,
    .I0 ( U1310.AB ) ,
    .I1 ( U1310.CD ) ) ;
and ( 
    .Z ( U1311.AB ) ,
    .I0 ( masks_shift_reg_1_0 ) ,
    .I1 ( n44 ) ) ;
not ( 
    .O1 ( U1311.CN ) ,
    .IN ( n13 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_1 ) ,
    .I0 ( U1311.AB ) ,
    .I1 ( U1311.CN ) ) ;
and ( 
    .Z ( U764.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_92 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U764.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_39 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U764.EF ) ,
    .I0 ( xor_decoded_masks_4_39 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_39 ) ,
    .I0 ( U764.AB ) ,
    .I1 ( U764.CD ) ,
    .I2 ( U764.EF ) ) ;
and ( 
    .Z ( U765.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_62 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U765.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_9 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U765.EF ) ,
    .I0 ( xor_decoded_masks_4_9 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_9 ) ,
    .I0 ( U765.AB ) ,
    .I1 ( U765.CD ) ,
    .I2 ( U765.EF ) ) ;
and ( 
    .Z ( U1015.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_67 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1015.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_14 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1015.EF ) ,
    .I0 ( xor_decoded_masks_10_14 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_14 ) ,
    .I0 ( U1015.AB ) ,
    .I1 ( U1015.CD ) ,
    .I2 ( U1015.EF ) ) ;
and ( 
    .Z ( U429.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_7 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U429.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_7 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U429.EF ) ,
    .I0 ( xor_decoded_masks_5_7 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_7 ) ,
    .I0 ( U429.AB ) ,
    .I1 ( U429.CD ) ,
    .I2 ( U429.EF ) ) ;
and ( 
    .Z ( U744.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_78 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U744.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_25 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U744.EF ) ,
    .I0 ( xor_decoded_masks_14_25 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_25 ) ,
    .I0 ( U744.AB ) ,
    .I1 ( U744.CD ) ,
    .I2 ( U744.EF ) ) ;
and ( 
    .Z ( U1014.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_89 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1014.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_36 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1014.EF ) ,
    .I0 ( xor_decoded_masks_10_36 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_36 ) ,
    .I0 ( U1014.AB ) ,
    .I1 ( U1014.CD ) ,
    .I2 ( U1014.EF ) ) ;
and ( 
    .Z ( U428.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_55 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U428.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_2 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U428.EF ) ,
    .I0 ( xor_decoded_masks_4_2 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_2 ) ,
    .I0 ( U428.AB ) ,
    .I1 ( U428.CD ) ,
    .I2 ( U428.EF ) ) ;
and ( 
    .Z ( U745.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_90 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U745.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_37 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U745.EF ) ,
    .I0 ( xor_decoded_masks_14_37 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_37 ) ,
    .I0 ( U745.AB ) ,
    .I1 ( U745.CD ) ,
    .I2 ( U745.EF ) ) ;
and ( 
    .Z ( U1017.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_69 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1017.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_16 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1017.EF ) ,
    .I0 ( xor_decoded_masks_10_16 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_16 ) ,
    .I0 ( U1017.AB ) ,
    .I1 ( U1017.CD ) ,
    .I2 ( U1017.EF ) ) ;
and ( 
    .Z ( U742.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_82 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U742.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_29 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U742.EF ) ,
    .I0 ( xor_decoded_masks_14_29 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_29 ) ,
    .I0 ( U742.AB ) ,
    .I1 ( U742.CD ) ,
    .I2 ( U742.EF ) ) ;
and ( 
    .Z ( U1016.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_63 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1016.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_10 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1016.EF ) ,
    .I0 ( xor_decoded_masks_10_10 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_10 ) ,
    .I0 ( U1016.AB ) ,
    .I1 ( U1016.CD ) ,
    .I2 ( U1016.EF ) ) ;
and ( 
    .Z ( U743.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_86 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U743.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_33 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U743.EF ) ,
    .I0 ( xor_decoded_masks_14_33 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_33 ) ,
    .I0 ( U743.AB ) ,
    .I1 ( U743.CD ) ,
    .I2 ( U743.EF ) ) ;
and ( 
    .Z ( U1011.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_36 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1011.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_36 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1011.EF ) ,
    .I0 ( xor_decoded_masks_9_36 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_36 ) ,
    .I0 ( U1011.AB ) ,
    .I1 ( U1011.CD ) ,
    .I2 ( U1011.EF ) ) ;
and ( 
    .Z ( U740.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_78 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U740.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_25 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U740.EF ) ,
    .I0 ( xor_decoded_masks_12_25 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_25 ) ,
    .I0 ( U740.AB ) ,
    .I1 ( U740.CD ) ,
    .I2 ( U740.EF ) ) ;
and ( 
    .Z ( U1010.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_32 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1010.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_32 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1010.EF ) ,
    .I0 ( xor_decoded_masks_9_32 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_32 ) ,
    .I0 ( U1010.AB ) ,
    .I1 ( U1010.CD ) ,
    .I2 ( U1010.EF ) ) ;
and ( 
    .Z ( U741.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_90 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U741.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_37 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U741.EF ) ,
    .I0 ( xor_decoded_masks_12_37 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_37 ) ,
    .I0 ( U741.AB ) ,
    .I1 ( U741.CD ) ,
    .I2 ( U741.EF ) ) ;
and ( 
    .Z ( U1013.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_10 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1013.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_10 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1013.EF ) ,
    .I0 ( xor_decoded_masks_9_10 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_10 ) ,
    .I0 ( U1013.AB ) ,
    .I1 ( U1013.CD ) ,
    .I2 ( U1013.EF ) ) ;
and ( 
    .Z ( U1012.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_20 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1012.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_20 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1012.EF ) ,
    .I0 ( xor_decoded_masks_9_20 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_20 ) ,
    .I0 ( U1012.AB ) ,
    .I1 ( U1012.CD ) ,
    .I2 ( U1012.EF ) ) ;
and ( 
    .Z ( U665.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_133 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U665.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_26 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U665.EF ) ,
    .I0 ( xor_decoded_masks_2_26 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_26 ) ,
    .I0 ( U665.AB ) ,
    .I1 ( U665.CD ) ,
    .I2 ( U665.EF ) ) ;
and ( 
    .Z ( U664.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_64 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U664.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_10 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U664.EF ) ,
    .I0 ( xor_decoded_masks_1_10 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_10 ) ,
    .I0 ( U664.AB ) ,
    .I1 ( U664.CD ) ,
    .I2 ( U664.EF ) ) ;
and ( 
    .Z ( U1136.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_11 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1136.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_11 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1136.EF ) ,
    .I0 ( xor_decoded_masks_7_11 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_11 ) ,
    .I0 ( U1136.AB ) ,
    .I1 ( U1136.CD ) ,
    .I2 ( U1136.EF ) ) ;
and ( 
    .Z ( U667.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_145 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U667.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_38 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U667.EF ) ,
    .I0 ( xor_decoded_masks_2_38 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_38 ) ,
    .I0 ( U667.AB ) ,
    .I1 ( U667.CD ) ,
    .I2 ( U667.EF ) ) ;
and ( 
    .Z ( U1137.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_29 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1137.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_29 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1137.EF ) ,
    .I0 ( xor_decoded_masks_9_29 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_29 ) ,
    .I0 ( U1137.AB ) ,
    .I1 ( U1137.CD ) ,
    .I2 ( U1137.EF ) ) ;
and ( 
    .Z ( U666.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_141 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U666.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_34 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U666.EF ) ,
    .I0 ( xor_decoded_masks_2_34 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_34 ) ,
    .I0 ( U666.AB ) ,
    .I1 ( U666.CD ) ,
    .I2 ( U666.EF ) ) ;
and ( 
    .Z ( U1134.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_21 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1134.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_21 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1134.EF ) ,
    .I0 ( xor_decoded_masks_7_21 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_21 ) ,
    .I0 ( U1134.AB ) ,
    .I1 ( U1134.CD ) ,
    .I2 ( U1134.EF ) ) ;
and ( 
    .Z ( U1019.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_36 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1019.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_36 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1019.EF ) ,
    .I0 ( xor_decoded_masks_11_36 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_36 ) ,
    .I0 ( U1019.AB ) ,
    .I1 ( U1019.CD ) ,
    .I2 ( U1019.EF ) ) ;
and ( 
    .Z ( U968.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_58 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U968.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_5 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U968.EF ) ,
    .I0 ( xor_decoded_masks_14_5 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_5 ) ,
    .I0 ( U968.AB ) ,
    .I1 ( U968.CD ) ,
    .I2 ( U968.EF ) ) ;
and ( 
    .Z ( U661.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_86 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U661.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_32 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U661.EF ) ,
    .I0 ( xor_decoded_masks_1_32 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_32 ) ,
    .I0 ( U661.AB ) ,
    .I1 ( U661.CD ) ,
    .I2 ( U661.EF ) ) ;
and ( 
    .Z ( U1135.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_15 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1135.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_15 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1135.EF ) ,
    .I0 ( xor_decoded_masks_7_15 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_15 ) ,
    .I0 ( U1135.AB ) ,
    .I1 ( U1135.CD ) ,
    .I2 ( U1135.EF ) ) ;
and ( 
    .Z ( U748.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_79 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U748.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_25 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U748.EF ) ,
    .I0 ( xor_decoded_masks_1_25 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_25 ) ,
    .I0 ( U748.AB ) ,
    .I1 ( U748.CD ) ,
    .I2 ( U748.EF ) ) ;
and ( 
    .Z ( U511.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_101 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U511.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_48 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U511.EF ) ,
    .I0 ( xor_decoded_masks_10_48 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_48 ) ,
    .I0 ( U511.AB ) ,
    .I1 ( U511.CD ) ,
    .I2 ( U511.EF ) ) ;
or ( 
    .Z ( U969.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_6 ) ) ;
not ( 
    .O1 ( U969.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_12 ) ) ;
not ( 
    .O1 ( U969.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U969.not_c_tempD ) ,
    .I0 ( U969.not_c_temp ) ,
    .I1 ( U969.ND ) ) ;
and ( 
    .Z ( U969.ZN ) ,
    .I0 ( U969.AB ) ,
    .I1 ( U969.not_c_tempD ) ) ;
not ( 
    .O1 ( N234 ) ,
    .IN ( U969.ZN ) ) ;
and ( 
    .Z ( U660.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_78 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U660.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_24 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U660.EF ) ,
    .I0 ( xor_decoded_masks_1_24 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_24 ) ,
    .I0 ( U660.AB ) ,
    .I1 ( U660.CD ) ,
    .I2 ( U660.EF ) ) ;
and ( 
    .Z ( U1132.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_37 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1132.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_37 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1132.EF ) ,
    .I0 ( xor_decoded_masks_7_37 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_37 ) ,
    .I0 ( U1132.AB ) ,
    .I1 ( U1132.CD ) ,
    .I2 ( U1132.EF ) ) ;
and ( 
    .Z ( U749.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_87 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U749.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_33 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U749.EF ) ,
    .I0 ( xor_decoded_masks_1_33 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_33 ) ,
    .I0 ( U749.AB ) ,
    .I1 ( U749.CD ) ,
    .I2 ( U749.EF ) ) ;
and ( 
    .Z ( U510.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_48 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U510.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_48 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U510.EF ) ,
    .I0 ( xor_decoded_masks_9_48 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_48 ) ,
    .I0 ( U510.AB ) ,
    .I1 ( U510.CD ) ,
    .I2 ( U510.EF ) ) ;
and ( 
    .Z ( U1242.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_43 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1242.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_43 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1242.EF ) ,
    .I0 ( xor_decoded_masks_7_43 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_43 ) ,
    .I0 ( U1242.AB ) ,
    .I1 ( U1242.CD ) ,
    .I2 ( U1242.EF ) ) ;
and ( 
    .Z ( U663.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_74 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U663.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_20 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U663.EF ) ,
    .I0 ( xor_decoded_masks_1_20 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_20 ) ,
    .I0 ( U663.AB ) ,
    .I1 ( U663.CD ) ,
    .I2 ( U663.EF ) ) ;
and ( 
    .Z ( U1133.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_17 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1133.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_17 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1133.EF ) ,
    .I0 ( xor_decoded_masks_7_17 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_17 ) ,
    .I0 ( U1133.AB ) ,
    .I1 ( U1133.CD ) ,
    .I2 ( U1133.EF ) ) ;
and ( 
    .Z ( U513.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_101 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U513.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_48 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U513.EF ) ,
    .I0 ( xor_decoded_masks_14_48 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_48 ) ,
    .I0 ( U513.AB ) ,
    .I1 ( U513.CD ) ,
    .I2 ( U513.EF ) ) ;
and ( 
    .Z ( U1243.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_96 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1243.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_43 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1243.EF ) ,
    .I0 ( xor_decoded_masks_8_43 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_43 ) ,
    .I0 ( U1243.AB ) ,
    .I1 ( U1243.CD ) ,
    .I2 ( U1243.EF ) ) ;
and ( 
    .Z ( U662.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_90 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U662.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_36 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U662.EF ) ,
    .I0 ( xor_decoded_masks_1_36 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_36 ) ,
    .I0 ( U662.AB ) ,
    .I1 ( U662.CD ) ,
    .I2 ( U662.EF ) ) ;
and ( 
    .Z ( U1130.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_25 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1130.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_25 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1130.EF ) ,
    .I0 ( xor_decoded_masks_7_25 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_25 ) ,
    .I0 ( U1130.AB ) ,
    .I1 ( U1130.CD ) ,
    .I2 ( U1130.EF ) ) ;
and ( 
    .Z ( U512.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_48 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U512.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_48 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U512.EF ) ,
    .I0 ( xor_decoded_masks_13_48 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_48 ) ,
    .I0 ( U512.AB ) ,
    .I1 ( U512.CD ) ,
    .I2 ( U512.EF ) ) ;
and ( 
    .Z ( U1240.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_43 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1240.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_43 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1240.EF ) ,
    .I0 ( xor_decoded_masks_5_43 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_43 ) ,
    .I0 ( U1240.AB ) ,
    .I1 ( U1240.CD ) ,
    .I2 ( U1240.EF ) ) ;
and ( 
    .Z ( U1131.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_33 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1131.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_33 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1131.EF ) ,
    .I0 ( xor_decoded_masks_7_33 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_33 ) ,
    .I0 ( U1131.AB ) ,
    .I1 ( U1131.CD ) ,
    .I2 ( U1131.EF ) ) ;
and ( 
    .Z ( U515.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_156 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U515.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_49 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U515.EF ) ,
    .I0 ( xor_decoded_masks_2_49 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_49 ) ,
    .I0 ( U515.AB ) ,
    .I1 ( U515.CD ) ,
    .I2 ( U515.EF ) ) ;
and ( 
    .Z ( U1241.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_96 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1241.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_43 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1241.EF ) ,
    .I0 ( xor_decoded_masks_6_43 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_43 ) ,
    .I0 ( U1241.AB ) ,
    .I1 ( U1241.CD ) ,
    .I2 ( U1241.EF ) ) ;
and ( 
    .Z ( U514.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_102 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U514.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_48 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U514.EF ) ,
    .I0 ( xor_decoded_masks_1_48 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_48 ) ,
    .I0 ( U514.AB ) ,
    .I1 ( U514.CD ) ,
    .I2 ( U514.EF ) ) ;
and ( 
    .Z ( U1246.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_43 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1246.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_43 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1246.EF ) ,
    .I0 ( xor_decoded_masks_11_43 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_43 ) ,
    .I0 ( U1246.AB ) ,
    .I1 ( U1246.CD ) ,
    .I2 ( U1246.EF ) ) ;
and ( 
    .Z ( U962.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_1 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U962.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_1 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U962.EF ) ,
    .I0 ( xor_decoded_masks_11_1 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_1 ) ,
    .I0 ( U962.AB ) ,
    .I1 ( U962.CD ) ,
    .I2 ( U962.EF ) ) ;
and ( 
    .Z ( U517.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_49 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U517.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_49 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U517.EF ) ,
    .I0 ( xor_decoded_masks_5_49 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_49 ) ,
    .I0 ( U517.AB ) ,
    .I1 ( U517.CD ) ,
    .I2 ( U517.EF ) ) ;
and ( 
    .Z ( U1247.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_96 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1247.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_43 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1247.EF ) ,
    .I0 ( xor_decoded_masks_12_43 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_43 ) ,
    .I0 ( U1247.AB ) ,
    .I1 ( U1247.CD ) ,
    .I2 ( U1247.EF ) ) ;
and ( 
    .Z ( U963.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_98 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U963.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_45 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U963.EF ) ,
    .I0 ( xor_decoded_masks_12_45 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_45 ) ,
    .I0 ( U963.AB ) ,
    .I1 ( U963.CD ) ,
    .I2 ( U963.EF ) ) ;
and ( 
    .Z ( U516.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_102 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U516.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_49 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U516.EF ) ,
    .I0 ( xor_decoded_masks_4_49 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_49 ) ,
    .I0 ( U516.AB ) ,
    .I1 ( U516.CD ) ,
    .I2 ( U516.EF ) ) ;
and ( 
    .Z ( U1244.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_43 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1244.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_43 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1244.EF ) ,
    .I0 ( xor_decoded_masks_9_43 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_43 ) ,
    .I0 ( U1244.AB ) ,
    .I1 ( U1244.CD ) ,
    .I2 ( U1244.EF ) ) ;
and ( 
    .Z ( U960.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_45 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U960.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_45 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U960.EF ) ,
    .I0 ( xor_decoded_masks_11_45 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_45 ) ,
    .I0 ( U960.AB ) ,
    .I1 ( U960.CD ) ,
    .I2 ( U960.EF ) ) ;
and ( 
    .Z ( U669.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_115 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U669.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_8 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U669.EF ) ,
    .I0 ( xor_decoded_masks_2_8 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_8 ) ,
    .I0 ( U669.AB ) ,
    .I1 ( U669.CD ) ,
    .I2 ( U669.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_9_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_1.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_1.CD ) ,
    .IN ( masks_shift_reg_9_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_1 ) ) ;
and ( 
    .Z ( U519.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_49 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U519.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_49 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U519.EF ) ,
    .I0 ( xor_decoded_masks_7_49 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_49 ) ,
    .I0 ( U519.AB ) ,
    .I1 ( U519.CD ) ,
    .I2 ( U519.EF ) ) ;
and ( 
    .Z ( U1245.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_96 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1245.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_43 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1245.EF ) ,
    .I0 ( xor_decoded_masks_10_43 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_43 ) ,
    .I0 ( U1245.AB ) ,
    .I1 ( U1245.CD ) ,
    .I2 ( U1245.EF ) ) ;
and ( 
    .Z ( U961.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_5 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U961.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_5 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U961.EF ) ,
    .I0 ( xor_decoded_masks_11_5 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_5 ) ,
    .I0 ( U961.AB ) ,
    .I1 ( U961.CD ) ,
    .I2 ( U961.EF ) ) ;
and ( 
    .Z ( U668.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_125 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U668.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_18 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U668.EF ) ,
    .I0 ( xor_decoded_masks_2_18 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_18 ) ,
    .I0 ( U668.AB ) ,
    .I1 ( U668.CD ) ,
    .I2 ( U668.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_9_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_0.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_0.CD ) ,
    .IN ( masks_shift_reg_9_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_0 ) ) ;
and ( 
    .Z ( U518.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_102 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U518.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_49 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U518.EF ) ,
    .I0 ( xor_decoded_masks_6_49 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_49 ) ,
    .I0 ( U518.AB ) ,
    .I1 ( U518.CD ) ,
    .I2 ( U518.EF ) ) ;
and ( 
    .Z ( U966.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_1 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U966.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_1 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U966.EF ) ,
    .I0 ( xor_decoded_masks_13_1 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_1 ) ,
    .I0 ( U966.AB ) ,
    .I1 ( U966.CD ) ,
    .I2 ( U966.EF ) ) ;
and ( 
    .Z ( U432.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_3 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U432.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_3 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U432.EF ) ,
    .I0 ( xor_decoded_masks_5_3 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_3 ) ,
    .I0 ( U432.AB ) ,
    .I1 ( U432.CD ) ,
    .I2 ( U432.EF ) ) ;
and ( 
    .Z ( U1261.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_51 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1261.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_51 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1261.EF ) ,
    .I0 ( xor_decoded_masks_9_51 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_51 ) ,
    .I0 ( U1261.AB ) ,
    .I1 ( U1261.CD ) ,
    .I2 ( U1261.EF ) ) ;
and ( 
    .Z ( U530.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_73 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U530.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_20 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U530.EF ) ,
    .I0 ( xor_decoded_masks_6_20 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_20 ) ,
    .I0 ( U530.AB ) ,
    .I1 ( U530.CD ) ,
    .I2 ( U530.EF ) ) ;
and ( 
    .Z ( U1262.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_104 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1262.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_51 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1262.EF ) ,
    .I0 ( xor_decoded_masks_10_51 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_51 ) ,
    .I0 ( U1262.AB ) ,
    .I1 ( U1262.CD ) ,
    .I2 ( U1262.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_0_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_8.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_8.CD ) ,
    .IN ( masks_shift_reg_0_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_8 ) ) ;
and ( 
    .Z ( U537.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_2 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U537.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_2 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U537.EF ) ,
    .I0 ( xor_decoded_masks_11_2 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_2 ) ,
    .I0 ( U537.AB ) ,
    .I1 ( U537.CD ) ,
    .I2 ( U537.EF ) ) ;
and ( 
    .Z ( U1263.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_51 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1263.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_51 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1263.EF ) ,
    .I0 ( xor_decoded_masks_13_51 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_51 ) ,
    .I0 ( U1263.AB ) ,
    .I1 ( U1263.CD ) ,
    .I2 ( U1263.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_0_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_9.CPI_ ) ,
    .IN ( edt_clock ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_9.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_9.CD ) ,
    .IN ( masks_shift_reg_0_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_9 ) ) ;
and ( 
    .Z ( U536.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_19 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U536.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_19 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U536.EF ) ,
    .I0 ( xor_decoded_masks_7_19 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_19 ) ,
    .I0 ( U536.AB ) ,
    .I1 ( U536.CD ) ,
    .I2 ( U536.EF ) ) ;
and ( 
    .Z ( U1264.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_159 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1264.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_52 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1264.EF ) ,
    .I0 ( xor_decoded_masks_2_52 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_52 ) ,
    .I0 ( U1264.AB ) ,
    .I1 ( U1264.CD ) ,
    .I2 ( U1264.EF ) ) ;
and ( 
    .Z ( U535.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_19 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U535.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_19 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U535.EF ) ,
    .I0 ( xor_decoded_masks_5_19 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_19 ) ,
    .I0 ( U535.AB ) ,
    .I1 ( U535.CD ) ,
    .I2 ( U535.EF ) ) ;
and ( 
    .Z ( U1265.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_52 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1265.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_52 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1265.EF ) ,
    .I0 ( xor_decoded_masks_3_52 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_52 ) ,
    .I0 ( U1265.AB ) ,
    .I1 ( U1265.CD ) ,
    .I2 ( U1265.EF ) ) ;
and ( 
    .Z ( U534.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_73 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U534.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_20 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U534.EF ) ,
    .I0 ( xor_decoded_masks_14_20 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_20 ) ,
    .I0 ( U534.AB ) ,
    .I1 ( U534.CD ) ,
    .I2 ( U534.EF ) ) ;
and ( 
    .Z ( U1266.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_105 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1266.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_52 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1266.EF ) ,
    .I0 ( xor_decoded_masks_4_52 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_52 ) ,
    .I0 ( U1266.AB ) ,
    .I1 ( U1266.CD ) ,
    .I2 ( U1266.EF ) ) ;
and ( 
    .Z ( U1267.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_52 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1267.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_52 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1267.EF ) ,
    .I0 ( xor_decoded_masks_5_52 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_52 ) ,
    .I0 ( U1267.AB ) ,
    .I1 ( U1267.CD ) ,
    .I2 ( U1267.EF ) ) ;
and ( 
    .Z ( U1268.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_105 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1268.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_52 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1268.EF ) ,
    .I0 ( xor_decoded_masks_6_52 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_52 ) ,
    .I0 ( U1268.AB ) ,
    .I1 ( U1268.CD ) ,
    .I2 ( U1268.EF ) ) ;
and ( 
    .Z ( U454.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_3 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U454.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_3 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U454.EF ) ,
    .I0 ( xor_decoded_masks_9_3 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_3 ) ,
    .I0 ( U454.AB ) ,
    .I1 ( U454.CD ) ,
    .I2 ( U454.EF ) ) ;
and ( 
    .Z ( U539.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_6 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U539.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_6 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U539.EF ) ,
    .I0 ( xor_decoded_masks_7_6 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_6 ) ,
    .I0 ( U539.AB ) ,
    .I1 ( U539.CD ) ,
    .I2 ( U539.EF ) ) ;
and ( 
    .Z ( U1269.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_52 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1269.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_52 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1269.EF ) ,
    .I0 ( xor_decoded_masks_7_52 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_52 ) ,
    .I0 ( U1269.AB ) ,
    .I1 ( U1269.CD ) ,
    .I2 ( U1269.EF ) ) ;
and ( 
    .Z ( U455.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_2 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U455.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_2 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U455.EF ) ,
    .I0 ( xor_decoded_masks_9_2 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_2 ) ,
    .I0 ( U455.AB ) ,
    .I1 ( U455.CD ) ,
    .I2 ( U455.EF ) ) ;
and ( 
    .Z ( U1307.AB ) ,
    .I0 ( edt_configuration_hfs_netlink_29290 ) ,
    .I1 ( masks_shift_reg_9_9 ) ) ;
and ( 
    .Z ( U1307.CD ) ,
    .I0 ( masks_shift_reg_9_0 ) ,
    .I1 ( n45 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_9 ) ,
    .I0 ( U1307.AB ) ,
    .I1 ( U1307.CD ) ) ;
and ( 
    .Z ( U538.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_4 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U538.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_4 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U538.EF ) ,
    .I0 ( xor_decoded_masks_5_4 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_4 ) ,
    .I0 ( U538.AB ) ,
    .I1 ( U538.CD ) ,
    .I2 ( U538.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_0_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_0.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_0.CD ) ,
    .IN ( masks_shift_reg_0_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_0 ) ) ;
and ( 
    .Z ( U456.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_57 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U456.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_4 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U456.EF ) ,
    .I0 ( xor_decoded_masks_10_4 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_4 ) ,
    .I0 ( U456.AB ) ,
    .I1 ( U456.CD ) ,
    .I2 ( U456.EF ) ) ;
and ( 
    .Z ( U1306.AB ) ,
    .I0 ( edt_configuration_hfs_netlink_29290 ) ,
    .I1 ( masks_shift_reg_11_9 ) ) ;
and ( 
    .Z ( U1306.CD ) ,
    .I0 ( masks_shift_reg_11_0 ) ,
    .I1 ( n45 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_11 ) ,
    .I0 ( U1306.AB ) ,
    .I1 ( U1306.CD ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_0_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_0_reg_1.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_1.CD ) ,
    .IN ( masks_shift_reg_0_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_0_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_0_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_0_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_0_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_0_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_0_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_0_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_0_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_0_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_0_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_0_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_0_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_0_1 ) ) ;
and ( 
    .Z ( U457.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_60 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U457.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_7 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U457.EF ) ,
    .I0 ( xor_decoded_masks_10_7 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_7 ) ,
    .I0 ( U457.AB ) ,
    .I1 ( U457.CD ) ,
    .I2 ( U457.EF ) ) ;
and ( 
    .Z ( U1305.AB ) ,
    .I0 ( edt_configuration_hfs_netlink_29290 ) ,
    .I1 ( masks_shift_reg_11_9 ) ) ;
and ( 
    .Z ( U1305.CD ) ,
    .I0 ( masks_shift_reg_12_0 ) ,
    .I1 ( n45 ) ) ;
or ( 
    .Z ( edt_channels_out_from_controller_12 ) ,
    .I0 ( U1305.AB ) ,
    .I1 ( U1305.CD ) ) ;
and ( 
    .Z ( U965.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_5 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U965.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_5 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U965.EF ) ,
    .I0 ( xor_decoded_masks_13_5 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_5 ) ,
    .I0 ( U965.AB ) ,
    .I1 ( U965.CD ) ,
    .I2 ( U965.EF ) ) ;
and ( 
    .Z ( U431.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_0 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U431.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_0 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U431.EF ) ,
    .I0 ( xor_decoded_masks_5_0 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_0 ) ,
    .I0 ( U431.AB ) ,
    .I1 ( U431.CD ) ,
    .I2 ( U431.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_9_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_4.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_4.CD ) ,
    .IN ( masks_shift_reg_9_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_4 ) ) ;
and ( 
    .Z ( U436.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_59 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U436.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_6 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U436.EF ) ,
    .I0 ( xor_decoded_masks_6_6 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_6 ) ,
    .I0 ( U436.AB ) ,
    .I1 ( U436.CD ) ,
    .I2 ( U436.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_7.DI_ ) ,
    .IN ( n77 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_7.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_7.CD ) ,
    .IN ( masks_shift_reg_9_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_7 ) ) ;
and ( 
    .Z ( U437.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_53 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U437.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_0 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U437.EF ) ,
    .I0 ( xor_decoded_masks_6_0 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_0 ) ,
    .I0 ( U437.AB ) ,
    .I1 ( U437.CD ) ,
    .I2 ( U437.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_9_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_6.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_6.CD ) ,
    .IN ( masks_shift_reg_9_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_3_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_9.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_9.CD ) ,
    .IN ( masks_shift_reg_3_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_9 ) ) ;
and ( 
    .Z ( U434.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_58 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U434.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_5 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U434.EF ) ,
    .I0 ( xor_decoded_masks_6_5 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_5 ) ,
    .I0 ( U434.AB ) ,
    .I1 ( U434.CD ) ,
    .I2 ( U434.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_9_10 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_9.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_9.CD ) ,
    .IN ( masks_shift_reg_9_reg_9.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_9.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_9.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_9.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_9.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_9.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_9.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_9.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_9.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_9.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_9.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_9.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_9.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_9 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_8.DI_ ) ,
    .IN ( n48 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_8.CDNI_ ) ,
    .IN ( masks_shift_reg_3_9 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_8.CD ) ,
    .IN ( masks_shift_reg_3_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_8 ) ) ;
and ( 
    .Z ( U435.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_60 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U435.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_7 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U435.EF ) ,
    .I0 ( xor_decoded_masks_6_7 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_7 ) ,
    .I0 ( U435.AB ) ,
    .I1 ( U435.CD ) ,
    .I2 ( U435.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_8.DI_ ) ,
    .IN ( n51 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_8.CDNI_ ) ,
    .IN ( masks_shift_reg_9_9 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_8.CD ) ,
    .IN ( masks_shift_reg_9_reg_8.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_8.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_8.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_8.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_8.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_8.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_8.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_8.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_8.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_8.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_8.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_8.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_8.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_8 ) ) ;
and ( 
    .Z ( U757.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_142 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U757.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_35 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U757.EF ) ,
    .I0 ( xor_decoded_masks_2_35 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_35 ) ,
    .I0 ( U757.AB ) ,
    .I1 ( U757.CD ) ,
    .I2 ( U757.EF ) ) ;
and ( 
    .Z ( U756.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_134 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U756.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_27 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U756.EF ) ,
    .I0 ( xor_decoded_masks_2_27 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_27 ) ,
    .I0 ( U756.AB ) ,
    .I1 ( U756.CD ) ,
    .I2 ( U756.EF ) ) ;
and ( 
    .Z ( U1004.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_32 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1004.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_32 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1004.EF ) ,
    .I0 ( xor_decoded_masks_7_32 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_32 ) ,
    .I0 ( U1004.AB ) ,
    .I1 ( U1004.CD ) ,
    .I2 ( U1004.EF ) ) ;
and ( 
    .Z ( U438.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_56 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U438.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_3 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U438.EF ) ,
    .I0 ( xor_decoded_masks_6_3 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_3 ) ,
    .I0 ( U438.AB ) ,
    .I1 ( U438.CD ) ,
    .I2 ( U438.EF ) ) ;
and ( 
    .Z ( U755.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_35 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U755.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_35 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U755.EF ) ,
    .I0 ( xor_decoded_masks_0_35 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_35 ) ,
    .I0 ( U755.AB ) ,
    .I1 ( U755.CD ) ,
    .I2 ( U755.EF ) ) ;
and ( 
    .Z ( U1005.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_36 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1005.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_36 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1005.EF ) ,
    .I0 ( xor_decoded_masks_7_36 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_36 ) ,
    .I0 ( U1005.AB ) ,
    .I1 ( U1005.CD ) ,
    .I2 ( U1005.EF ) ) ;
and ( 
    .Z ( U439.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_55 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U439.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_2 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U439.EF ) ,
    .I0 ( xor_decoded_masks_6_2 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_2 ) ,
    .I0 ( U439.AB ) ,
    .I1 ( U439.CD ) ,
    .I2 ( U439.EF ) ) ;
and ( 
    .Z ( U754.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_65 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U754.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_11 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U754.EF ) ,
    .I0 ( xor_decoded_masks_1_11 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_11 ) ,
    .I0 ( U754.AB ) ,
    .I1 ( U754.CD ) ,
    .I2 ( U754.EF ) ) ;
and ( 
    .Z ( U1006.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_20 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1006.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_20 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1006.EF ) ,
    .I0 ( xor_decoded_masks_7_20 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_20 ) ,
    .I0 ( U1006.AB ) ,
    .I1 ( U1006.CD ) ,
    .I2 ( U1006.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_3_4 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_3.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_3.CD ) ,
    .IN ( masks_shift_reg_3_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_3 ) ) ;
and ( 
    .Z ( U753.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_75 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U753.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_21 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U753.EF ) ,
    .I0 ( xor_decoded_masks_1_21 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_21 ) ,
    .I0 ( U753.AB ) ,
    .I1 ( U753.CD ) ,
    .I2 ( U753.EF ) ) ;
and ( 
    .Z ( U1007.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_14 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1007.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_14 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1007.EF ) ,
    .I0 ( xor_decoded_masks_7_14 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_14 ) ,
    .I0 ( U1007.AB ) ,
    .I1 ( U1007.CD ) ,
    .I2 ( U1007.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_3_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_2.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_2.CD ) ,
    .IN ( masks_shift_reg_3_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_2 ) ) ;
and ( 
    .Z ( U752.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_69 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U752.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_15 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U752.EF ) ,
    .I0 ( xor_decoded_masks_1_15 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_15 ) ,
    .I0 ( U752.AB ) ,
    .I1 ( U752.CD ) ,
    .I2 ( U752.EF ) ) ;
and ( 
    .Z ( U1000.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_20 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1000.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_20 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1000.EF ) ,
    .I0 ( xor_decoded_masks_5_20 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_20 ) ,
    .I0 ( U1000.AB ) ,
    .I1 ( U1000.CD ) ,
    .I2 ( U1000.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_3_2 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_1.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_1.CD ) ,
    .IN ( masks_shift_reg_3_reg_1.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_1.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_1.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_1.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_1.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_1.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_1.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_1.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_1.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_1.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_1.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_1.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_1.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_1 ) ) ;
and ( 
    .Z ( U751.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_71 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U751.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_17 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U751.EF ) ,
    .I0 ( xor_decoded_masks_1_17 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_17 ) ,
    .I0 ( U751.AB ) ,
    .I1 ( U751.CD ) ,
    .I2 ( U751.EF ) ) ;
and ( 
    .Z ( U1001.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_14 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1001.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_14 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1001.EF ) ,
    .I0 ( xor_decoded_masks_5_14 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_14 ) ,
    .I0 ( U1001.AB ) ,
    .I1 ( U1001.CD ) ,
    .I2 ( U1001.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_3_1 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_0.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_0.CD ) ,
    .IN ( masks_shift_reg_3_reg_0.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_0.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_0.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_0.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_0.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_0.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_0.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_0.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_0.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_0.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_0.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_0.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_0.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_0 ) ) ;
and ( 
    .Z ( U750.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_91 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U750.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_37 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U750.EF ) ,
    .I0 ( xor_decoded_masks_1_37 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_37 ) ,
    .I0 ( U750.AB ) ,
    .I1 ( U750.CD ) ,
    .I2 ( U750.EF ) ) ;
and ( 
    .Z ( U1002.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_10 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1002.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_10 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1002.EF ) ,
    .I0 ( xor_decoded_masks_5_10 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_10 ) ,
    .I0 ( U1002.AB ) ,
    .I1 ( U1002.CD ) ,
    .I2 ( U1002.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_3_8 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_7.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_7.CD ) ,
    .IN ( masks_shift_reg_3_reg_7.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_7.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_7.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_7.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_7.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_7.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_7.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_7.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_7.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_7.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_7.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_7.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_7.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_7 ) ) ;
and ( 
    .Z ( U1003.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_24 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1003.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_24 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1003.EF ) ,
    .I0 ( xor_decoded_masks_7_24 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_24 ) ,
    .I0 ( U1003.AB ) ,
    .I1 ( U1003.CD ) ,
    .I2 ( U1003.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_3_7 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_6.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_6.CD ) ,
    .IN ( masks_shift_reg_3_reg_6.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_6.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_6.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_6.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_6.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_6.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_6.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_6.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_6.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_6.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_6.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_6.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_6.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_3_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_5.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_5.CD ) ,
    .IN ( masks_shift_reg_3_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_5 ) ) ;
and ( 
    .Z ( U674.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_65 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U674.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_12 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U674.EF ) ,
    .I0 ( xor_decoded_masks_4_12 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_12 ) ,
    .I0 ( U674.AB ) ,
    .I1 ( U674.CD ) ,
    .I2 ( U674.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_3_5 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2961 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_3_reg_4.CDNI_ ) ,
    .IN ( n48 ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_4.CD ) ,
    .IN ( masks_shift_reg_3_reg_4.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_3_reg_4.U5.CD_ ) ,
    .IN ( masks_shift_reg_3_reg_4.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_3_reg_4.U5.D_1 ) ,
    .I0 ( masks_shift_reg_3_reg_4.DI_ ) ,
    .I1 ( masks_shift_reg_3_reg_4.U5.CD_ ) ) ;
MUX21 masks_shift_reg_3_reg_4.U5.I2 ( 
    .I0 ( masks_shift_reg_3_reg_4.U5.D_1 ) ,
    .I1 ( masks_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_3_reg_4.U5.Q1 ) ,
    .S ( masks_shift_reg_3_reg_4.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_3_reg_4.U5.I3 ( 
    .CK ( masks_shift_reg_3_reg_4.CPI_ ) ,
    .D ( masks_shift_reg_3_reg_4.U5.Q1 ) ,
    .Q ( masks_shift_reg_3_4 ) ) ;
and ( 
    .Z ( U675.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_87 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U675.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_34 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U675.EF ) ,
    .I0 ( xor_decoded_masks_6_34 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_34 ) ,
    .I0 ( U675.AB ) ,
    .I1 ( U675.CD ) ,
    .I2 ( U675.EF ) ) ;
and ( 
    .Z ( U1127.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_15 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1127.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_15 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1127.EF ) ,
    .I0 ( xor_decoded_masks_5_15 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_15 ) ,
    .I0 ( U1127.AB ) ,
    .I1 ( U1127.CD ) ,
    .I2 ( U1127.EF ) ) ;
and ( 
    .Z ( U676.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_79 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U676.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_26 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U676.EF ) ,
    .I0 ( xor_decoded_masks_6_26 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_26 ) ,
    .I0 ( U676.AB ) ,
    .I1 ( U676.CD ) ,
    .I2 ( U676.EF ) ) ;
and ( 
    .Z ( U1126.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_21 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1126.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_21 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1126.EF ) ,
    .I0 ( xor_decoded_masks_5_21 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_21 ) ,
    .I0 ( U1126.AB ) ,
    .I1 ( U1126.CD ) ,
    .I2 ( U1126.EF ) ) ;
and ( 
    .Z ( U677.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_91 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U677.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_38 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U677.EF ) ,
    .I0 ( xor_decoded_masks_6_38 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_38 ) ,
    .I0 ( U677.AB ) ,
    .I1 ( U677.CD ) ,
    .I2 ( U677.EF ) ) ;
and ( 
    .Z ( U1125.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_17 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1125.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_17 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1125.EF ) ,
    .I0 ( xor_decoded_masks_5_17 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_17 ) ,
    .I0 ( U1125.AB ) ,
    .I1 ( U1125.CD ) ,
    .I2 ( U1125.EF ) ) ;
and ( 
    .Z ( U1008.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_10 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1008.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_10 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1008.EF ) ,
    .I0 ( xor_decoded_masks_7_10 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_10 ) ,
    .I0 ( U1008.AB ) ,
    .I1 ( U1008.CD ) ,
    .I2 ( U1008.EF ) ) ;
and ( 
    .Z ( U979.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_25 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U979.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_25 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U979.EF ) ,
    .I0 ( xor_decoded_masks_0_25 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_25 ) ,
    .I0 ( U979.AB ) ,
    .I1 ( U979.CD ) ,
    .I2 ( U979.EF ) ) ;
and ( 
    .Z ( U670.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_119 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U670.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_12 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U670.EF ) ,
    .I0 ( xor_decoded_masks_2_12 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_12 ) ,
    .I0 ( U670.AB ) ,
    .I1 ( U670.CD ) ,
    .I2 ( U670.EF ) ) ;
and ( 
    .Z ( U1124.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_37 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1124.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_37 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1124.EF ) ,
    .I0 ( xor_decoded_masks_5_37 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_37 ) ,
    .I0 ( U1124.AB ) ,
    .I1 ( U1124.CD ) ,
    .I2 ( U1124.EF ) ) ;
and ( 
    .Z ( U759.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_126 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U759.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_19 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U759.EF ) ,
    .I0 ( xor_decoded_masks_2_19 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_19 ) ,
    .I0 ( U759.AB ) ,
    .I1 ( U759.CD ) ,
    .I2 ( U759.EF ) ) ;
and ( 
    .Z ( U1009.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_24 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1009.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_24 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1009.EF ) ,
    .I0 ( xor_decoded_masks_9_24 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_24 ) ,
    .I0 ( U1009.AB ) ,
    .I1 ( U1009.CD ) ,
    .I2 ( U1009.EF ) ) ;
and ( 
    .Z ( U978.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_17 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U978.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_17 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U978.EF ) ,
    .I0 ( xor_decoded_masks_0_17 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_17 ) ,
    .I0 ( U978.AB ) ,
    .I1 ( U978.CD ) ,
    .I2 ( U978.EF ) ) ;
and ( 
    .Z ( U671.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_87 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U671.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_34 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U671.EF ) ,
    .I0 ( xor_decoded_masks_4_34 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_34 ) ,
    .I0 ( U671.AB ) ,
    .I1 ( U671.CD ) ,
    .I2 ( U671.EF ) ) ;
and ( 
    .Z ( U1123.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_33 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1123.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_33 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1123.EF ) ,
    .I0 ( xor_decoded_masks_5_33 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_33 ) ,
    .I0 ( U1123.AB ) ,
    .I1 ( U1123.CD ) ,
    .I2 ( U1123.EF ) ) ;
and ( 
    .Z ( U758.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_146 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U758.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_39 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U758.EF ) ,
    .I0 ( xor_decoded_masks_2_39 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_39 ) ,
    .I0 ( U758.AB ) ,
    .I1 ( U758.CD ) ,
    .I2 ( U758.EF ) ) ;
and ( 
    .Z ( U672.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_79 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U672.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_26 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U672.EF ) ,
    .I0 ( xor_decoded_masks_4_26 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_26 ) ,
    .I0 ( U672.AB ) ,
    .I1 ( U672.CD ) ,
    .I2 ( U672.EF ) ) ;
and ( 
    .Z ( U1122.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_25 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1122.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_25 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1122.EF ) ,
    .I0 ( xor_decoded_masks_5_25 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_25 ) ,
    .I0 ( U1122.AB ) ,
    .I1 ( U1122.CD ) ,
    .I2 ( U1122.EF ) ) ;
and ( 
    .Z ( U673.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_91 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U673.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_38 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U673.EF ) ,
    .I0 ( xor_decoded_masks_4_38 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_38 ) ,
    .I0 ( U673.AB ) ,
    .I1 ( U673.CD ) ,
    .I2 ( U673.EF ) ) ;
and ( 
    .Z ( U1121.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_29 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1121.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_29 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1121.EF ) ,
    .I0 ( xor_decoded_masks_5_29 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_29 ) ,
    .I0 ( U1121.AB ) ,
    .I1 ( U1121.CD ) ,
    .I2 ( U1121.EF ) ) ;
and ( 
    .Z ( U1120.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_11 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1120.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_11 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1120.EF ) ,
    .I0 ( xor_decoded_masks_3_11 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_11 ) ,
    .I0 ( U1120.AB ) ,
    .I1 ( U1120.CD ) ,
    .I2 ( U1120.EF ) ) ;
or ( 
    .Z ( U973.AB ) ,
    .I0 ( n7 ) ,
    .I1 ( n18 ) ) ;
not ( 
    .O1 ( U973.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_9 ) ) ;
not ( 
    .O1 ( U973.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U973.not_c_tempD ) ,
    .I0 ( U973.not_c_temp ) ,
    .I1 ( U973.ND ) ) ;
and ( 
    .Z ( U973.ZN ) ,
    .I0 ( U973.AB ) ,
    .I1 ( U973.not_c_tempD ) ) ;
not ( 
    .O1 ( N201 ) ,
    .IN ( U973.ZN ) ) ;
or ( 
    .Z ( U972.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_5 ) ) ;
not ( 
    .O1 ( U972.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_10 ) ) ;
not ( 
    .O1 ( U972.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U972.not_c_tempD ) ,
    .I0 ( U972.not_c_temp ) ,
    .I1 ( U972.ND ) ) ;
and ( 
    .Z ( U972.ZN ) ,
    .I0 ( U972.AB ) ,
    .I1 ( U972.not_c_tempD ) ) ;
not ( 
    .O1 ( N212 ) ,
    .IN ( U972.ZN ) ) ;
and ( 
    .Z ( U971.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_54 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U971.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_1 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U971.EF ) ,
    .I0 ( xor_decoded_masks_14_1 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_1 ) ,
    .I0 ( U971.AB ) ,
    .I1 ( U971.CD ) ,
    .I2 ( U971.EF ) ) ;
and ( 
    .Z ( U678.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_61 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U678.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_8 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U678.EF ) ,
    .I0 ( xor_decoded_masks_6_8 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_8 ) ,
    .I0 ( U678.AB ) ,
    .I1 ( U678.CD ) ,
    .I2 ( U678.EF ) ) ;
or ( 
    .Z ( U970.AB ) ,
    .I0 ( n15 ) ,
    .I1 ( n18 ) ) ;
not ( 
    .O1 ( U970.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_11 ) ) ;
not ( 
    .O1 ( U970.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U970.not_c_tempD ) ,
    .I0 ( U970.not_c_temp ) ,
    .I1 ( U970.ND ) ) ;
and ( 
    .Z ( U970.ZN ) ,
    .I0 ( U970.AB ) ,
    .I1 ( U970.not_c_tempD ) ) ;
not ( 
    .O1 ( N223 ) ,
    .IN ( U970.ZN ) ) ;
and ( 
    .Z ( U679.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_65 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U679.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_12 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U679.EF ) ,
    .I0 ( xor_decoded_masks_6_12 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_12 ) ,
    .I0 ( U679.AB ) ,
    .I1 ( U679.CD ) ,
    .I2 ( U679.EF ) ) ;
or ( 
    .Z ( U977.AB ) ,
    .I0 ( n9 ) ,
    .I1 ( n18 ) ) ;
not ( 
    .O1 ( U977.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_7 ) ) ;
not ( 
    .O1 ( U977.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U977.not_c_tempD ) ,
    .I0 ( U977.not_c_temp ) ,
    .I1 ( U977.ND ) ) ;
and ( 
    .Z ( U977.ZN ) ,
    .I0 ( U977.AB ) ,
    .I1 ( U977.not_c_tempD ) ) ;
not ( 
    .O1 ( N179 ) ,
    .IN ( U977.ZN ) ) ;
and ( 
    .Z ( U401.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_19 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U401.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_19 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U401.EF ) ,
    .I0 ( xor_decoded_masks_11_19 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_19 ) ,
    .I0 ( U401.AB ) ,
    .I1 ( U401.CD ) ,
    .I2 ( U401.EF ) ) ;
or ( 
    .Z ( U976.AB ) ,
    .I0 ( n18 ) ,
    .I1 ( edt_channels_out_from_constant_shift_control_4 ) ) ;
not ( 
    .O1 ( U976.not_c_temp ) ,
    .IN ( edt_channels_out_from_constant_shift_control_8 ) ) ;
not ( 
    .O1 ( U976.ND ) ,
    .IN ( n20 ) ) ;
or ( 
    .Z ( U976.not_c_tempD ) ,
    .I0 ( U976.not_c_temp ) ,
    .I1 ( U976.ND ) ) ;
and ( 
    .Z ( U976.ZN ) ,
    .I0 ( U976.AB ) ,
    .I1 ( U976.not_c_tempD ) ) ;
not ( 
    .O1 ( N190 ) ,
    .IN ( U976.ZN ) ) ;
and ( 
    .Z ( U1129.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_29 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1129.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_29 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1129.EF ) ,
    .I0 ( xor_decoded_masks_7_29 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_29 ) ,
    .I0 ( U1129.AB ) ,
    .I1 ( U1129.CD ) ,
    .I2 ( U1129.EF ) ) ;
and ( 
    .Z ( U400.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_18 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U400.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_18 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U400.EF ) ,
    .I0 ( xor_decoded_masks_11_18 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_18 ) ,
    .I0 ( U400.AB ) ,
    .I1 ( U400.CD ) ,
    .I2 ( U400.EF ) ) ;
and ( 
    .Z ( U506.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_48 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U506.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_48 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U506.EF ) ,
    .I0 ( xor_decoded_masks_5_48 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_48 ) ,
    .I0 ( U506.AB ) ,
    .I1 ( U506.CD ) ,
    .I2 ( U506.EF ) ) ;
and ( 
    .Z ( U1256.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_158 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1256.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_51 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1256.EF ) ,
    .I0 ( xor_decoded_masks_2_51 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_51 ) ,
    .I0 ( U1256.AB ) ,
    .I1 ( U1256.CD ) ,
    .I2 ( U1256.EF ) ) ;
and ( 
    .Z ( U507.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_101 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U507.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_48 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U507.EF ) ,
    .I0 ( xor_decoded_masks_6_48 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_48 ) ,
    .I0 ( U507.AB ) ,
    .I1 ( U507.CD ) ,
    .I2 ( U507.EF ) ) ;
and ( 
    .Z ( U1255.AB ) ,
    .I0 ( masks_hold_reg_8_5 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U1255.CD ) ,
    .I0 ( config1_xor_encoded_masks_92 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_92 ) ,
    .I0 ( U1255.AB ) ,
    .I1 ( U1255.CD ) ) ;
and ( 
    .Z ( U508.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_48 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U508.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_48 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U508.EF ) ,
    .I0 ( xor_decoded_masks_7_48 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_48 ) ,
    .I0 ( U508.AB ) ,
    .I1 ( U508.CD ) ,
    .I2 ( U508.EF ) ) ;
and ( 
    .Z ( U1254.AB ) ,
    .I0 ( masks_hold_reg_6_3 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U1254.CD ) ,
    .I0 ( config1_xor_encoded_masks_72 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_72 ) ,
    .I0 ( U1254.AB ) ,
    .I1 ( U1254.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_2_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_10.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_10 ) ,
    .IN ( masks_hold_reg_2_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_2_reg_10.QT ) ,
    .I1 ( masks_hold_reg_2_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_10.ED ) ,
    .S ( masks_hold_reg_2_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_10.ED ) ,
    .I1 ( masks_hold_reg_2_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_2_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_2_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_10.QT ) ) ;
and ( 
    .Z ( U509.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_101 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U509.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_48 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U509.EF ) ,
    .I0 ( xor_decoded_masks_8_48 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_48 ) ,
    .I0 ( U509.AB ) ,
    .I1 ( U509.CD ) ,
    .I2 ( U509.EF ) ) ;
and ( 
    .Z ( U423.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_58 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U423.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_5 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U423.EF ) ,
    .I0 ( xor_decoded_masks_4_5 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_5 ) ,
    .I0 ( U423.AB ) ,
    .I1 ( U423.CD ) ,
    .I2 ( U423.EF ) ) ;
and ( 
    .Z ( U422.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_2 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U422.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_2 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U422.EF ) ,
    .I0 ( xor_decoded_masks_3_2 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_2 ) ,
    .I0 ( U422.AB ) ,
    .I1 ( U422.CD ) ,
    .I2 ( U422.EF ) ) ;
and ( 
    .Z ( U1259.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_51 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1259.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_51 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1259.EF ) ,
    .I0 ( xor_decoded_masks_5_51 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_51 ) ,
    .I0 ( U1259.AB ) ,
    .I1 ( U1259.CD ) ,
    .I2 ( U1259.EF ) ) ;
and ( 
    .Z ( U421.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_3 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U421.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_3 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U421.EF ) ,
    .I0 ( xor_decoded_masks_3_3 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_3 ) ,
    .I0 ( U421.AB ) ,
    .I1 ( U421.CD ) ,
    .I2 ( U421.EF ) ) ;
and ( 
    .Z ( U1258.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_104 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1258.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_51 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1258.EF ) ,
    .I0 ( xor_decoded_masks_4_51 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_51 ) ,
    .I0 ( U1258.AB ) ,
    .I1 ( U1258.CD ) ,
    .I2 ( U1258.EF ) ) ;
and ( 
    .Z ( U420.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_0 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U420.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_0 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U420.EF ) ,
    .I0 ( xor_decoded_masks_3_0 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_0 ) ,
    .I0 ( U420.AB ) ,
    .I1 ( U420.CD ) ,
    .I2 ( U420.EF ) ) ;
and ( 
    .Z ( U427.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_56 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U427.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_3 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U427.EF ) ,
    .I0 ( xor_decoded_masks_4_3 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_3 ) ,
    .I0 ( U427.AB ) ,
    .I1 ( U427.CD ) ,
    .I2 ( U427.EF ) ) ;
and ( 
    .Z ( U426.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_53 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U426.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_0 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U426.EF ) ,
    .I0 ( xor_decoded_masks_4_0 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_0 ) ,
    .I0 ( U426.AB ) ,
    .I1 ( U426.CD ) ,
    .I2 ( U426.EF ) ) ;
and ( 
    .Z ( U425.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_59 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U425.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_6 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U425.EF ) ,
    .I0 ( xor_decoded_masks_4_6 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_6 ) ,
    .I0 ( U425.AB ) ,
    .I1 ( U425.CD ) ,
    .I2 ( U425.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_10.DI_ ) ,
    .IN ( N234 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_12_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
DFF masks_shift_reg_12_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_12_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_12_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_12_10 ) ) ;
and ( 
    .Z ( U424.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_60 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U424.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_7 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U424.EF ) ,
    .I0 ( xor_decoded_masks_4_7 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_7 ) ,
    .I0 ( U424.AB ) ,
    .I1 ( U424.CD ) ,
    .I2 ( U424.EF ) ) ;
and ( 
    .Z ( U746.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_74 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U746.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_21 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U746.EF ) ,
    .I0 ( xor_decoded_masks_14_21 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_21 ) ,
    .I0 ( U746.AB ) ,
    .I1 ( U746.CD ) ,
    .I2 ( U746.EF ) ) ;
and ( 
    .Z ( U747.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_83 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U747.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_29 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U747.EF ) ,
    .I0 ( xor_decoded_masks_1_29 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_29 ) ,
    .I0 ( U747.AB ) ,
    .I1 ( U747.CD ) ,
    .I2 ( U747.EF ) ) ;
and ( 
    .Z ( U1128.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_11 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1128.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_11 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1128.EF ) ,
    .I0 ( xor_decoded_masks_5_11 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_11 ) ,
    .I0 ( U1128.AB ) ,
    .I1 ( U1128.CD ) ,
    .I2 ( U1128.EF ) ) ;
and ( 
    .Z ( U403.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_75 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U403.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_22 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U403.EF ) ,
    .I0 ( xor_decoded_masks_12_22 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_22 ) ,
    .I0 ( U403.AB ) ,
    .I1 ( U403.CD ) ,
    .I2 ( U403.EF ) ) ;
and ( 
    .Z ( U974.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_99 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U974.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_45 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U974.EF ) ,
    .I0 ( xor_decoded_masks_1_45 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_45 ) ,
    .I0 ( U974.AB ) ,
    .I1 ( U974.CD ) ,
    .I2 ( U974.EF ) ) ;
and ( 
    .Z ( U402.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_83 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U402.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_30 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U402.EF ) ,
    .I0 ( xor_decoded_masks_12_30 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_30 ) ,
    .I0 ( U402.AB ) ,
    .I1 ( U402.CD ) ,
    .I2 ( U402.EF ) ) ;
and ( 
    .Z ( U405.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_28 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U405.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_28 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U405.EF ) ,
    .I0 ( xor_decoded_masks_13_28 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_28 ) ,
    .I0 ( U405.AB ) ,
    .I1 ( U405.CD ) ,
    .I2 ( U405.EF ) ) ;
and ( 
    .Z ( U404.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_76 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U404.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_23 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U404.EF ) ,
    .I0 ( xor_decoded_masks_12_23 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_23 ) ,
    .I0 ( U404.AB ) ,
    .I1 ( U404.CD ) ,
    .I2 ( U404.EF ) ) ;
and ( 
    .Z ( U407.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_31 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U407.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_31 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U407.EF ) ,
    .I0 ( xor_decoded_masks_13_31 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_31 ) ,
    .I0 ( U407.AB ) ,
    .I1 ( U407.CD ) ,
    .I2 ( U407.EF ) ) ;
and ( 
    .Z ( U406.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_30 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U406.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_30 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U406.EF ) ,
    .I0 ( xor_decoded_masks_13_30 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_30 ) ,
    .I0 ( U406.AB ) ,
    .I1 ( U406.CD ) ,
    .I2 ( U406.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_5_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29282 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_5_10 ) ,
    .IN ( masks_hold_reg_5_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_27 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_28 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_29 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_5_reg_10.SYNTEST_VL_LSI_MUX21_26786.I0 ( 
    .I0 ( masks_hold_reg_5_reg_10.QT ) ,
    .I1 ( masks_hold_reg_5_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_5_reg_10.ED ) ,
    .S ( masks_hold_reg_5_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_5_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_29 ) ) ;
and ( 
    .Z ( masks_hold_reg_5_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_5_reg_10.ED ) ,
    .I1 ( masks_hold_reg_5_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_5_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_5_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_27 ) ,
    .Q ( masks_hold_reg_5_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_5_reg_10.SYNTEST_EXP_ADDED_NET_28 ) ) ;
DFF masks_hold_reg_5_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_5_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_5_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_5_reg_10.QT ) ) ;
and ( 
    .Z ( U409.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_19 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U409.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_19 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U409.EF ) ,
    .I0 ( xor_decoded_masks_13_19 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_19 ) ,
    .I0 ( U409.AB ) ,
    .I1 ( U409.CD ) ,
    .I2 ( U409.EF ) ) ;
and ( 
    .Z ( U408.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_18 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U408.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_18 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U408.EF ) ,
    .I0 ( xor_decoded_masks_13_18 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_18 ) ,
    .I0 ( U408.AB ) ,
    .I1 ( U408.CD ) ,
    .I2 ( U408.EF ) ) ;
and ( 
    .Z ( U720.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_78 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U720.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_25 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U720.EF ) ,
    .I0 ( xor_decoded_masks_6_25 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_25 ) ,
    .I0 ( U720.AB ) ,
    .I1 ( U720.CD ) ,
    .I2 ( U720.EF ) ) ;
and ( 
    .Z ( U1073.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_22 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1073.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_22 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1073.EF ) ,
    .I0 ( xor_decoded_masks_9_22 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_22 ) ,
    .I0 ( U1073.AB ) ,
    .I1 ( U1073.CD ) ,
    .I2 ( U1073.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_11_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_7.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_7 ) ,
    .IN ( masks_hold_reg_11_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_7.QT ) ,
    .I1 ( masks_hold_reg_11_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_7.ED ) ,
    .S ( masks_hold_reg_11_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_7.ED ) ,
    .I1 ( masks_hold_reg_11_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_7.QT ) ) ;
and ( 
    .Z ( U721.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_90 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U721.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_37 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U721.EF ) ,
    .I0 ( xor_decoded_masks_6_37 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_37 ) ,
    .I0 ( U721.AB ) ,
    .I1 ( U721.CD ) ,
    .I2 ( U721.EF ) ) ;
and ( 
    .Z ( U1072.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_38 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1072.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_38 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1072.EF ) ,
    .I0 ( xor_decoded_masks_9_38 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_38 ) ,
    .I0 ( U1072.AB ) ,
    .I1 ( U1072.CD ) ,
    .I2 ( U1072.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_11_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_6.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_6 ) ,
    .IN ( masks_hold_reg_11_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_6.QT ) ,
    .I1 ( masks_hold_reg_11_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_6.ED ) ,
    .S ( masks_hold_reg_11_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_6.ED ) ,
    .I1 ( masks_hold_reg_11_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_6.QT ) ) ;
and ( 
    .Z ( U722.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_74 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U722.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_21 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U722.EF ) ,
    .I0 ( xor_decoded_masks_6_21 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_21 ) ,
    .I0 ( U722.AB ) ,
    .I1 ( U722.CD ) ,
    .I2 ( U722.EF ) ) ;
and ( 
    .Z ( U1071.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_34 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1071.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_34 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1071.EF ) ,
    .I0 ( xor_decoded_masks_9_34 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_34 ) ,
    .I0 ( U1071.AB ) ,
    .I1 ( U1071.CD ) ,
    .I2 ( U1071.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_11_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_5.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_5 ) ,
    .IN ( masks_hold_reg_11_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_5.QT ) ,
    .I1 ( masks_hold_reg_11_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_5.ED ) ,
    .S ( masks_hold_reg_11_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_5.ED ) ,
    .I1 ( masks_hold_reg_11_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_5.QT ) ) ;
and ( 
    .Z ( U723.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_68 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U723.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_15 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U723.EF ) ,
    .I0 ( xor_decoded_masks_6_15 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_15 ) ,
    .I0 ( U723.AB ) ,
    .I1 ( U723.CD ) ,
    .I2 ( U723.EF ) ) ;
and ( 
    .Z ( U1070.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_26 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1070.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_26 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1070.EF ) ,
    .I0 ( xor_decoded_masks_9_26 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_26 ) ,
    .I0 ( U1070.AB ) ,
    .I1 ( U1070.CD ) ,
    .I2 ( U1070.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_11_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_4.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_4.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_4 ) ,
    .IN ( masks_hold_reg_11_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_4.QT ) ,
    .I1 ( masks_hold_reg_11_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_4.ED ) ,
    .S ( masks_hold_reg_11_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_4.ED ) ,
    .I1 ( masks_hold_reg_11_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_4.QT ) ) ;
and ( 
    .Z ( U724.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_64 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U724.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_11 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U724.EF ) ,
    .I0 ( xor_decoded_masks_6_11 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_11 ) ,
    .I0 ( U724.AB ) ,
    .I1 ( U724.CD ) ,
    .I2 ( U724.EF ) ) ;
and ( 
    .Z ( U1077.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_61 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1077.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_8 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1077.EF ) ,
    .I0 ( xor_decoded_masks_10_8 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_8 ) ,
    .I0 ( U1077.AB ) ,
    .I1 ( U1077.CD ) ,
    .I2 ( U1077.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_11_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_3.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_3 ) ,
    .IN ( masks_hold_reg_11_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_3.QT ) ,
    .I1 ( masks_hold_reg_11_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_3.ED ) ,
    .S ( masks_hold_reg_11_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_3.ED ) ,
    .I1 ( masks_hold_reg_11_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_3.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_1_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_10.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_10 ) ,
    .IN ( masks_hold_reg_1_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_10.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_10.QT ) ,
    .I1 ( masks_hold_reg_1_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_10.ED ) ,
    .S ( masks_hold_reg_1_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_10.ED ) ,
    .I1 ( masks_hold_reg_1_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_10.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_10.QT ) ) ;
and ( 
    .Z ( U725.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_70 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U725.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_17 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U725.EF ) ,
    .I0 ( xor_decoded_masks_6_17 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_17 ) ,
    .I0 ( U725.AB ) ,
    .I1 ( U725.CD ) ,
    .I2 ( U725.EF ) ) ;
and ( 
    .Z ( U1076.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_79 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1076.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_26 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1076.EF ) ,
    .I0 ( xor_decoded_masks_10_26 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_26 ) ,
    .I0 ( U1076.AB ) ,
    .I1 ( U1076.CD ) ,
    .I2 ( U1076.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_10.DI_ ) ,
    .IN ( N223 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_11_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_3_1 ) ) ;
DFF masks_shift_reg_11_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_11_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_11_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_11_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_11_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_2.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_2 ) ,
    .IN ( masks_hold_reg_11_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_2.QT ) ,
    .I1 ( masks_hold_reg_11_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_2.ED ) ,
    .S ( masks_hold_reg_11_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_2.ED ) ,
    .I1 ( masks_hold_reg_11_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_2.QT ) ) ;
and ( 
    .Z ( U726.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_82 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U726.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_29 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U726.EF ) ,
    .I0 ( xor_decoded_masks_8_29 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_29 ) ,
    .I0 ( U726.AB ) ,
    .I1 ( U726.CD ) ,
    .I2 ( U726.EF ) ) ;
and ( 
    .Z ( U1075.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_12 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1075.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_12 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1075.EF ) ,
    .I0 ( xor_decoded_masks_9_12 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_12 ) ,
    .I0 ( U1075.AB ) ,
    .I1 ( U1075.CD ) ,
    .I2 ( U1075.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_11_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_1.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_1.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_1 ) ,
    .IN ( masks_hold_reg_11_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_1.QT ) ,
    .I1 ( masks_hold_reg_11_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_1.ED ) ,
    .S ( masks_hold_reg_11_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_1.ED ) ,
    .I1 ( masks_hold_reg_11_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_1.QT ) ) ;
and ( 
    .Z ( U727.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_86 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U727.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_33 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U727.EF ) ,
    .I0 ( xor_decoded_masks_8_33 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_33 ) ,
    .I0 ( U727.AB ) ,
    .I1 ( U727.CD ) ,
    .I2 ( U727.EF ) ) ;
and ( 
    .Z ( U1074.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_8 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1074.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_8 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1074.EF ) ,
    .I0 ( xor_decoded_masks_9_8 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_8 ) ,
    .I0 ( U1074.AB ) ,
    .I1 ( U1074.CD ) ,
    .I2 ( U1074.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_11_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_0.CPI_ ) ,
    .IN ( edt_clock_cts_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_0.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_0 ) ,
    .IN ( masks_hold_reg_11_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_0.QT ) ,
    .I1 ( masks_hold_reg_11_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_0.ED ) ,
    .S ( masks_hold_reg_11_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_0.ED ) ,
    .I1 ( masks_hold_reg_11_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_0.QT ) ) ;
and ( 
    .Z ( U728.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_78 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U728.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_25 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U728.EF ) ,
    .I0 ( xor_decoded_masks_8_25 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_25 ) ,
    .I0 ( U728.AB ) ,
    .I1 ( U728.CD ) ,
    .I2 ( U728.EF ) ) ;
and ( 
    .Z ( U647.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_63 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U647.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_10 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U647.EF ) ,
    .I0 ( xor_decoded_masks_6_10 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_10 ) ,
    .I0 ( U647.AB ) ,
    .I1 ( U647.CD ) ,
    .I2 ( U647.EF ) ) ;
and ( 
    .Z ( U729.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_90 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U729.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_37 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U729.EF ) ,
    .I0 ( xor_decoded_masks_8_37 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_37 ) ,
    .I0 ( U729.AB ) ,
    .I1 ( U729.CD ) ,
    .I2 ( U729.EF ) ) ;
and ( 
    .Z ( U646.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_67 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U646.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_14 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U646.EF ) ,
    .I0 ( xor_decoded_masks_6_14 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_14 ) ,
    .I0 ( U646.AB ) ,
    .I1 ( U646.CD ) ,
    .I2 ( U646.EF ) ) ;
and ( 
    .Z ( U1114.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_25 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1114.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_25 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1114.EF ) ,
    .I0 ( xor_decoded_masks_3_25 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_25 ) ,
    .I0 ( U1114.AB ) ,
    .I1 ( U1114.CD ) ,
    .I2 ( U1114.EF ) ) ;
and ( 
    .Z ( U1079.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_71 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1079.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_18 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1079.EF ) ,
    .I0 ( xor_decoded_masks_10_18 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_18 ) ,
    .I0 ( U1079.AB ) ,
    .I1 ( U1079.CD ) ,
    .I2 ( U1079.EF ) ) ;
and ( 
    .Z ( U948.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_1 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U948.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_1 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U948.EF ) ,
    .I0 ( xor_decoded_masks_5_1 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_1 ) ,
    .I0 ( U948.AB ) ,
    .I1 ( U948.CD ) ,
    .I2 ( U948.EF ) ) ;
and ( 
    .Z ( U645.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_89 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U645.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_36 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U645.EF ) ,
    .I0 ( xor_decoded_masks_6_36 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_36 ) ,
    .I0 ( U645.AB ) ,
    .I1 ( U645.CD ) ,
    .I2 ( U645.EF ) ) ;
and ( 
    .Z ( U1115.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_29 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1115.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_29 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1115.EF ) ,
    .I0 ( xor_decoded_masks_3_29 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_29 ) ,
    .I0 ( U1115.AB ) ,
    .I1 ( U1115.CD ) ,
    .I2 ( U1115.EF ) ) ;
and ( 
    .Z ( U1078.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_65 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1078.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_12 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1078.EF ) ,
    .I0 ( xor_decoded_masks_10_12 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_12 ) ,
    .I0 ( U1078.AB ) ,
    .I1 ( U1078.CD ) ,
    .I2 ( U1078.EF ) ) ;
and ( 
    .Z ( U949.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_98 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U949.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_45 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U949.EF ) ,
    .I0 ( xor_decoded_masks_6_45 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_45 ) ,
    .I0 ( U949.AB ) ,
    .I1 ( U949.CD ) ,
    .I2 ( U949.EF ) ) ;
and ( 
    .Z ( U644.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_77 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U644.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_24 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U644.EF ) ,
    .I0 ( xor_decoded_masks_6_24 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_24 ) ,
    .I0 ( U644.AB ) ,
    .I1 ( U644.CD ) ,
    .I2 ( U644.EF ) ) ;
and ( 
    .Z ( U1116.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_37 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1116.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_37 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1116.EF ) ,
    .I0 ( xor_decoded_masks_3_37 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_37 ) ,
    .I0 ( U1116.AB ) ,
    .I1 ( U1116.CD ) ,
    .I2 ( U1116.EF ) ) ;
and ( 
    .Z ( U643.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_85 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U643.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_32 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U643.EF ) ,
    .I0 ( xor_decoded_masks_6_32 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_32 ) ,
    .I0 ( U643.AB ) ,
    .I1 ( U643.CD ) ,
    .I2 ( U643.EF ) ) ;
and ( 
    .Z ( U1117.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_21 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1117.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_21 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1117.EF ) ,
    .I0 ( xor_decoded_masks_3_21 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_21 ) ,
    .I0 ( U1117.AB ) ,
    .I1 ( U1117.CD ) ,
    .I2 ( U1117.EF ) ) ;
and ( 
    .Z ( U642.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_67 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U642.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_14 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U642.EF ) ,
    .I0 ( xor_decoded_masks_4_14 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_14 ) ,
    .I0 ( U642.AB ) ,
    .I1 ( U642.CD ) ,
    .I2 ( U642.EF ) ) ;
and ( 
    .Z ( U1110.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_42 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1110.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_42 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1110.EF ) ,
    .I0 ( xor_decoded_masks_13_42 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_42 ) ,
    .I0 ( U1110.AB ) ,
    .I1 ( U1110.CD ) ,
    .I2 ( U1110.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_11_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_4_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_9.E_ ) ,
    .IN ( edt_update_hfs_netlink_29288 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_9 ) ,
    .IN ( masks_hold_reg_11_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_9.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_11_reg_9.QT ) ,
    .I1 ( masks_hold_reg_11_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_9.ED ) ,
    .S ( masks_hold_reg_11_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_9.ED ) ,
    .I1 ( masks_hold_reg_11_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_11_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_9.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_11_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_9.QT ) ) ;
and ( 
    .Z ( U641.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_89 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U641.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_36 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U641.EF ) ,
    .I0 ( xor_decoded_masks_4_36 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_36 ) ,
    .I0 ( U641.AB ) ,
    .I1 ( U641.CD ) ,
    .I2 ( U641.EF ) ) ;
and ( 
    .Z ( U1111.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_95 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1111.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_42 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1111.EF ) ,
    .I0 ( xor_decoded_masks_14_42 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_42 ) ,
    .I0 ( U1111.AB ) ,
    .I1 ( U1111.CD ) ,
    .I2 ( U1111.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_11_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_8.E_ ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_8 ) ,
    .IN ( masks_hold_reg_11_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_11_reg_8.QT ) ,
    .I1 ( masks_hold_reg_11_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_8.ED ) ,
    .S ( masks_hold_reg_11_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_8.ED ) ,
    .I1 ( masks_hold_reg_11_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_11_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_11_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_8.QT ) ) ;
and ( 
    .Z ( U640.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_77 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U640.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_24 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U640.EF ) ,
    .I0 ( xor_decoded_masks_4_24 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_24 ) ,
    .I0 ( U640.AB ) ,
    .I1 ( U640.CD ) ,
    .I2 ( U640.EF ) ) ;
and ( 
    .Z ( U1112.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_96 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1112.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_42 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1112.EF ) ,
    .I0 ( xor_decoded_masks_1_42 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_42 ) ,
    .I0 ( U1112.AB ) ,
    .I1 ( U1112.CD ) ,
    .I2 ( U1112.EF ) ) ;
and ( 
    .Z ( U1113.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_52 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1113.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_52 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1113.EF ) ,
    .I0 ( xor_decoded_masks_0_52 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_52 ) ,
    .I0 ( U1113.AB ) ,
    .I1 ( U1113.CD ) ,
    .I2 ( U1113.EF ) ) ;
and ( 
    .Z ( U940.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_152 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U940.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_45 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U940.EF ) ,
    .I0 ( xor_decoded_masks_2_45 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_45 ) ,
    .I0 ( U940.AB ) ,
    .I1 ( U940.CD ) ,
    .I2 ( U940.EF ) ) ;
and ( 
    .Z ( U941.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_108 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U941.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_1 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U941.EF ) ,
    .I0 ( xor_decoded_masks_2_1 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_1 ) ,
    .I0 ( U941.AB ) ,
    .I1 ( U941.CD ) ,
    .I2 ( U941.EF ) ) ;
and ( 
    .Z ( U942.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_45 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U942.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_45 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U942.EF ) ,
    .I0 ( xor_decoded_masks_3_45 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_45 ) ,
    .I0 ( U942.AB ) ,
    .I1 ( U942.CD ) ,
    .I2 ( U942.EF ) ) ;
and ( 
    .Z ( U943.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_5 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U943.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_5 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U943.EF ) ,
    .I0 ( xor_decoded_masks_3_5 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_5 ) ,
    .I0 ( U943.AB ) ,
    .I1 ( U943.CD ) ,
    .I2 ( U943.EF ) ) ;
and ( 
    .Z ( U1118.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_15 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1118.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_15 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1118.EF ) ,
    .I0 ( xor_decoded_masks_3_15 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_15 ) ,
    .I0 ( U1118.AB ) ,
    .I1 ( U1118.CD ) ,
    .I2 ( U1118.EF ) ) ;
and ( 
    .Z ( U869.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_104 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U869.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_51 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U869.EF ) ,
    .I0 ( xor_decoded_masks_12_51 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_51 ) ,
    .I0 ( U869.AB ) ,
    .I1 ( U869.CD ) ,
    .I2 ( U869.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_10.DI_ ) ,
    .IN ( N201 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_10.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
DFF masks_shift_reg_9_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_9_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_9_10 ) ) ;
and ( 
    .Z ( U944.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_98 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U944.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_45 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U944.EF ) ,
    .I0 ( xor_decoded_masks_4_45 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_45 ) ,
    .I0 ( U944.AB ) ,
    .I1 ( U944.CD ) ,
    .I2 ( U944.EF ) ) ;
and ( 
    .Z ( U649.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_77 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U649.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_24 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U649.EF ) ,
    .I0 ( xor_decoded_masks_8_24 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_24 ) ,
    .I0 ( U649.AB ) ,
    .I1 ( U649.CD ) ,
    .I2 ( U649.EF ) ) ;
and ( 
    .Z ( U1119.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_17 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1119.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_17 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1119.EF ) ,
    .I0 ( xor_decoded_masks_3_17 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_17 ) ,
    .I0 ( U1119.AB ) ,
    .I1 ( U1119.CD ) ,
    .I2 ( U1119.EF ) ) ;
and ( 
    .Z ( U410.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_75 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U410.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_22 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U410.EF ) ,
    .I0 ( xor_decoded_masks_14_22 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_22 ) ,
    .I0 ( U410.AB ) ,
    .I1 ( U410.CD ) ,
    .I2 ( U410.EF ) ) ;
and ( 
    .Z ( U868.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_51 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U868.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_51 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U868.EF ) ,
    .I0 ( xor_decoded_masks_11_51 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_51 ) ,
    .I0 ( U868.AB ) ,
    .I1 ( U868.CD ) ,
    .I2 ( U868.EF ) ) ;
and ( 
    .Z ( U945.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_54 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U945.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_1 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U945.EF ) ,
    .I0 ( xor_decoded_masks_4_1 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_1 ) ,
    .I0 ( U945.AB ) ,
    .I1 ( U945.CD ) ,
    .I2 ( U945.EF ) ) ;
and ( 
    .Z ( U648.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_69 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U648.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_16 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U648.EF ) ,
    .I0 ( xor_decoded_masks_6_16 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_16 ) ,
    .I0 ( U648.AB ) ,
    .I1 ( U648.CD ) ,
    .I2 ( U648.EF ) ) ;
and ( 
    .Z ( U411.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_76 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U411.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_23 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U411.EF ) ,
    .I0 ( xor_decoded_masks_14_23 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_23 ) ,
    .I0 ( U411.AB ) ,
    .I1 ( U411.CD ) ,
    .I2 ( U411.EF ) ) ;
and ( 
    .Z ( U946.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_45 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U946.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_45 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U946.EF ) ,
    .I0 ( xor_decoded_masks_5_45 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_45 ) ,
    .I0 ( U946.AB ) ,
    .I1 ( U946.CD ) ,
    .I2 ( U946.EF ) ) ;
and ( 
    .Z ( U412.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_114 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U412.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_7 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U412.EF ) ,
    .I0 ( xor_decoded_masks_2_7 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_7 ) ,
    .I0 ( U412.AB ) ,
    .I1 ( U412.CD ) ,
    .I2 ( U412.EF ) ) ;
and ( 
    .Z ( U947.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_5 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U947.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_5 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U947.EF ) ,
    .I0 ( xor_decoded_masks_5_5 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_5 ) ,
    .I0 ( U947.AB ) ,
    .I1 ( U947.CD ) ,
    .I2 ( U947.EF ) ) ;
and ( 
    .Z ( U413.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_113 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U413.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_6 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U413.EF ) ,
    .I0 ( xor_decoded_masks_2_6 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_6 ) ,
    .I0 ( U413.AB ) ,
    .I1 ( U413.CD ) ,
    .I2 ( U413.EF ) ) ;
and ( 
    .Z ( U414.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_107 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U414.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_0 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U414.EF ) ,
    .I0 ( xor_decoded_masks_2_0 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_0 ) ,
    .I0 ( U414.AB ) ,
    .I1 ( U414.CD ) ,
    .I2 ( U414.EF ) ) ;
and ( 
    .Z ( U415.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_110 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U415.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_3 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U415.EF ) ,
    .I0 ( xor_decoded_masks_2_3 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_3 ) ,
    .I0 ( U415.AB ) ,
    .I1 ( U415.CD ) ,
    .I2 ( U415.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_3.DI_ ) ,
    .IN ( n96 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_3.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_3.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_3.CD ) ,
    .IN ( masks_shift_reg_9_reg_3.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_3.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_3.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_3.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_3.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_3.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_3.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_3.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_3.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_3.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_3.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_3.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_3.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_3 ) ) ;
and ( 
    .Z ( U967.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_98 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U967.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_45 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U967.EF ) ,
    .I0 ( xor_decoded_masks_14_45 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_45 ) ,
    .I0 ( U967.AB ) ,
    .I1 ( U967.CD ) ,
    .I2 ( U967.EF ) ) ;
and ( 
    .Z ( U1138.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_25 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1138.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_25 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1138.EF ) ,
    .I0 ( xor_decoded_masks_9_25 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_25 ) ,
    .I0 ( U1138.AB ) ,
    .I1 ( U1138.CD ) ,
    .I2 ( U1138.EF ) ) ;
and ( 
    .Z ( U433.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_2 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U433.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_2 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U433.EF ) ,
    .I0 ( xor_decoded_masks_5_2 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_2 ) ,
    .I0 ( U433.AB ) ,
    .I1 ( U433.CD ) ,
    .I2 ( U433.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_9_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_2.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_2.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_2.CD ) ,
    .IN ( masks_shift_reg_9_reg_2.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_2.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_2.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_2.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_2.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_2.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_2.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_2.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_2.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_2.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_2.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_2.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_2.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_2 ) ) ;
and ( 
    .Z ( U1248.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_43 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1248.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_43 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1248.EF ) ,
    .I0 ( xor_decoded_masks_13_43 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_43 ) ,
    .I0 ( U1248.AB ) ,
    .I1 ( U1248.CD ) ,
    .I2 ( U1248.EF ) ) ;
and ( 
    .Z ( U964.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_54 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U964.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_1 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U964.EF ) ,
    .I0 ( xor_decoded_masks_12_1 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_1 ) ,
    .I0 ( U964.AB ) ,
    .I1 ( U964.CD ) ,
    .I2 ( U964.EF ) ) ;
and ( 
    .Z ( U1139.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_33 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1139.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_33 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1139.EF ) ,
    .I0 ( xor_decoded_masks_9_33 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_33 ) ,
    .I0 ( U1139.AB ) ,
    .I1 ( U1139.CD ) ,
    .I2 ( U1139.EF ) ) ;
and ( 
    .Z ( U430.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_6 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U430.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_6 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U430.EF ) ,
    .I0 ( xor_decoded_masks_5_6 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_6 ) ,
    .I0 ( U430.AB ) ,
    .I1 ( U430.CD ) ,
    .I2 ( U430.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_9_6 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_5.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_9_reg_5.CDNI_ ) ,
    .IN ( n51 ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_5.CD ) ,
    .IN ( masks_shift_reg_9_reg_5.CDNI_ ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ,
    .A ( GND ) ) ;
not ( 
    .O1 ( masks_shift_reg_9_reg_5.U5.CD_ ) ,
    .IN ( masks_shift_reg_9_reg_5.CD ) ) ;
and ( 
    .Z ( masks_shift_reg_9_reg_5.U5.D_1 ) ,
    .I0 ( masks_shift_reg_9_reg_5.DI_ ) ,
    .I1 ( masks_shift_reg_9_reg_5.U5.CD_ ) ) ;
MUX21 masks_shift_reg_9_reg_5.U5.I2 ( 
    .I0 ( masks_shift_reg_9_reg_5.U5.D_1 ) ,
    .I1 ( masks_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_0 ) ,
    .Q ( masks_shift_reg_9_reg_5.U5.Q1 ) ,
    .S ( masks_shift_reg_9_reg_5.SYNTEST_EXP_ADDED_NET_1 ) ) ;
DFF masks_shift_reg_9_reg_5.U5.I3 ( 
    .CK ( masks_shift_reg_9_reg_5.CPI_ ) ,
    .D ( masks_shift_reg_9_reg_5.U5.Q1 ) ,
    .Q ( masks_shift_reg_9_5 ) ) ;
and ( 
    .Z ( U1249.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_96 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1249.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_43 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1249.EF ) ,
    .I0 ( xor_decoded_masks_14_43 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_43 ) ,
    .I0 ( U1249.AB ) ,
    .I1 ( U1249.CD ) ,
    .I2 ( U1249.EF ) ) ;
and ( 
    .Z ( U416.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_109 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U416.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_2 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U416.EF ) ,
    .I0 ( xor_decoded_masks_2_2 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_2 ) ,
    .I0 ( U416.AB ) ,
    .I1 ( U416.CD ) ,
    .I2 ( U416.EF ) ) ;
and ( 
    .Z ( U862.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_23 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U862.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_23 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U862.EF ) ,
    .I0 ( xor_decoded_masks_0_23 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_23 ) ,
    .I0 ( U862.AB ) ,
    .I1 ( U862.CD ) ,
    .I2 ( U862.EF ) ) ;
and ( 
    .Z ( U417.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_4 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U417.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_4 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U417.EF ) ,
    .I0 ( xor_decoded_masks_3_4 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_4 ) ,
    .I0 ( U417.AB ) ,
    .I1 ( U417.CD ) ,
    .I2 ( U417.EF ) ) ;
and ( 
    .Z ( U861.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_55 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U861.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_1 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U861.EF ) ,
    .I0 ( xor_decoded_masks_1_1 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_1 ) ,
    .I0 ( U861.AB ) ,
    .I1 ( U861.CD ) ,
    .I2 ( U861.EF ) ) ;
and ( 
    .Z ( U418.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_7 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U418.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_7 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U418.EF ) ,
    .I0 ( xor_decoded_masks_3_7 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_7 ) ,
    .I0 ( U418.AB ) ,
    .I1 ( U418.CD ) ,
    .I2 ( U418.EF ) ) ;
and ( 
    .Z ( U860.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_100 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U860.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_46 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U860.EF ) ,
    .I0 ( xor_decoded_masks_1_46 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_46 ) ,
    .I0 ( U860.AB ) ,
    .I1 ( U860.CD ) ,
    .I2 ( U860.EF ) ) ;
and ( 
    .Z ( U419.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_6 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U419.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_6 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U419.EF ) ,
    .I0 ( xor_decoded_masks_3_6 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_6 ) ,
    .I0 ( U419.AB ) ,
    .I1 ( U419.CD ) ,
    .I2 ( U419.EF ) ) ;
and ( 
    .Z ( U867.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_104 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U867.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_51 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U867.EF ) ,
    .I0 ( xor_decoded_masks_8_51 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_51 ) ,
    .I0 ( U867.AB ) ,
    .I1 ( U867.CD ) ,
    .I2 ( U867.EF ) ) ;
and ( 
    .Z ( U731.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_68 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U731.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_15 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U731.EF ) ,
    .I0 ( xor_decoded_masks_8_15 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_15 ) ,
    .I0 ( U731.AB ) ,
    .I1 ( U731.CD ) ,
    .I2 ( U731.EF ) ) ;
and ( 
    .Z ( U1062.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_12 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1062.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_12 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1062.EF ) ,
    .I0 ( xor_decoded_masks_5_12 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_12 ) ,
    .I0 ( U1062.AB ) ,
    .I1 ( U1062.CD ) ,
    .I2 ( U1062.EF ) ) ;
and ( 
    .Z ( U866.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_104 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U866.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_51 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U866.EF ) ,
    .I0 ( xor_decoded_masks_6_51 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_51 ) ,
    .I0 ( U866.AB ) ,
    .I1 ( U866.CD ) ,
    .I2 ( U866.EF ) ) ;
and ( 
    .Z ( U730.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_74 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U730.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_21 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U730.EF ) ,
    .I0 ( xor_decoded_masks_8_21 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_21 ) ,
    .I0 ( U730.AB ) ,
    .I1 ( U730.CD ) ,
    .I2 ( U730.EF ) ) ;
and ( 
    .Z ( U1063.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_26 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1063.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_26 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1063.EF ) ,
    .I0 ( xor_decoded_masks_7_26 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_26 ) ,
    .I0 ( U1063.AB ) ,
    .I1 ( U1063.CD ) ,
    .I2 ( U1063.EF ) ) ;
and ( 
    .Z ( U388.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_18 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U388.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_18 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U388.EF ) ,
    .I0 ( xor_decoded_masks_7_18 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_18 ) ,
    .I0 ( U388.AB ) ,
    .I1 ( U388.CD ) ,
    .I2 ( U388.EF ) ) ;
and ( 
    .Z ( U865.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_16 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U865.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_16 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U865.EF ) ,
    .I0 ( xor_decoded_masks_0_16 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_16 ) ,
    .I0 ( U865.AB ) ,
    .I1 ( U865.CD ) ,
    .I2 ( U865.EF ) ) ;
and ( 
    .Z ( U733.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_70 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U733.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_17 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U733.EF ) ,
    .I0 ( xor_decoded_masks_8_17 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_17 ) ,
    .I0 ( U733.AB ) ,
    .I1 ( U733.CD ) ,
    .I2 ( U733.EF ) ) ;
and ( 
    .Z ( U1060.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_22 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1060.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_22 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1060.EF ) ,
    .I0 ( xor_decoded_masks_5_22 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_22 ) ,
    .I0 ( U1060.AB ) ,
    .I1 ( U1060.CD ) ,
    .I2 ( U1060.EF ) ) ;
and ( 
    .Z ( U389.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_76 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U389.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_23 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U389.EF ) ,
    .I0 ( xor_decoded_masks_8_23 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_23 ) ,
    .I0 ( U389.AB ) ,
    .I1 ( U389.CD ) ,
    .I2 ( U389.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_10.DI_ ) ,
    .IN ( masks_shift_reg_11_10 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_1_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_reg_10.E_ ) ,
    .IN ( edt_update_hfs_netlink_29288 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_11_10 ) ,
    .IN ( masks_hold_reg_11_reg_10.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_11_reg_10.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_11_reg_10.QT ) ,
    .I1 ( masks_hold_reg_11_reg_10.DI_ ) ,
    .Q ( masks_hold_reg_11_reg_10.ED ) ,
    .S ( masks_hold_reg_11_reg_10.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_11_reg_10.U6.CD_ ) ,
    .IN ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_11_reg_10.U6.D_1 ) ,
    .I0 ( masks_hold_reg_11_reg_10.ED ) ,
    .I1 ( masks_hold_reg_11_reg_10.U6.CD_ ) ) ;
MUX21 masks_hold_reg_11_reg_10.U6.I2 ( 
    .I0 ( masks_hold_reg_11_reg_10.U6.D_1 ) ,
    .I1 ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_11_reg_10.U6.Q1 ) ,
    .S ( masks_hold_reg_11_reg_10.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_11_reg_10.U6.I3 ( 
    .CK ( masks_hold_reg_11_reg_10.CPI_ ) ,
    .D ( masks_hold_reg_11_reg_10.U6.Q1 ) ,
    .Q ( masks_hold_reg_11_reg_10.QT ) ) ;
and ( 
    .Z ( U864.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_19 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U864.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_19 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U864.EF ) ,
    .I0 ( xor_decoded_masks_0_19 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_19 ) ,
    .I0 ( U864.AB ) ,
    .I1 ( U864.CD ) ,
    .I2 ( U864.EF ) ) ;
and ( 
    .Z ( U732.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_64 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U732.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_11 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U732.EF ) ,
    .I0 ( xor_decoded_masks_8_11 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_11 ) ,
    .I0 ( U732.AB ) ,
    .I1 ( U732.CD ) ,
    .I2 ( U732.EF ) ) ;
and ( 
    .Z ( U1061.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_8 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1061.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_8 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1061.EF ) ,
    .I0 ( xor_decoded_masks_5_8 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_8 ) ,
    .I0 ( U1061.AB ) ,
    .I1 ( U1061.CD ) ,
    .I2 ( U1061.EF ) ) ;
and ( 
    .Z ( U386.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_31 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U386.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_31 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U386.EF ) ,
    .I0 ( xor_decoded_masks_7_31 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_31 ) ,
    .I0 ( U386.AB ) ,
    .I1 ( U386.CD ) ,
    .I2 ( U386.EF ) ) ;
and ( 
    .Z ( U735.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_86 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U735.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_33 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U735.EF ) ,
    .I0 ( xor_decoded_masks_10_33 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_33 ) ,
    .I0 ( U735.AB ) ,
    .I1 ( U735.CD ) ,
    .I2 ( U735.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_5.DI_ ) ,
    .IN ( n85 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_5.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_5 ) ,
    .IN ( masks_hold_reg_2_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_5.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_2_reg_5.QT ) ,
    .I1 ( masks_hold_reg_2_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_5.ED ) ,
    .S ( masks_hold_reg_2_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_5.ED ) ,
    .I1 ( masks_hold_reg_2_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_2_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_5.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_2_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_5.QT ) ) ;
and ( 
    .Z ( U1066.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_22 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1066.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_22 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1066.EF ) ,
    .I0 ( xor_decoded_masks_7_22 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_22 ) ,
    .I0 ( U1066.AB ) ,
    .I1 ( U1066.CD ) ,
    .I2 ( U1066.EF ) ) ;
and ( 
    .Z ( U387.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_16 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U387.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_16 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U387.EF ) ,
    .I0 ( xor_decoded_masks_7_16 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_16 ) ,
    .I0 ( U387.AB ) ,
    .I1 ( U387.CD ) ,
    .I2 ( U387.EF ) ) ;
and ( 
    .Z ( U734.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_82 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U734.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_29 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U734.EF ) ,
    .I0 ( xor_decoded_masks_10_29 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_29 ) ,
    .I0 ( U734.AB ) ,
    .I1 ( U734.CD ) ,
    .I2 ( U734.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_2_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_4.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_4 ) ,
    .IN ( masks_hold_reg_2_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_4.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_2_reg_4.QT ) ,
    .I1 ( masks_hold_reg_2_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_4.ED ) ,
    .S ( masks_hold_reg_2_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_4.ED ) ,
    .I1 ( masks_hold_reg_2_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_2_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_4.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_2_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_4.QT ) ) ;
and ( 
    .Z ( U1067.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_8 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1067.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_8 ) ,
    .I1 ( n66 ) ) ;
and ( 
    .Z ( U1067.EF ) ,
    .I0 ( xor_decoded_masks_7_8 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_8 ) ,
    .I0 ( U1067.AB ) ,
    .I1 ( U1067.CD ) ,
    .I2 ( U1067.EF ) ) ;
and ( 
    .Z ( U384.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_28 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U384.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_28 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U384.EF ) ,
    .I0 ( xor_decoded_masks_7_28 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_28 ) ,
    .I0 ( U384.AB ) ,
    .I1 ( U384.CD ) ,
    .I2 ( U384.EF ) ) ;
and ( 
    .Z ( U737.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_90 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U737.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_37 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U737.EF ) ,
    .I0 ( xor_decoded_masks_10_37 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_37 ) ,
    .I0 ( U737.AB ) ,
    .I1 ( U737.CD ) ,
    .I2 ( U737.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_2_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_7.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_7 ) ,
    .IN ( masks_hold_reg_2_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_7.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_2_reg_7.QT ) ,
    .I1 ( masks_hold_reg_2_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_7.ED ) ,
    .S ( masks_hold_reg_2_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_7.ED ) ,
    .I1 ( masks_hold_reg_2_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_2_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_7.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_2_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_7.QT ) ) ;
and ( 
    .Z ( U1064.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_34 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1064.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_34 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1064.EF ) ,
    .I0 ( xor_decoded_masks_7_34 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_34 ) ,
    .I0 ( U1064.AB ) ,
    .I1 ( U1064.CD ) ,
    .I2 ( U1064.EF ) ) ;
and ( 
    .Z ( U385.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_30 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U385.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_30 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U385.EF ) ,
    .I0 ( xor_decoded_masks_7_30 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_30 ) ,
    .I0 ( U385.AB ) ,
    .I1 ( U385.CD ) ,
    .I2 ( U385.EF ) ) ;
and ( 
    .Z ( U736.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_78 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U736.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_25 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U736.EF ) ,
    .I0 ( xor_decoded_masks_10_25 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_25 ) ,
    .I0 ( U736.AB ) ,
    .I1 ( U736.CD ) ,
    .I2 ( U736.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_6.DI_ ) ,
    .IN ( n84 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_6.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_6 ) ,
    .IN ( masks_hold_reg_2_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_6.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_2_reg_6.QT ) ,
    .I1 ( masks_hold_reg_2_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_6.ED ) ,
    .S ( masks_hold_reg_2_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_6.ED ) ,
    .I1 ( masks_hold_reg_2_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_2_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_6.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_2_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_6.QT ) ) ;
and ( 
    .Z ( U1065.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_38 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1065.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_38 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1065.EF ) ,
    .I0 ( xor_decoded_masks_7_38 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_38 ) ,
    .I0 ( U1065.AB ) ,
    .I1 ( U1065.CD ) ,
    .I2 ( U1065.EF ) ) ;
and ( 
    .Z ( U382.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_16 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U382.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_16 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U382.EF ) ,
    .I0 ( xor_decoded_masks_5_16 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_16 ) ,
    .I0 ( U382.AB ) ,
    .I1 ( U382.CD ) ,
    .I2 ( U382.EF ) ) ;
and ( 
    .Z ( U739.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_86 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U739.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_33 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U739.EF ) ,
    .I0 ( xor_decoded_masks_12_33 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_33 ) ,
    .I0 ( U739.AB ) ,
    .I1 ( U739.CD ) ,
    .I2 ( U739.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_1.DI_ ) ,
    .IN ( n97 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_1.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_1 ) ,
    .IN ( masks_hold_reg_2_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_1.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_2_reg_1.QT ) ,
    .I1 ( masks_hold_reg_2_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_1.ED ) ,
    .S ( masks_hold_reg_2_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_1.ED ) ,
    .I1 ( masks_hold_reg_2_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_2_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_1.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_2_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_1.QT ) ) ;
and ( 
    .Z ( U383.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_18 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U383.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_18 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U383.EF ) ,
    .I0 ( xor_decoded_masks_5_18 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_18 ) ,
    .I0 ( U383.AB ) ,
    .I1 ( U383.CD ) ,
    .I2 ( U383.EF ) ) ;
and ( 
    .Z ( U656.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_77 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U656.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_24 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U656.EF ) ,
    .I0 ( xor_decoded_masks_12_24 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_24 ) ,
    .I0 ( U656.AB ) ,
    .I1 ( U656.CD ) ,
    .I2 ( U656.EF ) ) ;
and ( 
    .Z ( U738.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_82 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U738.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_29 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U738.EF ) ,
    .I0 ( xor_decoded_masks_12_29 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_29 ) ,
    .I0 ( U738.AB ) ,
    .I1 ( U738.CD ) ,
    .I2 ( U738.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_2_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_0.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_0 ) ,
    .IN ( masks_hold_reg_2_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_0.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_2_reg_0.QT ) ,
    .I1 ( masks_hold_reg_2_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_0.ED ) ,
    .S ( masks_hold_reg_2_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_0.ED ) ,
    .I1 ( masks_hold_reg_2_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_2_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_0.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_2_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_0.QT ) ) ;
and ( 
    .Z ( U380.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_30 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U380.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_30 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U380.EF ) ,
    .I0 ( xor_decoded_masks_5_30 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_30 ) ,
    .I0 ( U380.AB ) ,
    .I1 ( U380.CD ) ,
    .I2 ( U380.EF ) ) ;
and ( 
    .Z ( U657.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_85 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U657.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_32 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U657.EF ) ,
    .I0 ( xor_decoded_masks_14_32 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_32 ) ,
    .I0 ( U657.AB ) ,
    .I1 ( U657.CD ) ,
    .I2 ( U657.EF ) ) ;
and ( 
    .Z ( U1105.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_95 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1105.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_42 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1105.EF ) ,
    .I0 ( xor_decoded_masks_8_42 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_42 ) ,
    .I0 ( U1105.AB ) ,
    .I1 ( U1105.CD ) ,
    .I2 ( U1105.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_3.DI_ ) ,
    .IN ( n78 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_3.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_3 ) ,
    .IN ( masks_hold_reg_2_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_3.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_2_reg_3.QT ) ,
    .I1 ( masks_hold_reg_2_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_3.ED ) ,
    .S ( masks_hold_reg_2_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_3.ED ) ,
    .I1 ( masks_hold_reg_2_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_2_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_3.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_2_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_3.QT ) ) ;
and ( 
    .Z ( U1068.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_12 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1068.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_12 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1068.EF ) ,
    .I0 ( xor_decoded_masks_7_12 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_12 ) ,
    .I0 ( U1068.AB ) ,
    .I1 ( U1068.CD ) ,
    .I2 ( U1068.EF ) ) ;
and ( 
    .Z ( U381.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_31 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U381.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_31 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U381.EF ) ,
    .I0 ( xor_decoded_masks_5_31 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_31 ) ,
    .I0 ( U381.AB ) ,
    .I1 ( U381.CD ) ,
    .I2 ( U381.EF ) ) ;
and ( 
    .Z ( U959.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_54 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U959.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_1 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U959.EF ) ,
    .I0 ( xor_decoded_masks_10_1 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_1 ) ,
    .I0 ( U959.AB ) ,
    .I1 ( U959.CD ) ,
    .I2 ( U959.EF ) ) ;
and ( 
    .Z ( U654.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_85 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U654.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_32 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U654.EF ) ,
    .I0 ( xor_decoded_masks_10_32 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_32 ) ,
    .I0 ( U654.AB ) ,
    .I1 ( U654.CD ) ,
    .I2 ( U654.EF ) ) ;
and ( 
    .Z ( U1104.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_42 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1104.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_42 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1104.EF ) ,
    .I0 ( xor_decoded_masks_7_42 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_42 ) ,
    .I0 ( U1104.AB ) ,
    .I1 ( U1104.CD ) ,
    .I2 ( U1104.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_2_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_2.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_2 ) ,
    .IN ( masks_hold_reg_2_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_2.SYNTEST_VL_LSI_MUX21_18873.I0 ( 
    .I0 ( masks_hold_reg_2_reg_2.QT ) ,
    .I1 ( masks_hold_reg_2_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_2.ED ) ,
    .S ( masks_hold_reg_2_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_14 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_2.ED ) ,
    .I1 ( masks_hold_reg_2_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_12 ) ,
    .Q ( masks_hold_reg_2_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_2.SYNTEST_EXP_ADDED_NET_13 ) ) ;
DFF masks_hold_reg_2_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_2.QT ) ) ;
and ( 
    .Z ( U1069.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_61 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1069.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_8 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1069.EF ) ,
    .I0 ( xor_decoded_masks_8_8 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_8 ) ,
    .I0 ( U1069.AB ) ,
    .I1 ( U1069.CD ) ,
    .I2 ( U1069.EF ) ) ;
and ( 
    .Z ( U958.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_58 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U958.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_5 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U958.EF ) ,
    .I0 ( xor_decoded_masks_10_5 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_5 ) ,
    .I0 ( U958.AB ) ,
    .I1 ( U958.CD ) ,
    .I2 ( U958.EF ) ) ;
and ( 
    .Z ( U655.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_85 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U655.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_32 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U655.EF ) ,
    .I0 ( xor_decoded_masks_12_32 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_32 ) ,
    .I0 ( U655.AB ) ,
    .I1 ( U655.CD ) ,
    .I2 ( U655.EF ) ) ;
and ( 
    .Z ( U1107.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_95 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1107.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_42 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1107.EF ) ,
    .I0 ( xor_decoded_masks_10_42 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_42 ) ,
    .I0 ( U1107.AB ) ,
    .I1 ( U1107.CD ) ,
    .I2 ( U1107.EF ) ) ;
and ( 
    .Z ( U652.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_63 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U652.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_10 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U652.EF ) ,
    .I0 ( xor_decoded_masks_8_10 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_10 ) ,
    .I0 ( U652.AB ) ,
    .I1 ( U652.CD ) ,
    .I2 ( U652.EF ) ) ;
and ( 
    .Z ( U1106.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_42 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1106.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_42 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1106.EF ) ,
    .I0 ( xor_decoded_masks_9_42 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_42 ) ,
    .I0 ( U1106.AB ) ,
    .I1 ( U1106.CD ) ,
    .I2 ( U1106.EF ) ) ;
and ( 
    .Z ( U653.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_69 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U653.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_16 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U653.EF ) ,
    .I0 ( xor_decoded_masks_8_16 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_16 ) ,
    .I0 ( U653.AB ) ,
    .I1 ( U653.CD ) ,
    .I2 ( U653.EF ) ) ;
and ( 
    .Z ( U1101.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_95 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1101.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_42 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1101.EF ) ,
    .I0 ( xor_decoded_masks_4_42 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_42 ) ,
    .I0 ( U1101.AB ) ,
    .I1 ( U1101.CD ) ,
    .I2 ( U1101.EF ) ) ;
and ( 
    .Z ( U650.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_89 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U650.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_36 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U650.EF ) ,
    .I0 ( xor_decoded_masks_8_36 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_36 ) ,
    .I0 ( U650.AB ) ,
    .I1 ( U650.CD ) ,
    .I2 ( U650.EF ) ) ;
and ( 
    .Z ( U1100.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_42 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1100.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_42 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1100.EF ) ,
    .I0 ( xor_decoded_masks_3_42 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_42 ) ,
    .I0 ( U1100.AB ) ,
    .I1 ( U1100.CD ) ,
    .I2 ( U1100.EF ) ) ;
and ( 
    .Z ( U651.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_67 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U651.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_14 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U651.EF ) ,
    .I0 ( xor_decoded_masks_8_14 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_14 ) ,
    .I0 ( U651.AB ) ,
    .I1 ( U651.CD ) ,
    .I2 ( U651.EF ) ) ;
and ( 
    .Z ( U1103.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_95 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1103.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_42 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1103.EF ) ,
    .I0 ( xor_decoded_masks_6_42 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_42 ) ,
    .I0 ( U1103.AB ) ,
    .I1 ( U1103.CD ) ,
    .I2 ( U1103.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_2_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_9.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_9 ) ,
    .IN ( masks_hold_reg_2_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_2_reg_9.QT ) ,
    .I1 ( masks_hold_reg_2_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_9.ED ) ,
    .S ( masks_hold_reg_2_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_9.ED ) ,
    .I1 ( masks_hold_reg_2_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_2_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_2_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_9.QT ) ) ;
and ( 
    .Z ( U1102.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_42 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1102.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_42 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1102.EF ) ,
    .I0 ( xor_decoded_masks_5_42 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_42 ) ,
    .I0 ( U1102.AB ) ,
    .I1 ( U1102.CD ) ,
    .I2 ( U1102.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_8_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_9.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_9.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_9 ) ,
    .IN ( masks_hold_reg_8_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_9.QT ) ,
    .I1 ( masks_hold_reg_8_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_9.ED ) ,
    .S ( masks_hold_reg_8_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_9.ED ) ,
    .I1 ( masks_hold_reg_8_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_9.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_2_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2641 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_reg_8.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_2_8 ) ,
    .IN ( masks_hold_reg_2_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_4 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_5 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_6 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_2_reg_8.SYNTEST_VL_LSI_MUX21_16157.I0 ( 
    .I0 ( masks_hold_reg_2_reg_8.QT ) ,
    .I1 ( masks_hold_reg_2_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_2_reg_8.ED ) ,
    .S ( masks_hold_reg_2_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_2_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_6 ) ) ;
and ( 
    .Z ( masks_hold_reg_2_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_2_reg_8.ED ) ,
    .I1 ( masks_hold_reg_2_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_2_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_2_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_4 ) ,
    .Q ( masks_hold_reg_2_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_2_reg_8.SYNTEST_EXP_ADDED_NET_5 ) ) ;
DFF masks_hold_reg_2_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_2_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_2_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_2_reg_8.QT ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_8_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_8.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_8.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_8 ) ,
    .IN ( masks_hold_reg_8_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_8.QT ) ,
    .I1 ( masks_hold_reg_8_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_8.ED ) ,
    .S ( masks_hold_reg_8_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_8.ED ) ,
    .I1 ( masks_hold_reg_8_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_8.QT ) ) ;
and ( 
    .Z ( U951.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_45 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U951.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_45 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U951.EF ) ,
    .I0 ( xor_decoded_masks_7_45 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_45 ) ,
    .I0 ( U951.AB ) ,
    .I1 ( U951.CD ) ,
    .I2 ( U951.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_8_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_7.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_7.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_7 ) ,
    .IN ( masks_hold_reg_8_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_7.QT ) ,
    .I1 ( masks_hold_reg_8_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_7.ED ) ,
    .S ( masks_hold_reg_8_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_7.ED ) ,
    .I1 ( masks_hold_reg_8_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_7.QT ) ) ;
and ( 
    .Z ( U950.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_54 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U950.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_1 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U950.EF ) ,
    .I0 ( xor_decoded_masks_6_1 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_1 ) ,
    .I0 ( U950.AB ) ,
    .I1 ( U950.CD ) ,
    .I2 ( U950.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_8_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_6.CPI_ ) ,
    .IN ( edt_clock_cts_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_6.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_6 ) ,
    .IN ( masks_hold_reg_8_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_6.QT ) ,
    .I1 ( masks_hold_reg_8_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_6.ED ) ,
    .S ( masks_hold_reg_8_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_6.ED ) ,
    .I1 ( masks_hold_reg_8_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_6.QT ) ) ;
not ( 
    .O1 ( n10 ) ,
    .IN ( masks_shift_reg_3_9 ) ) ;
and ( 
    .Z ( U953.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_1 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U953.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_1 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U953.EF ) ,
    .I0 ( xor_decoded_masks_7_1 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_1 ) ,
    .I0 ( U953.AB ) ,
    .I1 ( U953.CD ) ,
    .I2 ( U953.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_8_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_5.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_5 ) ,
    .IN ( masks_hold_reg_8_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_5.QT ) ,
    .I1 ( masks_hold_reg_8_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_5.ED ) ,
    .S ( masks_hold_reg_8_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_5.ED ) ,
    .I1 ( masks_hold_reg_8_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_5.QT ) ) ;
or ( 
    .Z ( U1298.AB ) ,
    .I0 ( n44 ) ,
    .I1 ( n10 ) ) ;
or ( 
    .Z ( U1298.CD ) ,
    .I0 ( n41 ) ,
    .I1 ( n11 ) ) ;
and ( 
    .Z ( U1298.ZN ) ,
    .I0 ( U1298.AB ) ,
    .I1 ( U1298.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_4 ) ,
    .IN ( U1298.ZN ) ) ;
and ( 
    .Z ( U952.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_5 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U952.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_5 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U952.EF ) ,
    .I0 ( xor_decoded_masks_7_5 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_5 ) ,
    .I0 ( U952.AB ) ,
    .I1 ( U952.CD ) ,
    .I2 ( U952.EF ) ) ;
and ( 
    .Z ( U1109.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_95 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1109.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_42 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1109.EF ) ,
    .I0 ( xor_decoded_masks_12_42 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_42 ) ,
    .I0 ( U1109.AB ) ,
    .I1 ( U1109.CD ) ,
    .I2 ( U1109.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_8_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_4.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_4 ) ,
    .IN ( masks_hold_reg_8_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_4.QT ) ,
    .I1 ( masks_hold_reg_8_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_4.ED ) ,
    .S ( masks_hold_reg_8_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_4.ED ) ,
    .I1 ( masks_hold_reg_8_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_4.QT ) ) ;
and ( 
    .Z ( U878.AB ) ,
    .I0 ( masks_hold_reg_12_1 ) ,
    .I1 ( edt_configuration_hfs_netlink_29292 ) ) ;
and ( 
    .Z ( U878.CD ) ,
    .I0 ( config1_xor_encoded_masks_140 ) ,
    .I1 ( edt_configuration_hfs_netlink_29291 ) ) ;
or ( 
    .Z ( xor_encoded_masks_140 ) ,
    .I0 ( U878.AB ) ,
    .I1 ( U878.CD ) ) ;
not ( 
    .O1 ( n6 ) ,
    .IN ( masks_shift_reg_7_9 ) ) ;
and ( 
    .Z ( U955.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_54 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U955.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_1 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U955.EF ) ,
    .I0 ( xor_decoded_masks_8_1 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_1 ) ,
    .I0 ( U955.AB ) ,
    .I1 ( U955.CD ) ,
    .I2 ( U955.EF ) ) ;
and ( 
    .Z ( U658.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_77 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U658.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_24 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U658.EF ) ,
    .I0 ( xor_decoded_masks_14_24 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_24 ) ,
    .I0 ( U658.AB ) ,
    .I1 ( U658.CD ) ,
    .I2 ( U658.EF ) ) ;
and ( 
    .Z ( U1108.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_42 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1108.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_42 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1108.EF ) ,
    .I0 ( xor_decoded_masks_11_42 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_42 ) ,
    .I0 ( U1108.AB ) ,
    .I1 ( U1108.CD ) ,
    .I2 ( U1108.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_8_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_3.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_3 ) ,
    .IN ( masks_hold_reg_8_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_3.QT ) ,
    .I1 ( masks_hold_reg_8_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_3.ED ) ,
    .S ( masks_hold_reg_8_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_3.ED ) ,
    .I1 ( masks_hold_reg_8_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_3.QT ) ) ;
and ( 
    .Z ( U879.AB ) ,
    .I0 ( masks_hold_reg_1_0 ) ,
    .I1 ( n39 ) ) ;
and ( 
    .Z ( U879.CD ) ,
    .I0 ( config1_xor_encoded_masks_20 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_20 ) ,
    .I0 ( U879.AB ) ,
    .I1 ( U879.CD ) ) ;
or ( 
    .Z ( U1296.AB ) ,
    .I0 ( n43 ) ,
    .I1 ( n6 ) ) ;
or ( 
    .Z ( U1296.CD ) ,
    .I0 ( n40 ) ,
    .I1 ( n7 ) ) ;
and ( 
    .Z ( U1296.ZN ) ,
    .I0 ( U1296.AB ) ,
    .I1 ( U1296.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_8 ) ,
    .IN ( U1296.ZN ) ) ;
and ( 
    .Z ( U954.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_98 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U954.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_45 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U954.EF ) ,
    .I0 ( xor_decoded_masks_8_45 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_45 ) ,
    .I0 ( U954.AB ) ,
    .I1 ( U954.CD ) ,
    .I2 ( U954.EF ) ) ;
and ( 
    .Z ( U975.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_59 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U975.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_5 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U975.EF ) ,
    .I0 ( xor_decoded_masks_1_5 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_5 ) ,
    .I0 ( U975.AB ) ,
    .I1 ( U975.CD ) ,
    .I2 ( U975.EF ) ) ;
and ( 
    .Z ( U848.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_47 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U848.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_47 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U848.EF ) ,
    .I0 ( xor_decoded_masks_11_47 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_47 ) ,
    .I0 ( U848.AB ) ,
    .I1 ( U848.CD ) ,
    .I2 ( U848.EF ) ) ;
and ( 
    .Z ( U1289.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_50 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1289.CD ) ,
    .I0 ( config0_onehot_decoded_masks_13_50 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1289.EF ) ,
    .I0 ( xor_decoded_masks_13_50 ) ,
    .I1 ( n30 ) ) ;
or ( 
    .Z ( masks_for_compactor_13_50 ) ,
    .I0 ( U1289.AB ) ,
    .I1 ( U1289.CD ) ,
    .I2 ( U1289.EF ) ) ;
and ( 
    .Z ( U925.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_18 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U925.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_18 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U925.EF ) ,
    .I0 ( xor_decoded_masks_0_18 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_18 ) ,
    .I0 ( U925.AB ) ,
    .I1 ( U925.CD ) ,
    .I2 ( U925.EF ) ) ;
and ( 
    .Z ( U1286.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_103 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1286.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_50 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1286.EF ) ,
    .I0 ( xor_decoded_masks_10_50 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_50 ) ,
    .I0 ( U1286.AB ) ,
    .I1 ( U1286.CD ) ,
    .I2 ( U1286.EF ) ) ;
and ( 
    .Z ( U922.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_46 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U922.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_46 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U922.EF ) ,
    .I0 ( xor_decoded_masks_11_46 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_46 ) ,
    .I0 ( U922.AB ) ,
    .I1 ( U922.CD ) ,
    .I2 ( U922.EF ) ) ;
and ( 
    .Z ( U1287.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_50 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1287.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_50 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1287.EF ) ,
    .I0 ( xor_decoded_masks_11_50 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_50 ) ,
    .I0 ( U1287.AB ) ,
    .I1 ( U1287.CD ) ,
    .I2 ( U1287.EF ) ) ;
and ( 
    .Z ( U923.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_99 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U923.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_46 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U923.EF ) ,
    .I0 ( xor_decoded_masks_12_46 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_46 ) ,
    .I0 ( U923.AB ) ,
    .I1 ( U923.CD ) ,
    .I2 ( U923.EF ) ) ;
and ( 
    .Z ( U1284.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_103 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1284.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_50 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1284.EF ) ,
    .I0 ( xor_decoded_masks_8_50 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_50 ) ,
    .I0 ( U1284.AB ) ,
    .I1 ( U1284.CD ) ,
    .I2 ( U1284.EF ) ) ;
and ( 
    .Z ( U920.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_46 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U920.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_46 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U920.EF ) ,
    .I0 ( xor_decoded_masks_9_46 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_46 ) ,
    .I0 ( U920.AB ) ,
    .I1 ( U920.CD ) ,
    .I2 ( U920.EF ) ) ;
and ( 
    .Z ( U659.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_89 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U659.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_36 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U659.EF ) ,
    .I0 ( xor_decoded_masks_14_36 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_36 ) ,
    .I0 ( U659.AB ) ,
    .I1 ( U659.CD ) ,
    .I2 ( U659.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_8_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_2.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_2 ) ,
    .IN ( masks_hold_reg_8_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_2.QT ) ,
    .I1 ( masks_hold_reg_8_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_2.ED ) ,
    .S ( masks_hold_reg_8_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_2.ED ) ,
    .I1 ( masks_hold_reg_8_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_2.QT ) ) ;
not ( 
    .O1 ( n14 ) ,
    .IN ( masks_shift_reg_9_9 ) ) ;
and ( 
    .Z ( U957.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_1 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U957.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_1 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U957.EF ) ,
    .I0 ( xor_decoded_masks_9_1 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_1 ) ,
    .I0 ( U957.AB ) ,
    .I1 ( U957.CD ) ,
    .I2 ( U957.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_8_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_1.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_1 ) ,
    .IN ( masks_hold_reg_8_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_1.QT ) ,
    .I1 ( masks_hold_reg_8_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_1.ED ) ,
    .S ( masks_hold_reg_8_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_1.ED ) ,
    .I1 ( masks_hold_reg_8_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_1.QT ) ) ;
or ( 
    .Z ( U1294.AB ) ,
    .I0 ( n45 ) ,
    .I1 ( n14 ) ) ;
or ( 
    .Z ( U1294.CD ) ,
    .I0 ( edt_configuration_hfs_netlink_29290 ) ,
    .I1 ( n15 ) ) ;
and ( 
    .Z ( U1294.ZN ) ,
    .I0 ( U1294.AB ) ,
    .I1 ( U1294.CD ) ) ;
not ( 
    .O1 ( edt_channels_out_from_controller_10 ) ,
    .IN ( U1294.ZN ) ) ;
and ( 
    .Z ( U956.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_45 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U956.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_45 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U956.EF ) ,
    .I0 ( xor_decoded_masks_9_45 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_45 ) ,
    .I0 ( U956.AB ) ,
    .I1 ( U956.CD ) ,
    .I2 ( U956.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_8_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2861 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_reg_0.E_ ) ,
    .IN ( n49 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_8_0 ) ,
    .IN ( masks_hold_reg_8_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_8_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_8_reg_0.QT ) ,
    .I1 ( masks_hold_reg_8_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_8_reg_0.ED ) ,
    .S ( masks_hold_reg_8_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_8_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_8_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_8_reg_0.ED ) ,
    .I1 ( masks_hold_reg_8_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_8_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_8_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_8_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_8_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_8_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_8_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_8_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_8_reg_0.QT ) ) ;
and ( 
    .Z ( U1293.AB ) ,
    .I0 ( n91 ) ,
    .I1 ( n38 ) ) ;
and ( 
    .Z ( U1293.CD ) ,
    .I0 ( config1_xor_encoded_masks_40 ) ,
    .I1 ( n37 ) ) ;
or ( 
    .Z ( xor_encoded_masks_40 ) ,
    .I0 ( U1293.AB ) ,
    .I1 ( U1293.CD ) ) ;
and ( 
    .Z ( U872.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_31 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U872.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_31 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U872.EF ) ,
    .I0 ( xor_decoded_masks_0_31 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_31 ) ,
    .I0 ( U872.AB ) ,
    .I1 ( U872.CD ) ,
    .I2 ( U872.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_6.DI_ ) ,
    .IN ( masks_shift_reg_1_6 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_6.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_6.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_6 ) ,
    .IN ( masks_hold_reg_1_reg_6.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_6.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_6.QT ) ,
    .I1 ( masks_hold_reg_1_reg_6.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_6.ED ) ,
    .S ( masks_hold_reg_1_reg_6.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_6.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_6.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_6.ED ) ,
    .I1 ( masks_hold_reg_1_reg_6.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_6.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_6.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_6.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_6.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_6.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_6.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_6.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_6.QT ) ) ;
and ( 
    .Z ( U1291.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_104 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U1291.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_50 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U1291.EF ) ,
    .I0 ( xor_decoded_masks_1_50 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_50 ) ,
    .I0 ( U1291.AB ) ,
    .I1 ( U1291.CD ) ,
    .I2 ( U1291.EF ) ) ;
and ( 
    .Z ( U873.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_29 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U873.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_29 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U873.EF ) ,
    .I0 ( xor_decoded_masks_0_29 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_29 ) ,
    .I0 ( U873.AB ) ,
    .I1 ( U873.CD ) ,
    .I2 ( U873.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_7.DI_ ) ,
    .IN ( masks_shift_reg_1_7 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_7.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_7.E_ ) ,
    .IN ( n47 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_7 ) ,
    .IN ( masks_hold_reg_1_reg_7.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_7.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_7.QT ) ,
    .I1 ( masks_hold_reg_1_reg_7.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_7.ED ) ,
    .S ( masks_hold_reg_1_reg_7.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_7.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_7.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_7.ED ) ,
    .I1 ( masks_hold_reg_1_reg_7.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_7.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_7.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_7.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_7.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_7.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_7.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_7.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_7.QT ) ) ;
and ( 
    .Z ( U1290.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_103 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U1290.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_50 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U1290.EF ) ,
    .I0 ( xor_decoded_masks_14_50 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_50 ) ,
    .I0 ( U1290.AB ) ,
    .I1 ( U1290.CD ) ,
    .I2 ( U1290.EF ) ) ;
and ( 
    .Z ( U870.AB ) ,
    .I0 ( config1_onehot_decoded_masks_6_104 ) ,
    .I1 ( n58 ) ) ;
and ( 
    .Z ( U870.CD ) ,
    .I0 ( config0_onehot_decoded_masks_14_51 ) ,
    .I1 ( n69 ) ) ;
and ( 
    .Z ( U870.EF ) ,
    .I0 ( xor_decoded_masks_14_51 ) ,
    .I1 ( n31 ) ) ;
or ( 
    .Z ( masks_for_compactor_14_51 ) ,
    .I0 ( U870.AB ) ,
    .I1 ( U870.CD ) ,
    .I2 ( U870.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_4.DI_ ) ,
    .IN ( masks_shift_reg_1_4 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_4.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_4.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_4 ) ,
    .IN ( masks_hold_reg_1_reg_4.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_4.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_4.QT ) ,
    .I1 ( masks_hold_reg_1_reg_4.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_4.ED ) ,
    .S ( masks_hold_reg_1_reg_4.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_4.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_4.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_4.ED ) ,
    .I1 ( masks_hold_reg_1_reg_4.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_4.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_4.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_4.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_4.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_4.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_4.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_4.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_4.QT ) ) ;
and ( 
    .Z ( U871.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_105 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U871.CD ) ,
    .I0 ( config0_onehot_decoded_masks_1_51 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U871.EF ) ,
    .I0 ( xor_decoded_masks_1_51 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_1_51 ) ,
    .I0 ( U871.AB ) ,
    .I1 ( U871.CD ) ,
    .I2 ( U871.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_5.DI_ ) ,
    .IN ( masks_shift_reg_1_5 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_5.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_5.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_5 ) ,
    .IN ( masks_hold_reg_1_reg_5.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_5.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_5.QT ) ,
    .I1 ( masks_hold_reg_1_reg_5.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_5.ED ) ,
    .S ( masks_hold_reg_1_reg_5.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_5.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_5.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_5.ED ) ,
    .I1 ( masks_hold_reg_1_reg_5.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_5.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_5.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_5.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_5.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_5.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_5.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_5.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_5.QT ) ) ;
and ( 
    .Z ( U876.AB ) ,
    .I0 ( masks_hold_reg_5_4 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U876.CD ) ,
    .I0 ( config1_xor_encoded_masks_60 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_60 ) ,
    .I0 ( U876.AB ) ,
    .I1 ( U876.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_2.DI_ ) ,
    .IN ( masks_shift_reg_1_2 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_2.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_2.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_2 ) ,
    .IN ( masks_hold_reg_1_reg_2.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_2.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_2.QT ) ,
    .I1 ( masks_hold_reg_1_reg_2.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_2.ED ) ,
    .S ( masks_hold_reg_1_reg_2.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_2.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_2.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_2.ED ) ,
    .I1 ( masks_hold_reg_1_reg_2.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_2.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_2.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_2.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_2.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_2.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_2.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_2.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_2.QT ) ) ;
and ( 
    .Z ( U702.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_136 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U702.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_29 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U702.EF ) ,
    .I0 ( xor_decoded_masks_2_29 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_29 ) ,
    .I0 ( U702.AB ) ,
    .I1 ( U702.CD ) ,
    .I2 ( U702.EF ) ) ;
and ( 
    .Z ( U1051.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_38 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1051.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_38 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1051.EF ) ,
    .I0 ( xor_decoded_masks_3_38 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_38 ) ,
    .I0 ( U1051.AB ) ,
    .I1 ( U1051.CD ) ,
    .I2 ( U1051.EF ) ) ;
and ( 
    .Z ( U877.AB ) ,
    .I0 ( masks_hold_reg_7_6 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U877.CD ) ,
    .I0 ( config1_xor_encoded_masks_80 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_80 ) ,
    .I0 ( U877.AB ) ,
    .I1 ( U877.CD ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_3.DI_ ) ,
    .IN ( masks_shift_reg_1_3 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_3.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_3.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_3 ) ,
    .IN ( masks_hold_reg_1_reg_3.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_3.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_3.QT ) ,
    .I1 ( masks_hold_reg_1_reg_3.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_3.ED ) ,
    .S ( masks_hold_reg_1_reg_3.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_3.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_3.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_3.ED ) ,
    .I1 ( masks_hold_reg_1_reg_3.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_3.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_3.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_3.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_3.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_3.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_3.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_3.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_3.QT ) ) ;
and ( 
    .Z ( U703.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_132 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U703.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_25 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U703.EF ) ,
    .I0 ( xor_decoded_masks_2_25 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_25 ) ,
    .I0 ( U703.AB ) ,
    .I1 ( U703.CD ) ,
    .I2 ( U703.EF ) ) ;
and ( 
    .Z ( U1050.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_30 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1050.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_30 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1050.EF ) ,
    .I0 ( xor_decoded_masks_3_30 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_30 ) ,
    .I0 ( U1050.AB ) ,
    .I1 ( U1050.CD ) ,
    .I2 ( U1050.EF ) ) ;
and ( 
    .Z ( U874.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_27 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U874.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_27 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U874.EF ) ,
    .I0 ( xor_decoded_masks_0_27 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_27 ) ,
    .I0 ( U874.AB ) ,
    .I1 ( U874.CD ) ,
    .I2 ( U874.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_0.DI_ ) ,
    .IN ( masks_shift_reg_1_0 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_0.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_0.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_0 ) ,
    .IN ( masks_hold_reg_1_reg_0.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_0.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_0.QT ) ,
    .I1 ( masks_hold_reg_1_reg_0.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_0.ED ) ,
    .S ( masks_hold_reg_1_reg_0.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_0.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_0.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_0.ED ) ,
    .I1 ( masks_hold_reg_1_reg_0.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_0.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_0.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_0.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_0.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_0.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_0.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_0.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_0.QT ) ) ;
and ( 
    .Z ( U700.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_45 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U700.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_45 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U700.EF ) ,
    .I0 ( xor_decoded_masks_0_45 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_45 ) ,
    .I0 ( U700.AB ) ,
    .I1 ( U700.CD ) ,
    .I2 ( U700.EF ) ) ;
and ( 
    .Z ( U1053.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_18 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1053.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_18 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1053.EF ) ,
    .I0 ( xor_decoded_masks_3_18 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_18 ) ,
    .I0 ( U1053.AB ) ,
    .I1 ( U1053.CD ) ,
    .I2 ( U1053.EF ) ) ;
and ( 
    .Z ( U875.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_24 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U875.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_24 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U875.EF ) ,
    .I0 ( xor_decoded_masks_0_24 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_24 ) ,
    .I0 ( U875.AB ) ,
    .I1 ( U875.CD ) ,
    .I2 ( U875.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_1.DI_ ) ,
    .IN ( masks_shift_reg_1_1 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_1.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_1.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_1 ) ,
    .IN ( masks_hold_reg_1_reg_1.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_1.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_1.QT ) ,
    .I1 ( masks_hold_reg_1_reg_1.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_1.ED ) ,
    .S ( masks_hold_reg_1_reg_1.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_1.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_1.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_1.ED ) ,
    .I1 ( masks_hold_reg_1_reg_1.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_1.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_1.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_1.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_1.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_1.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_1.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_1.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_1.QT ) ) ;
and ( 
    .Z ( U701.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_37 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U701.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_37 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U701.EF ) ,
    .I0 ( xor_decoded_masks_0_37 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_37 ) ,
    .I0 ( U701.AB ) ,
    .I1 ( U701.CD ) ,
    .I2 ( U701.EF ) ) ;
and ( 
    .Z ( U1052.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_8 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1052.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_8 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1052.EF ) ,
    .I0 ( xor_decoded_masks_3_8 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_8 ) ,
    .I0 ( U1052.AB ) ,
    .I1 ( U1052.CD ) ,
    .I2 ( U1052.EF ) ) ;
and ( 
    .Z ( U397.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_76 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U397.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_23 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U397.EF ) ,
    .I0 ( xor_decoded_masks_10_23 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_23 ) ,
    .I0 ( U397.AB ) ,
    .I1 ( U397.CD ) ,
    .I2 ( U397.EF ) ) ;
and ( 
    .Z ( U706.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_128 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U706.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_21 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U706.EF ) ,
    .I0 ( xor_decoded_masks_2_21 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_21 ) ,
    .I0 ( U706.AB ) ,
    .I1 ( U706.CD ) ,
    .I2 ( U706.EF ) ) ;
and ( 
    .Z ( U1055.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_61 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1055.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_8 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1055.EF ) ,
    .I0 ( xor_decoded_masks_4_8 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_8 ) ,
    .I0 ( U1055.AB ) ,
    .I1 ( U1055.CD ) ,
    .I2 ( U1055.EF ) ) ;
and ( 
    .Z ( U396.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_75 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U396.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_22 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U396.EF ) ,
    .I0 ( xor_decoded_masks_10_22 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_22 ) ,
    .I0 ( U396.AB ) ,
    .I1 ( U396.CD ) ,
    .I2 ( U396.EF ) ) ;
and ( 
    .Z ( U707.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_124 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U707.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_17 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U707.EF ) ,
    .I0 ( xor_decoded_masks_2_17 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_17 ) ,
    .I0 ( U707.AB ) ,
    .I1 ( U707.CD ) ,
    .I2 ( U707.EF ) ) ;
and ( 
    .Z ( U1054.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_12 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1054.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_12 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1054.EF ) ,
    .I0 ( xor_decoded_masks_3_12 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_12 ) ,
    .I0 ( U1054.AB ) ,
    .I1 ( U1054.CD ) ,
    .I2 ( U1054.EF ) ) ;
and ( 
    .Z ( U395.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_19 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U395.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_19 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U395.EF ) ,
    .I0 ( xor_decoded_masks_9_19 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_19 ) ,
    .I0 ( U395.AB ) ,
    .I1 ( U395.CD ) ,
    .I2 ( U395.EF ) ) ;
and ( 
    .Z ( U704.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_140 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U704.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_33 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U704.EF ) ,
    .I0 ( xor_decoded_masks_2_33 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_33 ) ,
    .I0 ( U704.AB ) ,
    .I1 ( U704.CD ) ,
    .I2 ( U704.EF ) ) ;
and ( 
    .Z ( U1057.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_26 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1057.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_26 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1057.EF ) ,
    .I0 ( xor_decoded_masks_5_26 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_26 ) ,
    .I0 ( U1057.AB ) ,
    .I1 ( U1057.CD ) ,
    .I2 ( U1057.EF ) ) ;
and ( 
    .Z ( U394.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_18 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U394.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_18 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U394.EF ) ,
    .I0 ( xor_decoded_masks_9_18 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_18 ) ,
    .I0 ( U394.AB ) ,
    .I1 ( U394.CD ) ,
    .I2 ( U394.EF ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_10.DI_ ) ,
    .IN ( N190 ) ) ;
buf ( 
    .O1 ( masks_shift_reg_8_reg_10.CPI_ ) ,
    .IN ( edt_clock_cts_0_1 ) ) ;
DFF masks_shift_reg_8_reg_10.udp1.I0 ( 
    .CK ( masks_shift_reg_8_reg_10.CPI_ ) ,
    .D ( masks_shift_reg_8_reg_10.DI_ ) ,
    .Q ( masks_shift_reg_8_10 ) ) ;
and ( 
    .Z ( U705.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_144 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U705.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_37 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U705.EF ) ,
    .I0 ( xor_decoded_masks_2_37 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_37 ) ,
    .I0 ( U705.AB ) ,
    .I1 ( U705.CD ) ,
    .I2 ( U705.EF ) ) ;
and ( 
    .Z ( U1056.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_71 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1056.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_18 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1056.EF ) ,
    .I0 ( xor_decoded_masks_4_18 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_18 ) ,
    .I0 ( U1056.AB ) ,
    .I1 ( U1056.CD ) ,
    .I2 ( U1056.EF ) ) ;
and ( 
    .Z ( U393.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_16 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U393.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_16 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U393.EF ) ,
    .I0 ( xor_decoded_masks_9_16 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_16 ) ,
    .I0 ( U393.AB ) ,
    .I1 ( U393.CD ) ,
    .I2 ( U393.EF ) ) ;
and ( 
    .Z ( U1059.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_38 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1059.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_38 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1059.EF ) ,
    .I0 ( xor_decoded_masks_5_38 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_38 ) ,
    .I0 ( U1059.AB ) ,
    .I1 ( U1059.CD ) ,
    .I2 ( U1059.EF ) ) ;
and ( 
    .Z ( U392.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_31 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U392.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_31 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U392.EF ) ,
    .I0 ( xor_decoded_masks_9_31 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_31 ) ,
    .I0 ( U392.AB ) ,
    .I1 ( U392.CD ) ,
    .I2 ( U392.EF ) ) ;
and ( 
    .Z ( U621.AB ) ,
    .I0 ( masks_hold_reg_6_9 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U621.CD ) ,
    .I0 ( config1_xor_encoded_masks_66 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_66 ) ,
    .I0 ( U621.AB ) ,
    .I1 ( U621.CD ) ) ;
and ( 
    .Z ( U1058.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_34 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1058.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_34 ) ,
    .I1 ( n68 ) ) ;
and ( 
    .Z ( U1058.EF ) ,
    .I0 ( xor_decoded_masks_5_34 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_34 ) ,
    .I0 ( U1058.AB ) ,
    .I1 ( U1058.CD ) ,
    .I2 ( U1058.EF ) ) ;
and ( 
    .Z ( U391.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_30 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U391.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_30 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U391.EF ) ,
    .I0 ( xor_decoded_masks_9_30 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_30 ) ,
    .I0 ( U391.AB ) ,
    .I1 ( U391.CD ) ,
    .I2 ( U391.EF ) ) ;
and ( 
    .Z ( U620.AB ) ,
    .I0 ( masks_hold_reg_7_2 ) ,
    .I1 ( n43 ) ) ;
and ( 
    .Z ( U620.CD ) ,
    .I0 ( config1_xor_encoded_masks_84 ) ,
    .I1 ( n40 ) ) ;
or ( 
    .Z ( xor_encoded_masks_84 ) ,
    .I0 ( U620.AB ) ,
    .I1 ( U620.CD ) ) ;
and ( 
    .Z ( U1172.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_94 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1172.CD ) ,
    .I0 ( config0_onehot_decoded_masks_4_41 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1172.EF ) ,
    .I0 ( xor_decoded_masks_4_41 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_4_41 ) ,
    .I0 ( U1172.AB ) ,
    .I1 ( U1172.CD ) ,
    .I2 ( U1172.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_8.DI_ ) ,
    .IN ( masks_shift_reg_1_8 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_8.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_8.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_8 ) ,
    .IN ( masks_hold_reg_1_reg_8.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_8.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_8.QT ) ,
    .I1 ( masks_hold_reg_1_reg_8.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_8.ED ) ,
    .S ( masks_hold_reg_1_reg_8.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_8.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_8.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_8.ED ) ,
    .I1 ( masks_hold_reg_1_reg_8.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_8.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_8.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_8.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_8.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_8.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_8.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_8.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_8.QT ) ) ;
and ( 
    .Z ( U708.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_122 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U708.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_15 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U708.EF ) ,
    .I0 ( xor_decoded_masks_2_15 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_15 ) ,
    .I0 ( U708.AB ) ,
    .I1 ( U708.CD ) ,
    .I2 ( U708.EF ) ) ;
and ( 
    .Z ( U390.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_28 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U390.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_28 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U390.EF ) ,
    .I0 ( xor_decoded_masks_9_28 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_28 ) ,
    .I0 ( U390.AB ) ,
    .I1 ( U390.CD ) ,
    .I2 ( U390.EF ) ) ;
and ( 
    .Z ( U623.AB ) ,
    .I0 ( masks_hold_reg_5_0 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U623.CD ) ,
    .I0 ( config1_xor_encoded_masks_64 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_64 ) ,
    .I0 ( U623.AB ) ,
    .I1 ( U623.CD ) ) ;
and ( 
    .Z ( U1173.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_41 ) ,
    .I1 ( n64 ) ) ;
and ( 
    .Z ( U1173.CD ) ,
    .I0 ( config0_onehot_decoded_masks_5_41 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1173.EF ) ,
    .I0 ( xor_decoded_masks_5_41 ) ,
    .I1 ( n17 ) ) ;
or ( 
    .Z ( masks_for_compactor_5_41 ) ,
    .I0 ( U1173.AB ) ,
    .I1 ( U1173.CD ) ,
    .I2 ( U1173.EF ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_9.DI_ ) ,
    .IN ( masks_shift_reg_1_9 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_9.CPI_ ) ,
    .IN ( CTS_lsi_ss_clk_delay2841 ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_reg_9.E_ ) ,
    .IN ( edt_update ) ) ;
buf ( 
    .O1 ( masks_hold_reg_1_9 ) ,
    .IN ( masks_hold_reg_1_reg_9.QT ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ,
    .A ( GND ) ) ;
buf ( 
    .Q ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ,
    .A ( GND ) ) ;
MUX21 masks_hold_reg_1_reg_9.SYNTEST_VL_LSI_MUX21_26796.I0 ( 
    .I0 ( masks_hold_reg_1_reg_9.QT ) ,
    .I1 ( masks_hold_reg_1_reg_9.DI_ ) ,
    .Q ( masks_hold_reg_1_reg_9.ED ) ,
    .S ( masks_hold_reg_1_reg_9.E_ ) ) ;
not ( 
    .O1 ( masks_hold_reg_1_reg_9.U6.CD_ ) ,
    .IN ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_22 ) ) ;
and ( 
    .Z ( masks_hold_reg_1_reg_9.U6.D_1 ) ,
    .I0 ( masks_hold_reg_1_reg_9.ED ) ,
    .I1 ( masks_hold_reg_1_reg_9.U6.CD_ ) ) ;
MUX21 masks_hold_reg_1_reg_9.U6.I2 ( 
    .I0 ( masks_hold_reg_1_reg_9.U6.D_1 ) ,
    .I1 ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_20 ) ,
    .Q ( masks_hold_reg_1_reg_9.U6.Q1 ) ,
    .S ( masks_hold_reg_1_reg_9.SYNTEST_EXP_ADDED_NET_21 ) ) ;
DFF masks_hold_reg_1_reg_9.U6.I3 ( 
    .CK ( masks_hold_reg_1_reg_9.CPI_ ) ,
    .D ( masks_hold_reg_1_reg_9.U6.Q1 ) ,
    .Q ( masks_hold_reg_1_reg_9.QT ) ) ;
and ( 
    .Z ( U709.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_118 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U709.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_11 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U709.EF ) ,
    .I0 ( xor_decoded_masks_2_11 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_11 ) ,
    .I0 ( U709.AB ) ,
    .I1 ( U709.CD ) ,
    .I2 ( U709.EF ) ) ;
and ( 
    .Z ( U622.AB ) ,
    .I0 ( masks_hold_reg_6_7 ) ,
    .I1 ( n44 ) ) ;
and ( 
    .Z ( U622.CD ) ,
    .I0 ( config1_xor_encoded_masks_68 ) ,
    .I1 ( n41 ) ) ;
or ( 
    .Z ( xor_encoded_masks_68 ) ,
    .I0 ( U622.AB ) ,
    .I1 ( U622.CD ) ) ;
and ( 
    .Z ( U1170.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_148 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U1170.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_41 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U1170.EF ) ,
    .I0 ( xor_decoded_masks_2_41 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_41 ) ,
    .I0 ( U1170.AB ) ,
    .I1 ( U1170.CD ) ,
    .I2 ( U1170.EF ) ) ;
and ( 
    .Z ( U625.AB ) ,
    .I0 ( masks_hold_reg_9_1 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U625.CD ) ,
    .I0 ( config1_xor_encoded_masks_107 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_107 ) ,
    .I0 ( U625.AB ) ,
    .I1 ( U625.CD ) ) ;
and ( 
    .Z ( U1171.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_41 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U1171.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_41 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U1171.EF ) ,
    .I0 ( xor_decoded_masks_3_41 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_41 ) ,
    .I0 ( U1171.AB ) ,
    .I1 ( U1171.CD ) ,
    .I2 ( U1171.EF ) ) ;
and ( 
    .Z ( U624.AB ) ,
    .I0 ( masks_hold_reg_11_3 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U624.CD ) ,
    .I0 ( config1_xor_encoded_masks_127 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_127 ) ,
    .I0 ( U624.AB ) ,
    .I1 ( U624.CD ) ) ;
and ( 
    .Z ( U1176.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_94 ) ,
    .I1 ( n56 ) ) ;
and ( 
    .Z ( U1176.CD ) ,
    .I0 ( config0_onehot_decoded_masks_8_41 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1176.EF ) ,
    .I0 ( xor_decoded_masks_8_41 ) ,
    .I1 ( n26 ) ) ;
or ( 
    .Z ( masks_for_compactor_8_41 ) ,
    .I0 ( U1176.AB ) ,
    .I1 ( U1176.CD ) ,
    .I2 ( U1176.EF ) ) ;
and ( 
    .Z ( U627.AB ) ,
    .I0 ( masks_hold_reg_9_3 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U627.CD ) ,
    .I0 ( config1_xor_encoded_masks_105 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_105 ) ,
    .I0 ( U627.AB ) ,
    .I1 ( U627.CD ) ) ;
and ( 
    .Z ( U1177.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_41 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1177.CD ) ,
    .I0 ( config0_onehot_decoded_masks_9_41 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1177.EF ) ,
    .I0 ( xor_decoded_masks_9_41 ) ,
    .I1 ( n27 ) ) ;
or ( 
    .Z ( masks_for_compactor_9_41 ) ,
    .I0 ( U1177.AB ) ,
    .I1 ( U1177.CD ) ,
    .I2 ( U1177.EF ) ) ;
and ( 
    .Z ( U626.AB ) ,
    .I0 ( masks_hold_reg_9_0 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U626.CD ) ,
    .I0 ( config1_xor_encoded_masks_108 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_108 ) ,
    .I0 ( U626.AB ) ,
    .I1 ( U626.CD ) ) ;
and ( 
    .Z ( U1174.AB ) ,
    .I0 ( config1_onehot_decoded_masks_2_94 ) ,
    .I1 ( n60 ) ) ;
and ( 
    .Z ( U1174.CD ) ,
    .I0 ( config0_onehot_decoded_masks_6_41 ) ,
    .I1 ( n71 ) ) ;
and ( 
    .Z ( U1174.EF ) ,
    .I0 ( xor_decoded_masks_6_41 ) ,
    .I1 ( n32 ) ) ;
or ( 
    .Z ( masks_for_compactor_6_41 ) ,
    .I0 ( U1174.AB ) ,
    .I1 ( U1174.CD ) ,
    .I2 ( U1174.EF ) ) ;
and ( 
    .Z ( U928.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_151 ) ,
    .I1 ( n57 ) ) ;
and ( 
    .Z ( U928.CD ) ,
    .I0 ( config0_onehot_decoded_masks_2_44 ) ,
    .I1 ( n75 ) ) ;
and ( 
    .Z ( U928.EF ) ,
    .I0 ( xor_decoded_masks_2_44 ) ,
    .I1 ( n21 ) ) ;
or ( 
    .Z ( masks_for_compactor_2_44 ) ,
    .I0 ( U928.AB ) ,
    .I1 ( U928.CD ) ,
    .I2 ( U928.EF ) ) ;
and ( 
    .Z ( U629.AB ) ,
    .I0 ( masks_hold_reg_11_1 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U629.CD ) ,
    .I0 ( config1_xor_encoded_masks_129 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_129 ) ,
    .I0 ( U629.AB ) ,
    .I1 ( U629.CD ) ) ;
and ( 
    .Z ( U1175.AB ) ,
    .I0 ( config1_onehot_decoded_masks_3_41 ) ,
    .I1 ( n61 ) ) ;
and ( 
    .Z ( U1175.CD ) ,
    .I0 ( config0_onehot_decoded_masks_7_41 ) ,
    .I1 ( n72 ) ) ;
and ( 
    .Z ( U1175.EF ) ,
    .I0 ( xor_decoded_masks_7_41 ) ,
    .I1 ( n25 ) ) ;
or ( 
    .Z ( masks_for_compactor_7_41 ) ,
    .I0 ( U1175.AB ) ,
    .I1 ( U1175.CD ) ,
    .I2 ( U1175.EF ) ) ;
and ( 
    .Z ( U929.AB ) ,
    .I0 ( config1_onehot_decoded_masks_1_44 ) ,
    .I1 ( n63 ) ) ;
and ( 
    .Z ( U929.CD ) ,
    .I0 ( config0_onehot_decoded_masks_3_44 ) ,
    .I1 ( n76 ) ) ;
and ( 
    .Z ( U929.EF ) ,
    .I0 ( xor_decoded_masks_3_44 ) ,
    .I1 ( n19 ) ) ;
or ( 
    .Z ( masks_for_compactor_3_44 ) ,
    .I0 ( U929.AB ) ,
    .I1 ( U929.CD ) ,
    .I2 ( U929.EF ) ) ;
and ( 
    .Z ( U628.AB ) ,
    .I0 ( masks_hold_reg_11_8 ) ,
    .I1 ( n45 ) ) ;
and ( 
    .Z ( U628.CD ) ,
    .I0 ( config1_xor_encoded_masks_122 ) ,
    .I1 ( edt_configuration_hfs_netlink_29290 ) ) ;
or ( 
    .Z ( xor_encoded_masks_122 ) ,
    .I0 ( U628.AB ) ,
    .I1 ( U628.CD ) ) ;
and ( 
    .Z ( U926.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_30 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U926.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_30 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U926.EF ) ,
    .I0 ( xor_decoded_masks_0_30 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_30 ) ,
    .I0 ( U926.AB ) ,
    .I1 ( U926.CD ) ,
    .I2 ( U926.EF ) ) ;
and ( 
    .Z ( U927.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_26 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U927.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_26 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U927.EF ) ,
    .I0 ( xor_decoded_masks_0_26 ) ,
    .I1 ( n23 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_26 ) ,
    .I0 ( U927.AB ) ,
    .I1 ( U927.CD ) ,
    .I2 ( U927.EF ) ) ;
and ( 
    .Z ( U863.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_21 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U863.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_21 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U863.EF ) ,
    .I0 ( xor_decoded_masks_0_21 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_21 ) ,
    .I0 ( U863.AB ) ,
    .I1 ( U863.CD ) ,
    .I2 ( U863.EF ) ) ;
and ( 
    .Z ( U1178.AB ) ,
    .I0 ( config1_onehot_decoded_masks_4_94 ) ,
    .I1 ( n59 ) ) ;
and ( 
    .Z ( U1178.CD ) ,
    .I0 ( config0_onehot_decoded_masks_10_41 ) ,
    .I1 ( n70 ) ) ;
and ( 
    .Z ( U1178.EF ) ,
    .I0 ( xor_decoded_masks_10_41 ) ,
    .I1 ( n28 ) ) ;
or ( 
    .Z ( masks_for_compactor_10_41 ) ,
    .I0 ( U1178.AB ) ,
    .I1 ( U1178.CD ) ,
    .I2 ( U1178.EF ) ) ;
and ( 
    .Z ( U849.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_44 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U849.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_44 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U849.EF ) ,
    .I0 ( xor_decoded_masks_11_44 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_44 ) ,
    .I0 ( U849.AB ) ,
    .I1 ( U849.CD ) ,
    .I2 ( U849.EF ) ) ;
and ( 
    .Z ( U1288.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_103 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1288.CD ) ,
    .I0 ( config0_onehot_decoded_masks_12_50 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1288.EF ) ,
    .I0 ( xor_decoded_masks_12_50 ) ,
    .I1 ( n34 ) ) ;
or ( 
    .Z ( masks_for_compactor_12_50 ) ,
    .I0 ( U1288.AB ) ,
    .I1 ( U1288.CD ) ,
    .I2 ( U1288.EF ) ) ;
and ( 
    .Z ( U924.AB ) ,
    .I0 ( config1_onehot_decoded_masks_0_22 ) ,
    .I1 ( n65 ) ) ;
and ( 
    .Z ( U924.CD ) ,
    .I0 ( config0_onehot_decoded_masks_0_22 ) ,
    .I1 ( n74 ) ) ;
and ( 
    .Z ( U924.EF ) ,
    .I0 ( xor_decoded_masks_0_22 ) ,
    .I1 ( n22 ) ) ;
or ( 
    .Z ( masks_for_compactor_0_22 ) ,
    .I0 ( U924.AB ) ,
    .I1 ( U924.CD ) ,
    .I2 ( U924.EF ) ) ;
and ( 
    .Z ( U1179.AB ) ,
    .I0 ( config1_onehot_decoded_masks_5_41 ) ,
    .I1 ( n62 ) ) ;
and ( 
    .Z ( U1179.CD ) ,
    .I0 ( config0_onehot_decoded_masks_11_41 ) ,
    .I1 ( n73 ) ) ;
and ( 
    .Z ( U1179.EF ) ,
    .I0 ( xor_decoded_masks_11_41 ) ,
    .I1 ( n33 ) ) ;
or ( 
    .Z ( masks_for_compactor_11_41 ) ,
    .I0 ( U1179.AB ) ,
    .I1 ( U1179.CD ) ,
    .I2 ( U1179.EF ) ) ;
buf ( 
    .O1 ( n42 ) ,
    .IN ( masks_shift_reg_12_8 ) ) ;
buf ( 
    .O1 ( n46 ) ,
    .IN ( masks_shift_reg_12_7 ) ) ;
buf ( 
    .O1 ( n67 ) ,
    .IN ( masks_shift_reg_12_9 ) ) ;
buf ( 
    .O1 ( n79 ) ,
    .IN ( masks_hold_reg_2_6 ) ) ;
buf ( 
    .O1 ( n86 ) ,
    .IN ( n79 ) ) ;
buf ( 
    .O1 ( n90 ) ,
    .IN ( masks_hold_reg_3_5 ) ) ;
buf ( 
    .O1 ( n91 ) ,
    .IN ( masks_hold_reg_3_2 ) ) ;
buf ( 
    .O1 ( n92 ) ,
    .IN ( masks_hold_reg_4_9 ) ) ;
buf ( 
    .O1 ( n93 ) ,
    .IN ( masks_shift_reg_8_8 ) ) ;
buf ( 
    .O1 ( n94 ) ,
    .IN ( masks_shift_reg_4_9 ) ) ;
buf ( 
    .O1 ( n95 ) ,
    .IN ( masks_shift_reg_6_6 ) ) ;
buf ( 
    .O1 ( n96 ) ,
    .IN ( masks_shift_reg_9_4 ) ) ;
buf ( 
    .O1 ( n97 ) ,
    .IN ( masks_shift_reg_2_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I9 ) ,
    .IN ( edt_clock_cts_6_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I11 ) ,
    .IN ( edt_clock_cts_7_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I3 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I23 ) ,
    .IN ( edt_clock_cts_6_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I24 ) ,
    .IN ( edt_clock_cts_6_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I27 ) ,
    .IN ( edt_clock_cts_6_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I25 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I34 ) ,
    .IN ( edt_clock_cts_6_1 ) ) ;
not ( 
    .O1 ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I1 ) ,
    .IN ( edt_clock_cts_5_1 ) ) ;
not ( 
    .O1 ( n44 ) ,
    .IN ( n41 ) ) ;
not ( 
    .O1 ( n38 ) ,
    .IN ( n37 ) ) ;
not ( 
    .O1 ( n43 ) ,
    .IN ( n40 ) ) ;
not ( 
    .O1 ( n29 ) ,
    .IN ( n5 ) ) ;
buf ( 
    .O1 ( n49 ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
not ( 
    .O1 ( n22 ) ,
    .IN ( n4 ) ) ;
buf ( 
    .O1 ( n37 ) ,
    .IN ( edt_configuration ) ) ;
not ( 
    .O1 ( n53 ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
not ( 
    .O1 ( n52 ) ,
    .IN ( edt_update_hfs_netlink_29280 ) ) ;
not ( 
    .O1 ( n17 ) ,
    .IN ( n4 ) ) ;
buf ( 
    .O1 ( n4 ) ,
    .IN ( n3 ) ) ;
not ( 
    .O1 ( n48 ) ,
    .IN ( n47 ) ) ;
not ( 
    .O1 ( n19 ) ,
    .IN ( n4 ) ) ;
buf ( 
    .O1 ( n47 ) ,
    .IN ( edt_update ) ) ;
not ( 
    .O1 ( n34 ) ,
    .IN ( n5 ) ) ;
buf ( 
    .O1 ( n40 ) ,
    .IN ( edt_configuration_hfs_netlink_29290 ) ) ;
buf ( 
    .O1 ( n41 ) ,
    .IN ( edt_configuration_hfs_netlink_29290 ) ) ;
buf ( 
    .O1 ( n56 ) ,
    .IN ( n55 ) ) ;
buf ( 
    .O1 ( n68 ) ,
    .IN ( n2 ) ) ;
buf ( 
    .O1 ( n5 ) ,
    .IN ( n3 ) ) ;
not ( 
    .O1 ( n51 ) ,
    .IN ( n49 ) ) ;
not ( 
    .O1 ( n54 ) ,
    .IN ( edt_update_hfs_netlink_29281 ) ) ;
not ( 
    .O1 ( n25 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n23 ) ,
    .IN ( n4 ) ) ;
not ( 
    .O1 ( n21 ) ,
    .IN ( n4 ) ) ;
not ( 
    .O1 ( n30 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n28 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n27 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n33 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n32 ) ,
    .IN ( n5 ) ) ;
not ( 
    .O1 ( n31 ) ,
    .IN ( n5 ) ) ;
buf ( 
    .O1 ( n60 ) ,
    .IN ( n56 ) ) ;
buf ( 
    .O1 ( n75 ) ,
    .IN ( n68 ) ) ;
buf ( 
    .O1 ( n71 ) ,
    .IN ( n66 ) ) ;
not ( 
    .O1 ( n26 ) ,
    .IN ( n5 ) ) ;
buf ( 
    .O1 ( n58 ) ,
    .IN ( n56 ) ) ;
buf ( 
    .O1 ( n72 ) ,
    .IN ( n66 ) ) ;
buf ( 
    .O1 ( n73 ) ,
    .IN ( n66 ) ) ;
buf ( 
    .O1 ( n59 ) ,
    .IN ( n56 ) ) ;
buf ( 
    .O1 ( n69 ) ,
    .IN ( n66 ) ) ;
buf ( 
    .O1 ( n70 ) ,
    .IN ( n66 ) ) ;
buf ( 
    .O1 ( n61 ) ,
    .IN ( n56 ) ) ;
buf ( 
    .O1 ( n62 ) ,
    .IN ( n56 ) ) ;
buf ( 
    .O1 ( n76 ) ,
    .IN ( n68 ) ) ;
buf ( 
    .O1 ( n74 ) ,
    .IN ( n68 ) ) ;
not ( 
    .O1 ( n45 ) ,
    .IN ( edt_configuration_hfs_netlink_29290 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2841 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I9 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2881 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I3 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2861 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I11 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2781 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I24 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2641 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I27 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay2961 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I23 ) ) ;
buf ( 
    .O1 ( CTS_lsi_ss_clk_delay1941 ) ,
    .IN ( net_LSI_EDT_CLOCK_power_clock_gate_G2B2I34 ) ) ;
buf ( 
    .O1 ( n2 ) ,
    .IN ( n66 ) ) ;
buf ( 
    .O1 ( n1 ) ,
    .IN ( n55 ) ) ;
endmodule

