module mtx_top(CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G487,G500,G513,G526,G539,G552,G565,G578,G591,G604,G617,G1289,G1310,G1331,G1352,G1373,G1394,G1415,G1436,G1497,G1518,G1539,G1560,G1581,G1602,G1623,G1644,G1705,G1726,G1747,G1768,G1789,G1810,G1831,G1852,G1913,G1934,G1955,G1976,G1997,G2018,G2039,G2060,G2121,G2142,G2163,G2184,G2205,G2226,G2247,G2268,G2329,G2350,G2371,G2392,G2413,G2434,G2455,G2476,G2537,G2558,G2579,G2600,G2621,G2642,G2663,G2684,G2745,G2766,G2787,G2808,G2829,G2850,G2871,G2892,G2953,G2974,G2995,G3016,G3037,G3058,G3079,G3100,G3161,G3182,G3203,G3224,G3245,G3266,G3287,G3308,G3369,G3390,G3411,G3432,G3453,G3474,G3495,G3516,G3537,G3598,G3619,G3640,G3661,G3682,G3703,G3724,G3745,G3806,G3827,G3848,G3869,G3890,G3911,G3932,G3953,G4014,G4035,G4056,G4077,G4098,G4119,G4140,G4161,G4222,G4243,G4264,G4285,G4306,G4327,G4348,G4369,G4390,G4451,G4472,G4493,G4514,G4535,G4556,G4577,G4598,G4659,G4680,G4701,G4722,G4743,G4764,G4785,G4806,G4867,G4888,G4909,G4930,G4951,G4972,G4993,G5014,G5075,G5096,G5117,G5138,G5159,G5180,G5201,G5222,G5243,G5304,G5325,G5346,G5367,G5388,G5409,G5430,G5451,G5512,G5533,G5554,G5575,G5596,G5617,G5638,G5659,G5720,G5741,G5762,G5783,G5804,G5825,G5846,G5867,G5928,G5949,G5970,G5991,G6012,G6033,G6054,G6075,G6136,G6157,G6178,G6199,G6220,G6241,G6262,G6283,G6344,G6365,G6386,G6407,G6428,G6449,G6470,G6491,G6552,G6573,G6594,G6615,G6636,G6657,G6678,G6699,G6760,G6781,G6802,G6823,G6844,G6865,G6886,G6907,G6968,G6989,G7010,G7031,G7052,G7073,G7094,G7115,G7176,G7197,G7218,G7239,G7260,G7281,G7302,G7323,G7384,G7405,G7426,G7447,G7468,G7489,G7510,G7531,G7592,G7613,G7634,G7655,G7676,G7697,G7718,G7739,G7800,G7821,G7842,G7863,G7884,G7905,G7926,G7947,G8008,G8029,G8050,G8071,G8092,G8113,G8134,G8155,G8216,G8237,G8258,G8279,G8300,G8321,G8342,G8363,G8424,G8445,G8466,G8487,G8508,G8529,G8550,G8571,G8632,G8653,G8674,G8695,G8716,G8737,G8758,G8779,G8840,G8861,G8882,G8903,G8924,G8945,G8966,G8987,G9048,G9069,G9090,G9111,G9132,G9153,G9174,G9195,G9256,G9277,G9298,G9319,G9340,G9361,G9382,G9403,G9464,G9485,G9506,G9527,G9548,G9569,G9590,G9611,G9672,G9693,G9714,G9735,G9756,G9777,G9798,G9819,G9880,G9901,G9922,G9943,G9964,G9985,G10006,G10027,G10088,G10109,G10130,G10151,G10172,G10193,G10214,G10235,G10296,G10317,G10338,G10359,G10380,G10401,G10422,G10443,G10504,G10525,G10546,G10567,G10588,G10609,G10630,G10651,G10712,G10733,G10754,G10775,G10796,G10817,G10838,G10859,G11327,G11348,G11369,G11390,G11411,G11432,G11453,G11475,G31621,G31634,G31647,G31660,G31673,G31686,G31699,G31712,G31725,G31738,G31751,G31764,G31777,G31790,G31803,G31816,G31829,G31842,G31855,G31868,G31881,G31894,G31907,G31920,G31933,G31946,G31959,G31972,G31985,G31998,G32011,G32024,G32037,G32050,G32063,G32076,G32089,G32102,G32115,G32128,G32141,G32154,G32167,G32180,G32193,G32206,G32219,G32232,G32245,G32258,G32271,G32284,G32297,G32310,G32323,G32336,G32349,G32362,G32375,G32388,G32401,G32414,G32427,G32440,G32453,G32466,G32479,G32492,G32505,G32518,G32531,G32544,G32557,G32570,G32583,G32596,G32609,G32622,G32635,G32648,G32661,G32674,G32687,G32700,G32713,G32726,G32739,G32752,G32765,G32778,G32791,G32804,G32817,G32830,G32843,G32856,G32869,G32882,G32895,G32908,G32921,G32934,G32947,G32960,G32973,G32986,G32999,G33012,G33025,G33038,G33051,G33064,G33077,G33090,G33103,G33116,G33129,G33142,G33155,G33168,G33181,G33194,G33207,G33220,G33233,G33246,G33259,G33272,G33285,G33298,G33311,G33324,G33337,G33350,G33363,G33376,G33389,G33402,G33415,G33428,G33441,G33454,G33467,G33480,G33493,G33506,G33519,G33532,G33545,G33558,G33571,G33584,G33597,G33610,G33623,G33636,G33649,G33662,G33675,G33688,G33701,G33714,G33727,G33740,G33753,G33766,G33779,G33792,G33805,G33818,G33831,G33844,G33857,G33870,G33883,G33896,G33909,G33922,G33935,G33948,G33961,G33974,G33987,G34000,G34013,G34026,G34039,G34052,G34065,G34078,G34091,G34104,G34117,G34130,G34143,G34156,G34169,G34182,G34195,G34208,G34221,G34234,G34247,G34260,G34273,G34286,G34299,G34312,G34325,G34338,G34351,G34364,G34377,G34390,G34403,G34416,G34429,G34442,G34455,G34468,G34481,G34494,G34507,G34520,G34533,G34546,G34559,G34572,G34585,G54748,G54761,G54774,G54787,G54800,G54813,G54826,G54839,G54852,G54865,G54878,G54891,G54904,G54917,G54930,G54943,G54956,G54969,G54982,G54995,G55008,G55021,G55034,G55047,G55060,G55073,G55086,G55099,G55112,G55125,G55138,G55151,G55164,G55177,G55190,G55203,G55216,G55229,G55242,G55255,G55268,G55281,G55294,G55307,G55320,G55333,G55346,G55359,G55372,G55385,G55398,G55411,G55424,G55437,G55450,G55463,G55476,G55489,G55502,G55515,G55528,G55541,G55554,G55567,G55580,G55593,G55606,G55619,G55632,G55645,G55658,G55671,G55684,G55697,G55710,G55723,G55736,G55749,G55762,G55775,G55788,G55801,G55814,G55827,G55840,G55853,G55866,G55879,G55892,G55905,G55918,G55931,G55944,G55957,G55970,G55983,G55996,G56009,G56022,G56035,G56048,G56061,G56074,G56087,G56100,G56113,G56126,G56139,G56152,G56165,G56178,G56191,G56204,G56217,G56230,G56243,G56256,G56269,G56282,G56295,G56308,G56321,G56334,G56347,G56360,G56373,G56386,G56399,G56412,G56425,G56438,G56451,G56464,G56477,G56490,G56503,G56516,G56529,G56542,G56555,G56568,G56581,G56594,G56607,G56620,G56633,G56646,G56659,G56672,G56685,G56698,G56711,G56724,G56737,G56750,G56763,G56776,G56789,G56802,G56815,G56828,G56841,G56854,G56867,G56880,G56893,G56906,G56919,G56932,G56945,G56958,G56971,G56984,G56997,G57010,G57023,G57036,G57049,G57062,G57075,G57088,G57101,G57114,G57127,G57140,G57153,G57166,G57179,G57192,G57205,G57218,G57231,G57244,G57257,G57270,G57283,G57296,G57309,G57322,G57335,G57348,G57361,G57374,G57387,G57400,G57413,G57426,G57439,G57452,G57465,G57478,G57491,G57504,G57517,G57530,G57543,G57556,G57569,G57582,G57595,G57608,G57621,G57634,G57647,G57660,G57673,G57686,G57699,G57712,G77875,G77888,G77901,G77914,G77927,G77940,G77953,G77966,G77979,G77992,G78005,G78018,G78031,G78044,G78057,G78070,G78083,G78096,G78109,G78122,G78135,G78148,G78161,G78174,G78187,G78200,G78213,G78226,G78239,G78252,G78265,G78278,G78291,G78304,G78317,G78330,G78343,G78356,G78369,G78382,G78395,G78408,G78421,G78434,G78447,G78460,G78473,G78486,G78499,G78512,G78525,G78538,G78551,G78564,G78577,G78590,G78603,G78616,G78629,G78642,G78655,G78668,G78681,G78694,G78707,G78720,G78733,G78746,G78759,G78772,G78785,G78798,G78811,G78824,G78837,G78850,G78863,G78876,G78889,G78902,G78915,G78928,G78941,G78954,G78967,G78980,G78993,G79006,G79019,G79032,G79045,G79058,G79071,G79084,G79097,G79110,G79123,G79136,G79149,G79162,G79175,G79188,G79201,G79214,G79227,G79240,G79253,G79266,G79279,G79292,G79305,G79318,G79331,G79344,G79357,G79370,G79383,G79396,G79409,G79422,G79435,G79448,G79461,G79474,G79487,G79500,G79513,G79526,G79539,G79552,G79565,G79578,G79591,G79604,G79617,G79630,G79643,G79656,G79669,G79682,G79695,G79708,G79721,G79734,G79747,G79760,G79773,G79786,G79799,G79812,G79825,G79838,G79851,G79864,G79877,G79890,G79903,G79916,G79929,G79942,G79955,G79968,G79981,G79994,G80007,G80020,G80033,G80046,G80059,G80072,G80085,G80098,G80111,G80124,G80137,G80150,G80163,G80176,G80189,G80202,G80215,G80228,G80241,G80254,G80267,G80280,G80293,G80306,G80319,G80332,G80345,G80358,G80371,G80384,G80397,G80410,G80423,G80436,G80449,G80462,G80475,G80488,G80501,G80514,G80527,G80540,G80553,G80566,G80579,G80592,G80605,G80618,G80631,G80644,G80657,G80670,G80683,G80696,G80709,G80722,G80735,G80748,G80761,G80774,G80787,G80800,G80813,G80826,G80839,G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G109,G110,G112,G114,G116,G118,G120,G122,G124,G126,G128,G130,G132,G134,G136,G138,G140,G142,G144,G146,G496,G509,G522,G535,G548,G561,G574,G587,G600,G613,G1306,G1327,G1348,G1369,G1390,G1411,G1432,G1453,G1514,G1535,G1556,G1577,G1598,G1619,G1640,G1661,G1722,G1743,G1764,G1785,G1806,G1827,G1848,G1869,G1930,G1951,G1972,G1993,G2014,G2035,G2056,G2077,G2138,G2159,G2180,G2201,G2222,G2243,G2264,G2285,G2346,G2367,G2388,G2409,G2430,G2451,G2472,G2493,G2554,G2575,G2596,G2617,G2638,G2659,G2680,G2701,G2762,G2783,G2804,G2825,G2846,G2867,G2888,G2909,G2970,G2991,G3012,G3033,G3054,G3075,G3096,G3117,G3178,G3199,G3220,G3241,G3262,G3283,G3304,G3325,G3386,G3407,G3428,G3449,G3470,G3491,G3512,G3533,G3554,G3615,G3636,G3657,G3678,G3699,G3720,G3741,G3762,G3823,G3844,G3865,G3886,G3907,G3928,G3949,G3970,G4031,G4052,G4073,G4094,G4115,G4136,G4157,G4178,G4239,G4260,G4281,G4302,G4323,G4344,G4365,G4386,G4407,G4468,G4489,G4510,G4531,G4552,G4573,G4594,G4615,G4676,G4697,G4718,G4739,G4760,G4781,G4802,G4823,G4884,G4905,G4926,G4947,G4968,G4989,G5010,G5031,G5092,G5113,G5134,G5155,G5176,G5197,G5239,G5260,G5321,G5342,G5363,G5384,G5405,G5426,G5447,G5468,G5529,G5550,G5571,G5592,G5613,G5634,G5655,G5676,G5737,G5758,G5779,G5800,G5821,G5842,G5863,G5884,G5945,G5966,G5987,G6008,G6029,G6050,G6071,G6092,G6153,G6174,G6195,G6216,G6237,G6258,G6279,G6300,G6361,G6382,G6403,G6424,G6445,G6466,G6487,G6508,G6569,G6590,G6611,G6632,G6653,G6674,G6695,G6716,G6777,G6798,G6819,G6840,G6861,G6882,G6903,G6924,G6985,G7006,G7027,G7048,G7069,G7090,G7111,G7132,G7193,G7214,G7235,G7256,G7277,G7298,G7319,G7340,G7401,G7422,G7443,G7464,G7485,G7506,G7527,G7548,G7609,G7630,G7651,G7672,G7693,G7714,G7735,G7756,G7817,G7838,G7859,G7880,G7901,G7922,G7943,G7964,G8025,G8046,G8067,G8088,G8109,G8130,G8151,G8172,G8233,G8254,G8275,G8296,G8317,G8338,G8359,G8380,G8441,G8462,G8483,G8504,G8525,G8546,G8567,G8588,G8649,G8691,G8712,G8733,G8754,G8775,G8796,G8857,G8878,G8899,G8920,G8941,G8962,G8983,G9004,G9065,G9086,G9107,G9128,G9149,G9170,G9191,G9212,G9273,G9294,G9315,G9336,G9357,G9378,G9399,G9420,G9481,G9502,G9523,G9544,G9565,G9586,G9607,G9628,G9689,G9710,G9731,G9752,G9773,G9794,G9815,G9836,G9897,G9918,G9939,G9960,G9981,G10002,G10023,G10044,G10105,G10126,G10147,G10168,G10189,G10210,G10231,G10252,G10313,G10334,G10355,G10376,G10397,G10418,G10439,G10460,G10521,G10542,G10563,G10584,G10605,G10626,G10647,G10668,G10729,G10750,G10771,G10792,G10813,G10834,G10855,G10876,G11344,G11365,G11386,G11407,G11428,G11449,G11470,G11492,G31630,G31643,G31656,G31669,G31682,G31695,G31708,G31721,G31734,G31747,G31760,G31773,G31786,G31799,G31812,G31825,G31838,G31851,G31864,G31877,G31890,G31903,G31916,G31929,G31942,G31955,G31968,G31981,G31994,G32007,G32020,G32033,G32046,G32059,G32072,G32085,G32098,G32111,G32124,G32137,G32150,G32163,G32176,G32189,G32202,G32215,G32228,G32241,G32254,G32267,G32280,G32293,G32306,G32319,G32332,G32345,G32358,G32371,G32384,G32397,G32410,G32423,G32436,G32449,G32462,G32475,G32488,G32501,G32514,G32527,G32540,G32553,G32566,G32579,G32592,G32605,G32618,G32631,G32644,G32657,G32670,G32683,G32696,G32709,G32722,G32735,G32748,G32761,G32774,G32787,G32800,G32813,G32826,G32839,G32852,G32865,G32878,G32891,G32904,G32917,G32930,G32943,G32956,G32969,G32982,G32995,G33008,G33021,G33034,G33047,G33060,G33073,G33086,G33099,G33112,G33125,G33138,G33151,G33164,G33177,G33190,G33203,G33216,G33229,G33242,G33255,G33268,G33281,G33294,G33307,G33320,G33333,G33346,G33359,G33372,G33385,G33398,G33411,G33424,G33437,G33450,G33463,G33476,G33489,G33502,G33515,G33528,G33541,G33554,G33567,G33580,G33593,G33606,G33619,G33632,G33645,G33658,G33671,G33684,G33697,G33710,G33723,G33736,G33749,G33762,G33775,G33788,G33801,G33814,G33827,G33840,G33853,G33866,G33879,G33892,G33905,G33918,G33931,G33944,G33957,G33970,G33983,G33996,G34009,G34022,G34035,G34048,G34061,G34074,G34087,G34100,G34113,G34126,G34139,G34152,G34165,G34178,G34191,G34204,G34217,G34230,G34243,G34256,G34269,G34282,G34295,G34308,G34321,G34334,G34347,G34373,G34386,G34399,G34412,G34425,G34438,G34451,G34464,G34477,G34490,G34503,G34516,G34529,G34542,G34555,G34568,G34581,G54757,G54770,G54783,G54796,G54809,G54822,G54835,G54848,G54861,G54874,G54887,G54900,G54913,G54926,G54939,G54952,G54965,G54978,G54991,G55004,G55017,G55030,G55043,G55056,G55069,G55082,G55095,G55108,G55121,G55134,G55147,G55160,G55173,G55186,G55199,G55212,G55225,G55238,G55251,G55264,G55277,G55290,G55303,G55316,G55329,G55342,G55355,G55368,G55381,G55394,G55407,G55420,G55433,G55446,G55459,G55472,G55485,G55498,G55511,G55524,G55537,G55550,G55563,G55576,G55589,G55602,G55615,G55628,G55641,G55654,G55667,G55680,G55693,G55706,G55719,G55732,G55745,G55758,G55771,G55784,G55797,G55810,G55823,G55836,G55849,G55862,G55875,G55888,G55901,G55914,G55927,G55940,G55953,G55966,G55979,G55992,G56005,G56018,G56031,G56044,G56057,G56070,G56083,G56096,G56109,G56122,G56135,G56148,G56161,G56174,G56187,G56200,G56213,G56226,G56239,G56252,G56265,G56278,G56291,G56304,G56317,G56330,G56343,G56356,G56369,G56382,G56395,G56408,G56421,G56434,G56447,G56460,G56473,G56486,G56499,G56512,G56525,G56538,G56551,G56564,G56577,G56590,G56603,G56616,G56629,G56642,G56655,G56668,G56681,G56694,G56707,G56720,G56733,G56746,G56759,G56772,G56785,G56798,G56811,G56824,G56837,G56850,G56863,G56876,G56889,G56902,G56915,G56928,G56941,G56954,G56967,G56980,G56993,G57006,G57019,G57032,G57045,G57058,G57071,G57084,G57097,G57110,G57123,G57136,G57149,G57162,G57175,G57188,G57201,G57214,G57227,G57240,G57253,G57266,G57279,G57292,G57305,G57318,G57331,G57357,G57370,G57383,G57396,G57409,G57422,G57435,G57448,G57461,G57474,G57487,G57500,G57513,G57526,G57539,G57552,G57578,G57591,G57604,G57617,G57630,G57643,G57656,G57669,G57682,G57695,G57708,G57721,G77884,G77897,G77910,G77923,G77936,G77949,G77962,G77975,G77988,G78001,G78014,G78027,G78040,G78053,G78066,G78079,G78092,G78105,G78118,G78131,G78144,G78157,G78170,G78183,G78196,G78209,G78222,G78235,G78248,G78261,G78274,G78287,G78300,G78313,G78326,G78339,G78352,G78365,G78378,G78391,G78404,G78417,G78430,G78443,G78456,G78469,G78482,G78495,G78508,G78521,G78534,G78547,G78560,G78573,G78586,G78599,G78612,G78625,G78638,G78651,G78664,G78677,G78690,G78703,G78716,G78729,G78742,G78755,G78768,G78781,G78794,G78807,G78820,G78833,G78846,G78859,G78872,G78885,G78898,G78911,G78924,G78937,G78950,G78963,G78976,G78989,G79002,G79015,G79028,G79041,G79054,G79067,G79080,G79093,G79106,G79119,G79132,G79145,G79158,G79171,G79184,G79197,G79210,G79223,G79236,G79249,G79262,G79275,G79288,G79301,G79314,G79327,G79340,G79353,G79366,G79379,G79392,G79405,G79418,G79431,G79444,G79457,G79470,G79483,G79496,G79509,G79522,G79535,G79548,G79561,G79574,G79587,G79600,G79613,G79626,G79639,G79652,G79665,G79678,G79691,G79704,G79717,G79730,G79743,G79756,G79769,G79782,G79795,G79808,G79821,G79834,G79847,G79860,G79873,G79886,G79899,G79912,G79925,G79938,G79951,G79964,G79977,G79990,G80003,G80016,G80029,G80042,G80055,G80068,G80081,G80094,G80107,G80120,G80133,G80146,G80159,G80172,G80185,G80211,G80224,G80237,G80250,G80263,G80276,G80289,G80302,G80315,G80328,G80341,G80354,G80367,G80380,G80393,G80406,G80419,G80432,G80445,G80458,G80471,G80484,G80497,G80510,G80523,G80536,G80549,G80562,G80575,G80588,G80601,G80614,G80627,G80640,G80653,G80679,G80692,G80705,G80731,G80744,G80757,G80770,G80783,G80796,G80809,G80822,G80835,G80848);
input CK,G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G487,G500,G513,G526,G539,G552,G565,G578,G591,G604,G617,G1289,G1310,G1331,G1352,G1373,G1394,G1415,G1436,G1497,G1518,G1539,G1560,G1581,G1602,G1623,G1644,G1705,G1726,G1747,G1768,G1789,G1810,G1831,G1852,G1913,G1934,G1955,G1976,G1997,G2018,G2039,G2060,G2121,G2142,G2163,G2184,G2205,G2226,G2247,G2268,G2329,G2350,G2371,G2392,G2413,G2434,G2455,G2476,G2537,G2558,G2579,G2600,G2621,G2642,G2663,G2684,G2745,G2766,G2787,G2808,G2829,G2850,G2871,G2892,G2953,G2974,G2995,G3016,G3037,G3058,G3079,G3100,G3161,G3182,G3203,G3224,G3245,G3266,G3287,G3308,G3369,G3390,G3411,G3432,G3453,G3474,G3495,G3516,G3537,G3598,G3619,G3640,G3661,G3682,G3703,G3724,G3745,G3806,G3827,G3848,G3869,G3890,G3911,G3932,G3953,G4014,G4035,G4056,G4077,G4098,G4119,G4140,G4161,G4222,G4243,G4264,G4285,G4306,G4327,G4348,G4369,G4390,G4451,G4472,G4493,G4514,G4535,G4556,G4577,G4598,G4659,G4680,G4701,G4722,G4743,G4764,G4785,G4806,G4867,G4888,G4909,G4930,G4951,G4972,G4993,G5014,G5075,G5096,G5117,G5138,G5159,G5180,G5201,G5222,G5243,G5304,G5325,G5346,G5367,G5388,G5409,G5430,G5451,G5512,G5533,G5554,G5575,G5596,G5617,G5638,G5659,G5720,G5741,G5762,G5783,G5804,G5825,G5846,G5867,G5928,G5949,G5970,G5991,G6012,G6033,G6054,G6075,G6136,G6157,G6178,G6199,G6220,G6241,G6262,G6283,G6344,G6365,G6386,G6407,G6428,G6449,G6470,G6491,G6552,G6573,G6594,G6615,G6636,G6657,G6678,G6699,G6760,G6781,G6802,G6823,G6844,G6865,G6886,G6907,G6968,G6989,G7010,G7031,G7052,G7073,G7094,G7115,G7176,G7197,G7218,G7239,G7260,G7281,G7302,G7323,G7384,G7405,G7426,G7447,G7468,G7489,G7510,G7531,G7592,G7613,G7634,G7655,G7676,G7697,G7718,G7739,G7800,G7821,G7842,G7863,G7884,G7905,G7926,G7947,G8008,G8029,G8050,G8071,G8092,G8113,G8134,G8155,G8216,G8237,G8258,G8279,G8300,G8321,G8342,G8363,G8424,G8445,G8466,G8487,G8508,G8529,G8550,G8571,G8632,G8653,G8674,G8695,G8716,G8737,G8758,G8779,G8840,G8861,G8882,G8903,G8924,G8945,G8966,G8987,G9048,G9069,G9090,G9111,G9132,G9153,G9174,G9195,G9256,G9277,G9298,G9319,G9340,G9361,G9382,G9403,G9464,G9485,G9506,G9527,G9548,G9569,G9590,G9611,G9672,G9693,G9714,G9735,G9756,G9777,G9798,G9819,G9880,G9901,G9922,G9943,G9964,G9985,G10006,G10027,G10088,G10109,G10130,G10151,G10172,G10193,G10214,G10235,G10296,G10317,G10338,G10359,G10380,G10401,G10422,G10443,G10504,G10525,G10546,G10567,G10588,G10609,G10630,G10651,G10712,G10733,G10754,G10775,G10796,G10817,G10838,G10859,G11327,G11348,G11369,G11390,G11411,G11432,G11453,G11475,G31621,G31634,G31647,G31660,G31673,G31686,G31699,G31712,G31725,G31738,G31751,G31764,G31777,G31790,G31803,G31816,G31829,G31842,G31855,G31868,G31881,G31894,G31907,G31920,G31933,G31946,G31959,G31972,G31985,G31998,G32011,G32024,G32037,G32050,G32063,G32076,G32089,G32102,G32115,G32128,G32141,G32154,G32167,G32180,G32193,G32206,G32219,G32232,G32245,G32258,G32271,G32284,G32297,G32310,G32323,G32336,G32349,G32362,G32375,G32388,G32401,G32414,G32427,G32440,G32453,G32466,G32479,G32492,G32505,G32518,G32531,G32544,G32557,G32570,G32583,G32596,G32609,G32622,G32635,G32648,G32661,G32674,G32687,G32700,G32713,G32726,G32739,G32752,G32765,G32778,G32791,G32804,G32817,G32830,G32843,G32856,G32869,G32882,G32895,G32908,G32921,G32934,G32947,G32960,G32973,G32986,G32999,G33012,G33025,G33038,G33051,G33064,G33077,G33090,G33103,G33116,G33129,G33142,G33155,G33168,G33181,G33194,G33207,G33220,G33233,G33246,G33259,G33272,G33285,G33298,G33311,G33324,G33337,G33350,G33363,G33376,G33389,G33402,G33415,G33428,G33441,G33454,G33467,G33480,G33493,G33506,G33519,G33532,G33545,G33558,G33571,G33584,G33597,G33610,G33623,G33636,G33649,G33662,G33675,G33688,G33701,G33714,G33727,G33740,G33753,G33766,G33779,G33792,G33805,G33818,G33831,G33844,G33857,G33870,G33883,G33896,G33909,G33922,G33935,G33948,G33961,G33974,G33987,G34000,G34013,G34026,G34039,G34052,G34065,G34078,G34091,G34104,G34117,G34130,G34143,G34156,G34169,G34182,G34195,G34208,G34221,G34234,G34247,G34260,G34273,G34286,G34299,G34312,G34325,G34338,G34351,G34364,G34377,G34390,G34403,G34416,G34429,G34442,G34455,G34468,G34481,G34494,G34507,G34520,G34533,G34546,G34559,G34572,G34585,G54748,G54761,G54774,G54787,G54800,G54813,G54826,G54839,G54852,G54865,G54878,G54891,G54904,G54917,G54930,G54943,G54956,G54969,G54982,G54995,G55008,G55021,G55034,G55047,G55060,G55073,G55086,G55099,G55112,G55125,G55138,G55151,G55164,G55177,G55190,G55203,G55216,G55229,G55242,G55255,G55268,G55281,G55294,G55307,G55320,G55333,G55346,G55359,G55372,G55385,G55398,G55411,G55424,G55437,G55450,G55463,G55476,G55489,G55502,G55515,G55528,G55541,G55554,G55567,G55580,G55593,G55606,G55619,G55632,G55645,G55658,G55671,G55684,G55697,G55710,G55723,G55736,G55749,G55762,G55775,G55788,G55801,G55814,G55827,G55840,G55853,G55866,G55879,G55892,G55905,G55918,G55931,G55944,G55957,G55970,G55983,G55996,G56009,G56022,G56035,G56048,G56061,G56074,G56087,G56100,G56113,G56126,G56139,G56152,G56165,G56178,G56191,G56204,G56217,G56230,G56243,G56256,G56269,G56282,G56295,G56308,G56321,G56334,G56347,G56360,G56373,G56386,G56399,G56412,G56425,G56438,G56451,G56464,G56477,G56490,G56503,G56516,G56529,G56542,G56555,G56568,G56581,G56594,G56607,G56620,G56633,G56646,G56659,G56672,G56685,G56698,G56711,G56724,G56737,G56750,G56763,G56776,G56789,G56802,G56815,G56828,G56841,G56854,G56867,G56880,G56893,G56906,G56919,G56932,G56945,G56958,G56971,G56984,G56997,G57010,G57023,G57036,G57049,G57062,G57075,G57088,G57101,G57114,G57127,G57140,G57153,G57166,G57179,G57192,G57205,G57218,G57231,G57244,G57257,G57270,G57283,G57296,G57309,G57322,G57335,G57348,G57361,G57374,G57387,G57400,G57413,G57426,G57439,G57452,G57465,G57478,G57491,G57504,G57517,G57530,G57543,G57556,G57569,G57582,G57595,G57608,G57621,G57634,G57647,G57660,G57673,G57686,G57699,G57712,G77875,G77888,G77901,G77914,G77927,G77940,G77953,G77966,G77979,G77992,G78005,G78018,G78031,G78044,G78057,G78070,G78083,G78096,G78109,G78122,G78135,G78148,G78161,G78174,G78187,G78200,G78213,G78226,G78239,G78252,G78265,G78278,G78291,G78304,G78317,G78330,G78343,G78356,G78369,G78382,G78395,G78408,G78421,G78434,G78447,G78460,G78473,G78486,G78499,G78512,G78525,G78538,G78551,G78564,G78577,G78590,G78603,G78616,G78629,G78642,G78655,G78668,G78681,G78694,G78707,G78720,G78733,G78746,G78759,G78772,G78785,G78798,G78811,G78824,G78837,G78850,G78863,G78876,G78889,G78902,G78915,G78928,G78941,G78954,G78967,G78980,G78993,G79006,G79019,G79032,G79045,G79058,G79071,G79084,G79097,G79110,G79123,G79136,G79149,G79162,G79175,G79188,G79201,G79214,G79227,G79240,G79253,G79266,G79279,G79292,G79305,G79318,G79331,G79344,G79357,G79370,G79383,G79396,G79409,G79422,G79435,G79448,G79461,G79474,G79487,G79500,G79513,G79526,G79539,G79552,G79565,G79578,G79591,G79604,G79617,G79630,G79643,G79656,G79669,G79682,G79695,G79708,G79721,G79734,G79747,G79760,G79773,G79786,G79799,G79812,G79825,G79838,G79851,G79864,G79877,G79890,G79903,G79916,G79929,G79942,G79955,G79968,G79981,G79994,G80007,G80020,G80033,G80046,G80059,G80072,G80085,G80098,G80111,G80124,G80137,G80150,G80163,G80176,G80189,G80202,G80215,G80228,G80241,G80254,G80267,G80280,G80293,G80306,G80319,G80332,G80345,G80358,G80371,G80384,G80397,G80410,G80423,G80436,G80449,G80462,G80475,G80488,G80501,G80514,G80527,G80540,G80553,G80566,G80579,G80592,G80605,G80618,G80631,G80644,G80657,G80670,G80683,G80696,G80709,G80722,G80735,G80748,G80761,G80774,G80787,G80800,G80813,G80826,G80839;
output G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G109,G110,G112,G114,G116,G118,G120,G122,G124,G126,G128,G130,G132,G134,G136,G138,G140,G142,G144,G146,G496,G509,G522,G535,G548,G561,G574,G587,G600,G613,G1306,G1327,G1348,G1369,G1390,G1411,G1432,G1453,G1514,G1535,G1556,G1577,G1598,G1619,G1640,G1661,G1722,G1743,G1764,G1785,G1806,G1827,G1848,G1869,G1930,G1951,G1972,G1993,G2014,G2035,G2056,G2077,G2138,G2159,G2180,G2201,G2222,G2243,G2264,G2285,G2346,G2367,G2388,G2409,G2430,G2451,G2472,G2493,G2554,G2575,G2596,G2617,G2638,G2659,G2680,G2701,G2762,G2783,G2804,G2825,G2846,G2867,G2888,G2909,G2970,G2991,G3012,G3033,G3054,G3075,G3096,G3117,G3178,G3199,G3220,G3241,G3262,G3283,G3304,G3325,G3386,G3407,G3428,G3449,G3470,G3491,G3512,G3533,G3554,G3615,G3636,G3657,G3678,G3699,G3720,G3741,G3762,G3823,G3844,G3865,G3886,G3907,G3928,G3949,G3970,G4031,G4052,G4073,G4094,G4115,G4136,G4157,G4178,G4239,G4260,G4281,G4302,G4323,G4344,G4365,G4386,G4407,G4468,G4489,G4510,G4531,G4552,G4573,G4594,G4615,G4676,G4697,G4718,G4739,G4760,G4781,G4802,G4823,G4884,G4905,G4926,G4947,G4968,G4989,G5010,G5031,G5092,G5113,G5134,G5155,G5176,G5197,G5239,G5260,G5321,G5342,G5363,G5384,G5405,G5426,G5447,G5468,G5529,G5550,G5571,G5592,G5613,G5634,G5655,G5676,G5737,G5758,G5779,G5800,G5821,G5842,G5863,G5884,G5945,G5966,G5987,G6008,G6029,G6050,G6071,G6092,G6153,G6174,G6195,G6216,G6237,G6258,G6279,G6300,G6361,G6382,G6403,G6424,G6445,G6466,G6487,G6508,G6569,G6590,G6611,G6632,G6653,G6674,G6695,G6716,G6777,G6798,G6819,G6840,G6861,G6882,G6903,G6924,G6985,G7006,G7027,G7048,G7069,G7090,G7111,G7132,G7193,G7214,G7235,G7256,G7277,G7298,G7319,G7340,G7401,G7422,G7443,G7464,G7485,G7506,G7527,G7548,G7609,G7630,G7651,G7672,G7693,G7714,G7735,G7756,G7817,G7838,G7859,G7880,G7901,G7922,G7943,G7964,G8025,G8046,G8067,G8088,G8109,G8130,G8151,G8172,G8233,G8254,G8275,G8296,G8317,G8338,G8359,G8380,G8441,G8462,G8483,G8504,G8525,G8546,G8567,G8588,G8649,G8691,G8712,G8733,G8754,G8775,G8796,G8857,G8878,G8899,G8920,G8941,G8962,G8983,G9004,G9065,G9086,G9107,G9128,G9149,G9170,G9191,G9212,G9273,G9294,G9315,G9336,G9357,G9378,G9399,G9420,G9481,G9502,G9523,G9544,G9565,G9586,G9607,G9628,G9689,G9710,G9731,G9752,G9773,G9794,G9815,G9836,G9897,G9918,G9939,G9960,G9981,G10002,G10023,G10044,G10105,G10126,G10147,G10168,G10189,G10210,G10231,G10252,G10313,G10334,G10355,G10376,G10397,G10418,G10439,G10460,G10521,G10542,G10563,G10584,G10605,G10626,G10647,G10668,G10729,G10750,G10771,G10792,G10813,G10834,G10855,G10876,G11344,G11365,G11386,G11407,G11428,G11449,G11470,G11492,G31630,G31643,G31656,G31669,G31682,G31695,G31708,G31721,G31734,G31747,G31760,G31773,G31786,G31799,G31812,G31825,G31838,G31851,G31864,G31877,G31890,G31903,G31916,G31929,G31942,G31955,G31968,G31981,G31994,G32007,G32020,G32033,G32046,G32059,G32072,G32085,G32098,G32111,G32124,G32137,G32150,G32163,G32176,G32189,G32202,G32215,G32228,G32241,G32254,G32267,G32280,G32293,G32306,G32319,G32332,G32345,G32358,G32371,G32384,G32397,G32410,G32423,G32436,G32449,G32462,G32475,G32488,G32501,G32514,G32527,G32540,G32553,G32566,G32579,G32592,G32605,G32618,G32631,G32644,G32657,G32670,G32683,G32696,G32709,G32722,G32735,G32748,G32761,G32774,G32787,G32800,G32813,G32826,G32839,G32852,G32865,G32878,G32891,G32904,G32917,G32930,G32943,G32956,G32969,G32982,G32995,G33008,G33021,G33034,G33047,G33060,G33073,G33086,G33099,G33112,G33125,G33138,G33151,G33164,G33177,G33190,G33203,G33216,G33229,G33242,G33255,G33268,G33281,G33294,G33307,G33320,G33333,G33346,G33359,G33372,G33385,G33398,G33411,G33424,G33437,G33450,G33463,G33476,G33489,G33502,G33515,G33528,G33541,G33554,G33567,G33580,G33593,G33606,G33619,G33632,G33645,G33658,G33671,G33684,G33697,G33710,G33723,G33736,G33749,G33762,G33775,G33788,G33801,G33814,G33827,G33840,G33853,G33866,G33879,G33892,G33905,G33918,G33931,G33944,G33957,G33970,G33983,G33996,G34009,G34022,G34035,G34048,G34061,G34074,G34087,G34100,G34113,G34126,G34139,G34152,G34165,G34178,G34191,G34204,G34217,G34230,G34243,G34256,G34269,G34282,G34295,G34308,G34321,G34334,G34347,G34373,G34386,G34399,G34412,G34425,G34438,G34451,G34464,G34477,G34490,G34503,G34516,G34529,G34542,G34555,G34568,G34581,G54757,G54770,G54783,G54796,G54809,G54822,G54835,G54848,G54861,G54874,G54887,G54900,G54913,G54926,G54939,G54952,G54965,G54978,G54991,G55004,G55017,G55030,G55043,G55056,G55069,G55082,G55095,G55108,G55121,G55134,G55147,G55160,G55173,G55186,G55199,G55212,G55225,G55238,G55251,G55264,G55277,G55290,G55303,G55316,G55329,G55342,G55355,G55368,G55381,G55394,G55407,G55420,G55433,G55446,G55459,G55472,G55485,G55498,G55511,G55524,G55537,G55550,G55563,G55576,G55589,G55602,G55615,G55628,G55641,G55654,G55667,G55680,G55693,G55706,G55719,G55732,G55745,G55758,G55771,G55784,G55797,G55810,G55823,G55836,G55849,G55862,G55875,G55888,G55901,G55914,G55927,G55940,G55953,G55966,G55979,G55992,G56005,G56018,G56031,G56044,G56057,G56070,G56083,G56096,G56109,G56122,G56135,G56148,G56161,G56174,G56187,G56200,G56213,G56226,G56239,G56252,G56265,G56278,G56291,G56304,G56317,G56330,G56343,G56356,G56369,G56382,G56395,G56408,G56421,G56434,G56447,G56460,G56473,G56486,G56499,G56512,G56525,G56538,G56551,G56564,G56577,G56590,G56603,G56616,G56629,G56642,G56655,G56668,G56681,G56694,G56707,G56720,G56733,G56746,G56759,G56772,G56785,G56798,G56811,G56824,G56837,G56850,G56863,G56876,G56889,G56902,G56915,G56928,G56941,G56954,G56967,G56980,G56993,G57006,G57019,G57032,G57045,G57058,G57071,G57084,G57097,G57110,G57123,G57136,G57149,G57162,G57175,G57188,G57201,G57214,G57227,G57240,G57253,G57266,G57279,G57292,G57305,G57318,G57331,G57357,G57370,G57383,G57396,G57409,G57422,G57435,G57448,G57461,G57474,G57487,G57500,G57513,G57526,G57539,G57552,G57578,G57591,G57604,G57617,G57630,G57643,G57656,G57669,G57682,G57695,G57708,G57721,G77884,G77897,G77910,G77923,G77936,G77949,G77962,G77975,G77988,G78001,G78014,G78027,G78040,G78053,G78066,G78079,G78092,G78105,G78118,G78131,G78144,G78157,G78170,G78183,G78196,G78209,G78222,G78235,G78248,G78261,G78274,G78287,G78300,G78313,G78326,G78339,G78352,G78365,G78378,G78391,G78404,G78417,G78430,G78443,G78456,G78469,G78482,G78495,G78508,G78521,G78534,G78547,G78560,G78573,G78586,G78599,G78612,G78625,G78638,G78651,G78664,G78677,G78690,G78703,G78716,G78729,G78742,G78755,G78768,G78781,G78794,G78807,G78820,G78833,G78846,G78859,G78872,G78885,G78898,G78911,G78924,G78937,G78950,G78963,G78976,G78989,G79002,G79015,G79028,G79041,G79054,G79067,G79080,G79093,G79106,G79119,G79132,G79145,G79158,G79171,G79184,G79197,G79210,G79223,G79236,G79249,G79262,G79275,G79288,G79301,G79314,G79327,G79340,G79353,G79366,G79379,G79392,G79405,G79418,G79431,G79444,G79457,G79470,G79483,G79496,G79509,G79522,G79535,G79548,G79561,G79574,G79587,G79600,G79613,G79626,G79639,G79652,G79665,G79678,G79691,G79704,G79717,G79730,G79743,G79756,G79769,G79782,G79795,G79808,G79821,G79834,G79847,G79860,G79873,G79886,G79899,G79912,G79925,G79938,G79951,G79964,G79977,G79990,G80003,G80016,G80029,G80042,G80055,G80068,G80081,G80094,G80107,G80120,G80133,G80146,G80159,G80172,G80185,G80211,G80224,G80237,G80250,G80263,G80276,G80289,G80302,G80315,G80328,G80341,G80354,G80367,G80380,G80393,G80406,G80419,G80432,G80445,G80458,G80471,G80484,G80497,G80510,G80523,G80536,G80549,G80562,G80575,G80588,G80601,G80614,G80627,G80640,G80653,G80679,G80692,G80705,G80731,G80744,G80757,G80770,G80783,G80796,G80809,G80822,G80835,G80848;

  wire G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
       G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,
       G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60,
       G61,G62,G63,G64,G65,G66,G67,G68,G80,
       G81,G82,G83,G84,G85,G86,G87,G88,G89,G90,G91,G92,G93,G94,G95,G96,G97,G98,G99,G100,
       G101,G102,G103,G104,G105,G106,G107,G108,G109,G110,G111,G112,G113,G114,G115,G116,G117,G118,G119,G120,
       G121,G122,G123,G124,G125,G126,G127,G128,G129,G130,G131,G132,G133,G134,G135,G136,G137,G138,G139,G140,
       G141,G142,G143,G144,G145,G146,G147,G148,G149,G150,G151,G152,G153,G154,G155,G156,G157,G158,G159,G160,
       G161,G162,G163,G164,G165,G166,G167,G168,G169,G170,G171,G172,G173,G174,G175,G176,G177,G178,G179,G180,
       G181,G182,G183,G184,G185,G186,G187,G188,G189,G190,G191,G192,G193,G194,G195,G196,G197,G198,G199,G200,
       G201,G202,G203,G204,G205,G206,G207,G208,G209,G210,G211,G212,G213,G214,G215,G216,G217,G218,G219,G220,
       G221,G222,G223,G224,G225,G226,G227,G228,G229,G230,G231,G232,G233,G234,G235,G236,G237,G238,G239,G240,
       G241,G242,G243,G244,G245,G246,G247,G248,G249,G250,G251,G252,G253,G254,G255,G256,G257,G258,G259,G260,
       G261,G262,G263,G264,G265,G266,G267,G268,G269,G270,G271,G272,G273,G274,G275,G276,G277,G278,G279,G280,
       G281,G282,G283,G284,G285,G286,G287,G288,G289,G290,G291,G292,G293,G294,G295,G296,G297,G298,G299,G300,
       G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G311,G312,G313,G314,G315,G316,G317,G318,G319,G320,
       G321,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,
       G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G358,G359,G360,
       G361,G362,G363,G364,G365,G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
       G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,G396,G397,G398,G399,G400,
       G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,
       G421,G422,G423,G424,G425,G426,G427,G428,G429,G430,G431,G432,G433,G434,G435,G436,G437,G438,G439,G440,
       G441,G442,G443,G444,G445,G446,G447,G448,G449,G450,G451,G452,G453,G454,G455,G456,G457,G458,G459,G460,
       G461,G462,G463,G464,G465,G466,G467,G468,G469,G470,G471,G472,G473,G474,G475,G476,G477,G478,G479,G480,
       G481,G482,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,
       G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G516,G517,G518,G519,G520,
       G521,G522,G523,G524,G525,G526,G527,G528,G529,G530,G531,G532,G533,G534,G535,G536,G537,G538,G539,G540,
       G541,G542,G543,G544,G545,G546,G547,G548,G549,G550,G551,G552,G553,G554,G555,G556,G557,G558,G559,G560,
       G561,G562,G563,G564,G565,G566,G567,G568,G569,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,
       G581,G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,G597,G598,G599,G600,
       G601,G602,G603,G604,G605,G606,G607,G608,G609,G610,G611,G612,G613,G614,G615,G616,G617,G618,G619,G620,
       G621,G622,G623,G624,G625,G626,G627,G628,G629,G630,G631,G632,G633,G634,G635,G636,G637,G638,G639,G640,
       G641,G642,G643,G644,G645,G646,G647,G648,G649,G650,G651,G652,G653,G654,G655,G656,G657,G658,G659,G660,
       G661,G662,G663,G664,G665,G666,G667,G668,G669,G670,G671,G672,G673,G674,G675,G676,G677,G678,G679,G680,
       G681,G682,G683,G684,G685,G686,G687,G688,G689,G690,G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,
       G701,G702,G703,G704,G705,G706,G707,G708,G709,G710,G711,G712,G713,G714,G715,G716,G717,G718,G719,G720,
       G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,
       G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G757,G758,G759,G760,
       G761,G762,G763,G764,G765,G766,G767,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G780,
       G781,G782,G783,G784,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G799,G800,
       G801,G802,G803,G804,G805,G806,G807,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,
       G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,
       G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854,G855,G856,G857,G858,G859,G860,
       G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,
       G881,G882,G883,G884,G885,G886,G887,G888,G889,G890,G891,G892,G893,G894,G895,G896,G897,G898,G899,G900,
       G901,G902,G903,G904,G905,G906,G907,G908,G909,G910,G911,G912,G913,G914,G915,G916,G917,G918,G919,G920,
       G921,G922,G923,G924,G925,G926,G927,G928,G929,G930,G931,G932,G933,G934,G935,G936,G937,G938,G939,G940,
       G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,G956,G957,G958,G959,G960,
       G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,
       G981,G982,G983,G984,G985,G986,G987,G988,G989,G990,G991,G992,G993,G994,G995,G996,G997,G998,G999,G1000,
       G1001,G1002,G1003,G1004,G1005,G1006,G1007,G1008,G1009,G1010,G1011,G1012,G1013,G1014,G1015,G1016,G1017,G1018,G1019,G1020,
       G1021,G1022,G1023,G1024,G1025,G1026,G1027,G1028,G1029,G1030,G1031,G1032,G1033,G1034,G1035,G1036,G1037,G1038,G1039,G1040,
       G1041,G1042,G1043,G1044,G1045,G1046,G1047,G1048,G1049,G1050,G1051,G1052,G1053,G1054,G1055,G1056,G1057,G1058,G1059,G1060,
       G1061,G1062,G1063,G1064,G1065,G1066,G1067,G1068,G1069,G1070,G1071,G1072,G1073,G1074,G1075,G1076,G1077,G1078,G1079,G1080,
       G1081,G1082,G1083,G1084,G1085,G1086,G1087,G1088,G1089,G1090,G1091,G1092,G1093,G1094,G1095,G1096,G1097,G1098,G1099,G1100,
       G1101,G1102,G1103,G1104,G1105,G1106,G1107,G1108,G1109,G1110,G1111,G1112,G1113,G1114,G1115,G1116,G1117,G1118,G1119,G1120,
       G1121,G1122,G1123,G1124,G1125,G1126,G1127,G1128,G1129,G1130,G1131,G1132,G1133,G1134,G1135,G1136,G1137,G1138,G1139,G1140,
       G1141,G1142,G1143,G1144,G1145,G1146,G1147,G1148,G1149,G1150,G1151,G1152,G1153,G1154,G1155,G1156,G1157,G1158,G1159,G1160,
       G1161,G1162,G1163,G1164,G1165,G1166,G1167,G1168,G1169,G1170,G1171,G1172,G1173,G1174,G1175,G1176,G1177,G1178,G1179,G1180,
       G1181,G1182,G1183,G1184,G1185,G1186,G1187,G1188,G1189,G1190,G1191,G1192,G1193,G1194,G1195,G1196,G1197,G1198,G1199,G1200,
       G1201,G1202,G1203,G1204,G1205,G1206,G1207,G1208,G1209,G1210,G1211,G1212,G1213,G1214,G1215,G1216,G1217,G1218,G1219,G1220,
       G1221,G1222,G1223,G1224,G1225,G1226,G1227,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,G1239,G1240,
       G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,
       G1261,G1262,G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,G1275,G1276,G1277,G1278,G1279,G1280,
       G1281,G1282,G1283,G1284,G1285,G1286,G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,G1299,G1300,
       G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,
       G1321,G1322,G1323,G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,
       G1341,G1342,G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355,G1356,G1357,G1358,G1359,G1360,
       G1361,G1362,G1363,G1364,G1365,G1366,G1367,G1368,G1369,G1370,G1371,G1372,G1373,G1374,G1375,G1376,G1377,G1378,G1379,G1380,
       G1381,G1382,G1383,G1384,G1385,G1386,G1387,G1388,G1389,G1390,G1391,G1392,G1393,G1394,G1395,G1396,G1397,G1398,G1399,G1400,
       G1401,G1402,G1403,G1404,G1405,G1406,G1407,G1408,G1409,G1410,G1411,G1412,G1413,G1414,G1415,G1416,G1417,G1418,G1419,G1420,
       G1421,G1422,G1423,G1424,G1425,G1426,G1427,G1428,G1429,G1430,G1431,G1432,G1433,G1434,G1435,G1436,G1437,G1438,G1439,G1440,
       G1441,G1442,G1443,G1444,G1445,G1446,G1447,G1448,G1449,G1450,G1451,G1452,G1453,G1454,G1455,G1456,G1457,G1458,G1459,G1460,
       G1461,G1462,G1463,G1464,G1465,G1466,G1467,G1468,G1469,G1470,G1471,G1472,G1473,G1474,G1475,G1476,G1477,G1478,G1479,G1480,
       G1481,G1482,G1483,G1484,G1485,G1486,G1487,G1488,G1489,G1490,G1491,G1492,G1493,G1494,G1495,G1496,G1497,G1498,G1499,G1500,
       G1501,G1502,G1503,G1504,G1505,G1506,G1507,G1508,G1509,G1510,G1511,G1512,G1513,G1514,G1515,G1516,G1517,G1518,G1519,G1520,
       G1521,G1522,G1523,G1524,G1525,G1526,G1527,G1528,G1529,G1530,G1531,G1532,G1533,G1534,G1535,G1536,G1537,G1538,G1539,G1540,
       G1541,G1542,G1543,G1544,G1545,G1546,G1547,G1548,G1549,G1550,G1551,G1552,G1553,G1554,G1555,G1556,G1557,G1558,G1559,G1560,
       G1561,G1562,G1563,G1564,G1565,G1566,G1567,G1568,G1569,G1570,G1571,G1572,G1573,G1574,G1575,G1576,G1577,G1578,G1579,G1580,
       G1581,G1582,G1583,G1584,G1585,G1586,G1587,G1588,G1589,G1590,G1591,G1592,G1593,G1594,G1595,G1596,G1597,G1598,G1599,G1600,
       G1601,G1602,G1603,G1604,G1605,G1606,G1607,G1608,G1609,G1610,G1611,G1612,G1613,G1614,G1615,G1616,G1617,G1618,G1619,G1620,
       G1621,G1622,G1623,G1624,G1625,G1626,G1627,G1628,G1629,G1630,G1631,G1632,G1633,G1634,G1635,G1636,G1637,G1638,G1639,G1640,
       G1641,G1642,G1643,G1644,G1645,G1646,G1647,G1648,G1649,G1650,G1651,G1652,G1653,G1654,G1655,G1656,G1657,G1658,G1659,G1660,
       G1661,G1662,G1663,G1664,G1665,G1666,G1667,G1668,G1669,G1670,G1671,G1672,G1673,G1674,G1675,G1676,G1677,G1678,G1679,G1680,
       G1681,G1682,G1683,G1684,G1685,G1686,G1687,G1688,G1689,G1690,G1691,G1692,G1693,G1694,G1695,G1696,G1697,G1698,G1699,G1700,
       G1701,G1702,G1703,G1704,G1705,G1706,G1707,G1708,G1709,G1710,G1711,G1712,G1713,G1714,G1715,G1716,G1717,G1718,G1719,G1720,
       G1721,G1722,G1723,G1724,G1725,G1726,G1727,G1728,G1729,G1730,G1731,G1732,G1733,G1734,G1735,G1736,G1737,G1738,G1739,G1740,
       G1741,G1742,G1743,G1744,G1745,G1746,G1747,G1748,G1749,G1750,G1751,G1752,G1753,G1754,G1755,G1756,G1757,G1758,G1759,G1760,
       G1761,G1762,G1763,G1764,G1765,G1766,G1767,G1768,G1769,G1770,G1771,G1772,G1773,G1774,G1775,G1776,G1777,G1778,G1779,G1780,
       G1781,G1782,G1783,G1784,G1785,G1786,G1787,G1788,G1789,G1790,G1791,G1792,G1793,G1794,G1795,G1796,G1797,G1798,G1799,G1800,
       G1801,G1802,G1803,G1804,G1805,G1806,G1807,G1808,G1809,G1810,G1811,G1812,G1813,G1814,G1815,G1816,G1817,G1818,G1819,G1820,
       G1821,G1822,G1823,G1824,G1825,G1826,G1827,G1828,G1829,G1830,G1831,G1832,G1833,G1834,G1835,G1836,G1837,G1838,G1839,G1840,
       G1841,G1842,G1843,G1844,G1845,G1846,G1847,G1848,G1849,G1850,G1851,G1852,G1853,G1854,G1855,G1856,G1857,G1858,G1859,G1860,
       G1861,G1862,G1863,G1864,G1865,G1866,G1867,G1868,G1869,G1870,G1871,G1872,G1873,G1874,G1875,G1876,G1877,G1878,G1879,G1880,
       G1881,G1882,G1883,G1884,G1885,G1886,G1887,G1888,G1889,G1890,G1891,G1892,G1893,G1894,G1895,G1896,G1897,G1898,G1899,G1900,
       G1901,G1902,G1903,G1904,G1905,G1906,G1907,G1908,G1909,G1910,G1911,G1912,G1913,G1914,G1915,G1916,G1917,G1918,G1919,G1920,
       G1921,G1922,G1923,G1924,G1925,G1926,G1927,G1928,G1929,G1930,G1931,G1932,G1933,G1934,G1935,G1936,G1937,G1938,G1939,G1940,
       G1941,G1942,G1943,G1944,G1945,G1946,G1947,G1948,G1949,G1950,G1951,G1952,G1953,G1954,G1955,G1956,G1957,G1958,G1959,G1960,
       G1961,G1962,G1963,G1964,G1965,G1966,G1967,G1968,G1969,G1970,G1971,G1972,G1973,G1974,G1975,G1976,G1977,G1978,G1979,G1980,
       G1981,G1982,G1983,G1984,G1985,G1986,G1987,G1988,G1989,G1990,G1991,G1992,G1993,G1994,G1995,G1996,G1997,G1998,G1999,G2000,
       G2001,G2002,G2003,G2004,G2005,G2006,G2007,G2008,G2009,G2010,G2011,G2012,G2013,G2014,G2015,G2016,G2017,G2018,G2019,G2020,
       G2021,G2022,G2023,G2024,G2025,G2026,G2027,G2028,G2029,G2030,G2031,G2032,G2033,G2034,G2035,G2036,G2037,G2038,G2039,G2040,
       G2041,G2042,G2043,G2044,G2045,G2046,G2047,G2048,G2049,G2050,G2051,G2052,G2053,G2054,G2055,G2056,G2057,G2058,G2059,G2060,
       G2061,G2062,G2063,G2064,G2065,G2066,G2067,G2068,G2069,G2070,G2071,G2072,G2073,G2074,G2075,G2076,G2077,G2078,G2079,G2080,
       G2081,G2082,G2083,G2084,G2085,G2086,G2087,G2088,G2089,G2090,G2091,G2092,G2093,G2094,G2095,G2096,G2097,G2098,G2099,G2100,
       G2101,G2102,G2103,G2104,G2105,G2106,G2107,G2108,G2109,G2110,G2111,G2112,G2113,G2114,G2115,G2116,G2117,G2118,G2119,G2120,
       G2121,G2122,G2123,G2124,G2125,G2126,G2127,G2128,G2129,G2130,G2131,G2132,G2133,G2134,G2135,G2136,G2137,G2138,G2139,G2140,
       G2141,G2142,G2143,G2144,G2145,G2146,G2147,G2148,G2149,G2150,G2151,G2152,G2153,G2154,G2155,G2156,G2157,G2158,G2159,G2160,
       G2161,G2162,G2163,G2164,G2165,G2166,G2167,G2168,G2169,G2170,G2171,G2172,G2173,G2174,G2175,G2176,G2177,G2178,G2179,G2180,
       G2181,G2182,G2183,G2184,G2185,G2186,G2187,G2188,G2189,G2190,G2191,G2192,G2193,G2194,G2195,G2196,G2197,G2198,G2199,G2200,
       G2201,G2202,G2203,G2204,G2205,G2206,G2207,G2208,G2209,G2210,G2211,G2212,G2213,G2214,G2215,G2216,G2217,G2218,G2219,G2220,
       G2221,G2222,G2223,G2224,G2225,G2226,G2227,G2228,G2229,G2230,G2231,G2232,G2233,G2234,G2235,G2236,G2237,G2238,G2239,G2240,
       G2241,G2242,G2243,G2244,G2245,G2246,G2247,G2248,G2249,G2250,G2251,G2252,G2253,G2254,G2255,G2256,G2257,G2258,G2259,G2260,
       G2261,G2262,G2263,G2264,G2265,G2266,G2267,G2268,G2269,G2270,G2271,G2272,G2273,G2274,G2275,G2276,G2277,G2278,G2279,G2280,
       G2281,G2282,G2283,G2284,G2285,G2286,G2287,G2288,G2289,G2290,G2291,G2292,G2293,G2294,G2295,G2296,G2297,G2298,G2299,G2300,
       G2301,G2302,G2303,G2304,G2305,G2306,G2307,G2308,G2309,G2310,G2311,G2312,G2313,G2314,G2315,G2316,G2317,G2318,G2319,G2320,
       G2321,G2322,G2323,G2324,G2325,G2326,G2327,G2328,G2329,G2330,G2331,G2332,G2333,G2334,G2335,G2336,G2337,G2338,G2339,G2340,
       G2341,G2342,G2343,G2344,G2345,G2346,G2347,G2348,G2349,G2350,G2351,G2352,G2353,G2354,G2355,G2356,G2357,G2358,G2359,G2360,
       G2361,G2362,G2363,G2364,G2365,G2366,G2367,G2368,G2369,G2370,G2371,G2372,G2373,G2374,G2375,G2376,G2377,G2378,G2379,G2380,
       G2381,G2382,G2383,G2384,G2385,G2386,G2387,G2388,G2389,G2390,G2391,G2392,G2393,G2394,G2395,G2396,G2397,G2398,G2399,G2400,
       G2401,G2402,G2403,G2404,G2405,G2406,G2407,G2408,G2409,G2410,G2411,G2412,G2413,G2414,G2415,G2416,G2417,G2418,G2419,G2420,
       G2421,G2422,G2423,G2424,G2425,G2426,G2427,G2428,G2429,G2430,G2431,G2432,G2433,G2434,G2435,G2436,G2437,G2438,G2439,G2440,
       G2441,G2442,G2443,G2444,G2445,G2446,G2447,G2448,G2449,G2450,G2451,G2452,G2453,G2454,G2455,G2456,G2457,G2458,G2459,G2460,
       G2461,G2462,G2463,G2464,G2465,G2466,G2467,G2468,G2469,G2470,G2471,G2472,G2473,G2474,G2475,G2476,G2477,G2478,G2479,G2480,
       G2481,G2482,G2483,G2484,G2485,G2486,G2487,G2488,G2489,G2490,G2491,G2492,G2493,G2494,G2495,G2496,G2497,G2498,G2499,G2500,
       G2501,G2502,G2503,G2504,G2505,G2506,G2507,G2508,G2509,G2510,G2511,G2512,G2513,G2514,G2515,G2516,G2517,G2518,G2519,G2520,
       G2521,G2522,G2523,G2524,G2525,G2526,G2527,G2528,G2529,G2530,G2531,G2532,G2533,G2534,G2535,G2536,G2537,G2538,G2539,G2540,
       G2541,G2542,G2543,G2544,G2545,G2546,G2547,G2548,G2549,G2550,G2551,G2552,G2553,G2554,G2555,G2556,G2557,G2558,G2559,G2560,
       G2561,G2562,G2563,G2564,G2565,G2566,G2567,G2568,G2569,G2570,G2571,G2572,G2573,G2574,G2575,G2576,G2577,G2578,G2579,G2580,
       G2581,G2582,G2583,G2584,G2585,G2586,G2587,G2588,G2589,G2590,G2591,G2592,G2593,G2594,G2595,G2596,G2597,G2598,G2599,G2600,
       G2601,G2602,G2603,G2604,G2605,G2606,G2607,G2608,G2609,G2610,G2611,G2612,G2613,G2614,G2615,G2616,G2617,G2618,G2619,G2620,
       G2621,G2622,G2623,G2624,G2625,G2626,G2627,G2628,G2629,G2630,G2631,G2632,G2633,G2634,G2635,G2636,G2637,G2638,G2639,G2640,
       G2641,G2642,G2643,G2644,G2645,G2646,G2647,G2648,G2649,G2650,G2651,G2652,G2653,G2654,G2655,G2656,G2657,G2658,G2659,G2660,
       G2661,G2662,G2663,G2664,G2665,G2666,G2667,G2668,G2669,G2670,G2671,G2672,G2673,G2674,G2675,G2676,G2677,G2678,G2679,G2680,
       G2681,G2682,G2683,G2684,G2685,G2686,G2687,G2688,G2689,G2690,G2691,G2692,G2693,G2694,G2695,G2696,G2697,G2698,G2699,G2700,
       G2701,G2702,G2703,G2704,G2705,G2706,G2707,G2708,G2709,G2710,G2711,G2712,G2713,G2714,G2715,G2716,G2717,G2718,G2719,G2720,
       G2721,G2722,G2723,G2724,G2725,G2726,G2727,G2728,G2729,G2730,G2731,G2732,G2733,G2734,G2735,G2736,G2737,G2738,G2739,G2740,
       G2741,G2742,G2743,G2744,G2745,G2746,G2747,G2748,G2749,G2750,G2751,G2752,G2753,G2754,G2755,G2756,G2757,G2758,G2759,G2760,
       G2761,G2762,G2763,G2764,G2765,G2766,G2767,G2768,G2769,G2770,G2771,G2772,G2773,G2774,G2775,G2776,G2777,G2778,G2779,G2780,
       G2781,G2782,G2783,G2784,G2785,G2786,G2787,G2788,G2789,G2790,G2791,G2792,G2793,G2794,G2795,G2796,G2797,G2798,G2799,G2800,
       G2801,G2802,G2803,G2804,G2805,G2806,G2807,G2808,G2809,G2810,G2811,G2812,G2813,G2814,G2815,G2816,G2817,G2818,G2819,G2820,
       G2821,G2822,G2823,G2824,G2825,G2826,G2827,G2828,G2829,G2830,G2831,G2832,G2833,G2834,G2835,G2836,G2837,G2838,G2839,G2840,
       G2841,G2842,G2843,G2844,G2845,G2846,G2847,G2848,G2849,G2850,G2851,G2852,G2853,G2854,G2855,G2856,G2857,G2858,G2859,G2860,
       G2861,G2862,G2863,G2864,G2865,G2866,G2867,G2868,G2869,G2870,G2871,G2872,G2873,G2874,G2875,G2876,G2877,G2878,G2879,G2880,
       G2881,G2882,G2883,G2884,G2885,G2886,G2887,G2888,G2889,G2890,G2891,G2892,G2893,G2894,G2895,G2896,G2897,G2898,G2899,G2900,
       G2901,G2902,G2903,G2904,G2905,G2906,G2907,G2908,G2909,G2910,G2911,G2912,G2913,G2914,G2915,G2916,G2917,G2918,G2919,G2920,
       G2921,G2922,G2923,G2924,G2925,G2926,G2927,G2928,G2929,G2930,G2931,G2932,G2933,G2934,G2935,G2936,G2937,G2938,G2939,G2940,
       G2941,G2942,G2943,G2944,G2945,G2946,G2947,G2948,G2949,G2950,G2951,G2952,G2953,G2954,G2955,G2956,G2957,G2958,G2959,G2960,
       G2961,G2962,G2963,G2964,G2965,G2966,G2967,G2968,G2969,G2970,G2971,G2972,G2973,G2974,G2975,G2976,G2977,G2978,G2979,G2980,
       G2981,G2982,G2983,G2984,G2985,G2986,G2987,G2988,G2989,G2990,G2991,G2992,G2993,G2994,G2995,G2996,G2997,G2998,G2999,G3000,
       G3001,G3002,G3003,G3004,G3005,G3006,G3007,G3008,G3009,G3010,G3011,G3012,G3013,G3014,G3015,G3016,G3017,G3018,G3019,G3020,
       G3021,G3022,G3023,G3024,G3025,G3026,G3027,G3028,G3029,G3030,G3031,G3032,G3033,G3034,G3035,G3036,G3037,G3038,G3039,G3040,
       G3041,G3042,G3043,G3044,G3045,G3046,G3047,G3048,G3049,G3050,G3051,G3052,G3053,G3054,G3055,G3056,G3057,G3058,G3059,G3060,
       G3061,G3062,G3063,G3064,G3065,G3066,G3067,G3068,G3069,G3070,G3071,G3072,G3073,G3074,G3075,G3076,G3077,G3078,G3079,G3080,
       G3081,G3082,G3083,G3084,G3085,G3086,G3087,G3088,G3089,G3090,G3091,G3092,G3093,G3094,G3095,G3096,G3097,G3098,G3099,G3100,
       G3101,G3102,G3103,G3104,G3105,G3106,G3107,G3108,G3109,G3110,G3111,G3112,G3113,G3114,G3115,G3116,G3117,G3118,G3119,G3120,
       G3121,G3122,G3123,G3124,G3125,G3126,G3127,G3128,G3129,G3130,G3131,G3132,G3133,G3134,G3135,G3136,G3137,G3138,G3139,G3140,
       G3141,G3142,G3143,G3144,G3145,G3146,G3147,G3148,G3149,G3150,G3151,G3152,G3153,G3154,G3155,G3156,G3157,G3158,G3159,G3160,
       G3161,G3162,G3163,G3164,G3165,G3166,G3167,G3168,G3169,G3170,G3171,G3172,G3173,G3174,G3175,G3176,G3177,G3178,G3179,G3180,
       G3181,G3182,G3183,G3184,G3185,G3186,G3187,G3188,G3189,G3190,G3191,G3192,G3193,G3194,G3195,G3196,G3197,G3198,G3199,G3200,
       G3201,G3202,G3203,G3204,G3205,G3206,G3207,G3208,G3209,G3210,G3211,G3212,G3213,G3214,G3215,G3216,G3217,G3218,G3219,G3220,
       G3221,G3222,G3223,G3224,G3225,G3226,G3227,G3228,G3229,G3230,G3231,G3232,G3233,G3234,G3235,G3236,G3237,G3238,G3239,G3240,
       G3241,G3242,G3243,G3244,G3245,G3246,G3247,G3248,G3249,G3250,G3251,G3252,G3253,G3254,G3255,G3256,G3257,G3258,G3259,G3260,
       G3261,G3262,G3263,G3264,G3265,G3266,G3267,G3268,G3269,G3270,G3271,G3272,G3273,G3274,G3275,G3276,G3277,G3278,G3279,G3280,
       G3281,G3282,G3283,G3284,G3285,G3286,G3287,G3288,G3289,G3290,G3291,G3292,G3293,G3294,G3295,G3296,G3297,G3298,G3299,G3300,
       G3301,G3302,G3303,G3304,G3305,G3306,G3307,G3308,G3309,G3310,G3311,G3312,G3313,G3314,G3315,G3316,G3317,G3318,G3319,G3320,
       G3321,G3322,G3323,G3324,G3325,G3326,G3327,G3328,G3329,G3330,G3331,G3332,G3333,G3334,G3335,G3336,G3337,G3338,G3339,G3340,
       G3341,G3342,G3343,G3344,G3345,G3346,G3347,G3348,G3349,G3350,G3351,G3352,G3353,G3354,G3355,G3356,G3357,G3358,G3359,G3360,
       G3361,G3362,G3363,G3364,G3365,G3366,G3367,G3368,G3369,G3370,G3371,G3372,G3373,G3374,G3375,G3376,G3377,G3378,G3379,G3380,
       G3381,G3382,G3383,G3384,G3385,G3386,G3387,G3388,G3389,G3390,G3391,G3392,G3393,G3394,G3395,G3396,G3397,G3398,G3399,G3400,
       G3401,G3402,G3403,G3404,G3405,G3406,G3407,G3408,G3409,G3410,G3411,G3412,G3413,G3414,G3415,G3416,G3417,G3418,G3419,G3420,
       G3421,G3422,G3423,G3424,G3425,G3426,G3427,G3428,G3429,G3430,G3431,G3432,G3433,G3434,G3435,G3436,G3437,G3438,G3439,G3440,
       G3441,G3442,G3443,G3444,G3445,G3446,G3447,G3448,G3449,G3450,G3451,G3452,G3453,G3454,G3455,G3456,G3457,G3458,G3459,G3460,
       G3461,G3462,G3463,G3464,G3465,G3466,G3467,G3468,G3469,G3470,G3471,G3472,G3473,G3474,G3475,G3476,G3477,G3478,G3479,G3480,
       G3481,G3482,G3483,G3484,G3485,G3486,G3487,G3488,G3489,G3490,G3491,G3492,G3493,G3494,G3495,G3496,G3497,G3498,G3499,G3500,
       G3501,G3502,G3503,G3504,G3505,G3506,G3507,G3508,G3509,G3510,G3511,G3512,G3513,G3514,G3515,G3516,G3517,G3518,G3519,G3520,
       G3521,G3522,G3523,G3524,G3525,G3526,G3527,G3528,G3529,G3530,G3531,G3532,G3533,G3534,G3535,G3536,G3537,G3538,G3539,G3540,
       G3541,G3542,G3543,G3544,G3545,G3546,G3547,G3548,G3549,G3550,G3551,G3552,G3553,G3554,G3555,G3556,G3557,G3558,G3559,G3560,
       G3561,G3562,G3563,G3564,G3565,G3566,G3567,G3568,G3569,G3570,G3571,G3572,G3573,G3574,G3575,G3576,G3577,G3578,G3579,G3580,
       G3581,G3582,G3583,G3584,G3585,G3586,G3587,G3588,G3589,G3590,G3591,G3592,G3593,G3594,G3595,G3596,G3597,G3598,G3599,G3600,
       G3601,G3602,G3603,G3604,G3605,G3606,G3607,G3608,G3609,G3610,G3611,G3612,G3613,G3614,G3615,G3616,G3617,G3618,G3619,G3620,
       G3621,G3622,G3623,G3624,G3625,G3626,G3627,G3628,G3629,G3630,G3631,G3632,G3633,G3634,G3635,G3636,G3637,G3638,G3639,G3640,
       G3641,G3642,G3643,G3644,G3645,G3646,G3647,G3648,G3649,G3650,G3651,G3652,G3653,G3654,G3655,G3656,G3657,G3658,G3659,G3660,
       G3661,G3662,G3663,G3664,G3665,G3666,G3667,G3668,G3669,G3670,G3671,G3672,G3673,G3674,G3675,G3676,G3677,G3678,G3679,G3680,
       G3681,G3682,G3683,G3684,G3685,G3686,G3687,G3688,G3689,G3690,G3691,G3692,G3693,G3694,G3695,G3696,G3697,G3698,G3699,G3700,
       G3701,G3702,G3703,G3704,G3705,G3706,G3707,G3708,G3709,G3710,G3711,G3712,G3713,G3714,G3715,G3716,G3717,G3718,G3719,G3720,
       G3721,G3722,G3723,G3724,G3725,G3726,G3727,G3728,G3729,G3730,G3731,G3732,G3733,G3734,G3735,G3736,G3737,G3738,G3739,G3740,
       G3741,G3742,G3743,G3744,G3745,G3746,G3747,G3748,G3749,G3750,G3751,G3752,G3753,G3754,G3755,G3756,G3757,G3758,G3759,G3760,
       G3761,G3762,G3763,G3764,G3765,G3766,G3767,G3768,G3769,G3770,G3771,G3772,G3773,G3774,G3775,G3776,G3777,G3778,G3779,G3780,
       G3781,G3782,G3783,G3784,G3785,G3786,G3787,G3788,G3789,G3790,G3791,G3792,G3793,G3794,G3795,G3796,G3797,G3798,G3799,G3800,
       G3801,G3802,G3803,G3804,G3805,G3806,G3807,G3808,G3809,G3810,G3811,G3812,G3813,G3814,G3815,G3816,G3817,G3818,G3819,G3820,
       G3821,G3822,G3823,G3824,G3825,G3826,G3827,G3828,G3829,G3830,G3831,G3832,G3833,G3834,G3835,G3836,G3837,G3838,G3839,G3840,
       G3841,G3842,G3843,G3844,G3845,G3846,G3847,G3848,G3849,G3850,G3851,G3852,G3853,G3854,G3855,G3856,G3857,G3858,G3859,G3860,
       G3861,G3862,G3863,G3864,G3865,G3866,G3867,G3868,G3869,G3870,G3871,G3872,G3873,G3874,G3875,G3876,G3877,G3878,G3879,G3880,
       G3881,G3882,G3883,G3884,G3885,G3886,G3887,G3888,G3889,G3890,G3891,G3892,G3893,G3894,G3895,G3896,G3897,G3898,G3899,G3900,
       G3901,G3902,G3903,G3904,G3905,G3906,G3907,G3908,G3909,G3910,G3911,G3912,G3913,G3914,G3915,G3916,G3917,G3918,G3919,G3920,
       G3921,G3922,G3923,G3924,G3925,G3926,G3927,G3928,G3929,G3930,G3931,G3932,G3933,G3934,G3935,G3936,G3937,G3938,G3939,G3940,
       G3941,G3942,G3943,G3944,G3945,G3946,G3947,G3948,G3949,G3950,G3951,G3952,G3953,G3954,G3955,G3956,G3957,G3958,G3959,G3960,
       G3961,G3962,G3963,G3964,G3965,G3966,G3967,G3968,G3969,G3970,G3971,G3972,G3973,G3974,G3975,G3976,G3977,G3978,G3979,G3980,
       G3981,G3982,G3983,G3984,G3985,G3986,G3987,G3988,G3989,G3990,G3991,G3992,G3993,G3994,G3995,G3996,G3997,G3998,G3999,G4000,
       G4001,G4002,G4003,G4004,G4005,G4006,G4007,G4008,G4009,G4010,G4011,G4012,G4013,G4014,G4015,G4016,G4017,G4018,G4019,G4020,
       G4021,G4022,G4023,G4024,G4025,G4026,G4027,G4028,G4029,G4030,G4031,G4032,G4033,G4034,G4035,G4036,G4037,G4038,G4039,G4040,
       G4041,G4042,G4043,G4044,G4045,G4046,G4047,G4048,G4049,G4050,G4051,G4052,G4053,G4054,G4055,G4056,G4057,G4058,G4059,G4060,
       G4061,G4062,G4063,G4064,G4065,G4066,G4067,G4068,G4069,G4070,G4071,G4072,G4073,G4074,G4075,G4076,G4077,G4078,G4079,G4080,
       G4081,G4082,G4083,G4084,G4085,G4086,G4087,G4088,G4089,G4090,G4091,G4092,G4093,G4094,G4095,G4096,G4097,G4098,G4099,G4100,
       G4101,G4102,G4103,G4104,G4105,G4106,G4107,G4108,G4109,G4110,G4111,G4112,G4113,G4114,G4115,G4116,G4117,G4118,G4119,G4120,
       G4121,G4122,G4123,G4124,G4125,G4126,G4127,G4128,G4129,G4130,G4131,G4132,G4133,G4134,G4135,G4136,G4137,G4138,G4139,G4140,
       G4141,G4142,G4143,G4144,G4145,G4146,G4147,G4148,G4149,G4150,G4151,G4152,G4153,G4154,G4155,G4156,G4157,G4158,G4159,G4160,
       G4161,G4162,G4163,G4164,G4165,G4166,G4167,G4168,G4169,G4170,G4171,G4172,G4173,G4174,G4175,G4176,G4177,G4178,G4179,G4180,
       G4181,G4182,G4183,G4184,G4185,G4186,G4187,G4188,G4189,G4190,G4191,G4192,G4193,G4194,G4195,G4196,G4197,G4198,G4199,G4200,
       G4201,G4202,G4203,G4204,G4205,G4206,G4207,G4208,G4209,G4210,G4211,G4212,G4213,G4214,G4215,G4216,G4217,G4218,G4219,G4220,
       G4221,G4222,G4223,G4224,G4225,G4226,G4227,G4228,G4229,G4230,G4231,G4232,G4233,G4234,G4235,G4236,G4237,G4238,G4239,G4240,
       G4241,G4242,G4243,G4244,G4245,G4246,G4247,G4248,G4249,G4250,G4251,G4252,G4253,G4254,G4255,G4256,G4257,G4258,G4259,G4260,
       G4261,G4262,G4263,G4264,G4265,G4266,G4267,G4268,G4269,G4270,G4271,G4272,G4273,G4274,G4275,G4276,G4277,G4278,G4279,G4280,
       G4281,G4282,G4283,G4284,G4285,G4286,G4287,G4288,G4289,G4290,G4291,G4292,G4293,G4294,G4295,G4296,G4297,G4298,G4299,G4300,
       G4301,G4302,G4303,G4304,G4305,G4306,G4307,G4308,G4309,G4310,G4311,G4312,G4313,G4314,G4315,G4316,G4317,G4318,G4319,G4320,
       G4321,G4322,G4323,G4324,G4325,G4326,G4327,G4328,G4329,G4330,G4331,G4332,G4333,G4334,G4335,G4336,G4337,G4338,G4339,G4340,
       G4341,G4342,G4343,G4344,G4345,G4346,G4347,G4348,G4349,G4350,G4351,G4352,G4353,G4354,G4355,G4356,G4357,G4358,G4359,G4360,
       G4361,G4362,G4363,G4364,G4365,G4366,G4367,G4368,G4369,G4370,G4371,G4372,G4373,G4374,G4375,G4376,G4377,G4378,G4379,G4380,
       G4381,G4382,G4383,G4384,G4385,G4386,G4387,G4388,G4389,G4390,G4391,G4392,G4393,G4394,G4395,G4396,G4397,G4398,G4399,G4400,
       G4401,G4402,G4403,G4404,G4405,G4406,G4407,G4408,G4409,G4410,G4411,G4412,G4413,G4414,G4415,G4416,G4417,G4418,G4419,G4420,
       G4421,G4422,G4423,G4424,G4425,G4426,G4427,G4428,G4429,G4430,G4431,G4432,G4433,G4434,G4435,G4436,G4437,G4438,G4439,G4440,
       G4441,G4442,G4443,G4444,G4445,G4446,G4447,G4448,G4449,G4450,G4451,G4452,G4453,G4454,G4455,G4456,G4457,G4458,G4459,G4460,
       G4461,G4462,G4463,G4464,G4465,G4466,G4467,G4468,G4469,G4470,G4471,G4472,G4473,G4474,G4475,G4476,G4477,G4478,G4479,G4480,
       G4481,G4482,G4483,G4484,G4485,G4486,G4487,G4488,G4489,G4490,G4491,G4492,G4493,G4494,G4495,G4496,G4497,G4498,G4499,G4500,
       G4501,G4502,G4503,G4504,G4505,G4506,G4507,G4508,G4509,G4510,G4511,G4512,G4513,G4514,G4515,G4516,G4517,G4518,G4519,G4520,
       G4521,G4522,G4523,G4524,G4525,G4526,G4527,G4528,G4529,G4530,G4531,G4532,G4533,G4534,G4535,G4536,G4537,G4538,G4539,G4540,
       G4541,G4542,G4543,G4544,G4545,G4546,G4547,G4548,G4549,G4550,G4551,G4552,G4553,G4554,G4555,G4556,G4557,G4558,G4559,G4560,
       G4561,G4562,G4563,G4564,G4565,G4566,G4567,G4568,G4569,G4570,G4571,G4572,G4573,G4574,G4575,G4576,G4577,G4578,G4579,G4580,
       G4581,G4582,G4583,G4584,G4585,G4586,G4587,G4588,G4589,G4590,G4591,G4592,G4593,G4594,G4595,G4596,G4597,G4598,G4599,G4600,
       G4601,G4602,G4603,G4604,G4605,G4606,G4607,G4608,G4609,G4610,G4611,G4612,G4613,G4614,G4615,G4616,G4617,G4618,G4619,G4620,
       G4621,G4622,G4623,G4624,G4625,G4626,G4627,G4628,G4629,G4630,G4631,G4632,G4633,G4634,G4635,G4636,G4637,G4638,G4639,G4640,
       G4641,G4642,G4643,G4644,G4645,G4646,G4647,G4648,G4649,G4650,G4651,G4652,G4653,G4654,G4655,G4656,G4657,G4658,G4659,G4660,
       G4661,G4662,G4663,G4664,G4665,G4666,G4667,G4668,G4669,G4670,G4671,G4672,G4673,G4674,G4675,G4676,G4677,G4678,G4679,G4680,
       G4681,G4682,G4683,G4684,G4685,G4686,G4687,G4688,G4689,G4690,G4691,G4692,G4693,G4694,G4695,G4696,G4697,G4698,G4699,G4700,
       G4701,G4702,G4703,G4704,G4705,G4706,G4707,G4708,G4709,G4710,G4711,G4712,G4713,G4714,G4715,G4716,G4717,G4718,G4719,G4720,
       G4721,G4722,G4723,G4724,G4725,G4726,G4727,G4728,G4729,G4730,G4731,G4732,G4733,G4734,G4735,G4736,G4737,G4738,G4739,G4740,
       G4741,G4742,G4743,G4744,G4745,G4746,G4747,G4748,G4749,G4750,G4751,G4752,G4753,G4754,G4755,G4756,G4757,G4758,G4759,G4760,
       G4761,G4762,G4763,G4764,G4765,G4766,G4767,G4768,G4769,G4770,G4771,G4772,G4773,G4774,G4775,G4776,G4777,G4778,G4779,G4780,
       G4781,G4782,G4783,G4784,G4785,G4786,G4787,G4788,G4789,G4790,G4791,G4792,G4793,G4794,G4795,G4796,G4797,G4798,G4799,G4800,
       G4801,G4802,G4803,G4804,G4805,G4806,G4807,G4808,G4809,G4810,G4811,G4812,G4813,G4814,G4815,G4816,G4817,G4818,G4819,G4820,
       G4821,G4822,G4823,G4824,G4825,G4826,G4827,G4828,G4829,G4830,G4831,G4832,G4833,G4834,G4835,G4836,G4837,G4838,G4839,G4840,
       G4841,G4842,G4843,G4844,G4845,G4846,G4847,G4848,G4849,G4850,G4851,G4852,G4853,G4854,G4855,G4856,G4857,G4858,G4859,G4860,
       G4861,G4862,G4863,G4864,G4865,G4866,G4867,G4868,G4869,G4870,G4871,G4872,G4873,G4874,G4875,G4876,G4877,G4878,G4879,G4880,
       G4881,G4882,G4883,G4884,G4885,G4886,G4887,G4888,G4889,G4890,G4891,G4892,G4893,G4894,G4895,G4896,G4897,G4898,G4899,G4900,
       G4901,G4902,G4903,G4904,G4905,G4906,G4907,G4908,G4909,G4910,G4911,G4912,G4913,G4914,G4915,G4916,G4917,G4918,G4919,G4920,
       G4921,G4922,G4923,G4924,G4925,G4926,G4927,G4928,G4929,G4930,G4931,G4932,G4933,G4934,G4935,G4936,G4937,G4938,G4939,G4940,
       G4941,G4942,G4943,G4944,G4945,G4946,G4947,G4948,G4949,G4950,G4951,G4952,G4953,G4954,G4955,G4956,G4957,G4958,G4959,G4960,
       G4961,G4962,G4963,G4964,G4965,G4966,G4967,G4968,G4969,G4970,G4971,G4972,G4973,G4974,G4975,G4976,G4977,G4978,G4979,G4980,
       G4981,G4982,G4983,G4984,G4985,G4986,G4987,G4988,G4989,G4990,G4991,G4992,G4993,G4994,G4995,G4996,G4997,G4998,G4999,G5000,
       G5001,G5002,G5003,G5004,G5005,G5006,G5007,G5008,G5009,G5010,G5011,G5012,G5013,G5014,G5015,G5016,G5017,G5018,G5019,G5020,
       G5021,G5022,G5023,G5024,G5025,G5026,G5027,G5028,G5029,G5030,G5031,G5032,G5033,G5034,G5035,G5036,G5037,G5038,G5039,G5040,
       G5041,G5042,G5043,G5044,G5045,G5046,G5047,G5048,G5049,G5050,G5051,G5052,G5053,G5054,G5055,G5056,G5057,G5058,G5059,G5060,
       G5061,G5062,G5063,G5064,G5065,G5066,G5067,G5068,G5069,G5070,G5071,G5072,G5073,G5074,G5075,G5076,G5077,G5078,G5079,G5080,
       G5081,G5082,G5083,G5084,G5085,G5086,G5087,G5088,G5089,G5090,G5091,G5092,G5093,G5094,G5095,G5096,G5097,G5098,G5099,G5100,
       G5101,G5102,G5103,G5104,G5105,G5106,G5107,G5108,G5109,G5110,G5111,G5112,G5113,G5114,G5115,G5116,G5117,G5118,G5119,G5120,
       G5121,G5122,G5123,G5124,G5125,G5126,G5127,G5128,G5129,G5130,G5131,G5132,G5133,G5134,G5135,G5136,G5137,G5138,G5139,G5140,
       G5141,G5142,G5143,G5144,G5145,G5146,G5147,G5148,G5149,G5150,G5151,G5152,G5153,G5154,G5155,G5156,G5157,G5158,G5159,G5160,
       G5161,G5162,G5163,G5164,G5165,G5166,G5167,G5168,G5169,G5170,G5171,G5172,G5173,G5174,G5175,G5176,G5177,G5178,G5179,G5180,
       G5181,G5182,G5183,G5184,G5185,G5186,G5187,G5188,G5189,G5190,G5191,G5192,G5193,G5194,G5195,G5196,G5197,G5198,G5199,G5200,
       G5201,G5202,G5203,G5204,G5205,G5206,G5207,G5208,G5209,G5210,G5211,G5212,G5213,G5214,G5215,G5216,G5217,G5218,G5219,G5220,
       G5221,G5222,G5223,G5224,G5225,G5226,G5227,G5228,G5229,G5230,G5231,G5232,G5233,G5234,G5235,G5236,G5237,G5238,G5239,G5240,
       G5241,G5242,G5243,G5244,G5245,G5246,G5247,G5248,G5249,G5250,G5251,G5252,G5253,G5254,G5255,G5256,G5257,G5258,G5259,G5260,
       G5261,G5262,G5263,G5264,G5265,G5266,G5267,G5268,G5269,G5270,G5271,G5272,G5273,G5274,G5275,G5276,G5277,G5278,G5279,G5280,
       G5281,G5282,G5283,G5284,G5285,G5286,G5287,G5288,G5289,G5290,G5291,G5292,G5293,G5294,G5295,G5296,G5297,G5298,G5299,G5300,
       G5301,G5302,G5303,G5304,G5305,G5306,G5307,G5308,G5309,G5310,G5311,G5312,G5313,G5314,G5315,G5316,G5317,G5318,G5319,G5320,
       G5321,G5322,G5323,G5324,G5325,G5326,G5327,G5328,G5329,G5330,G5331,G5332,G5333,G5334,G5335,G5336,G5337,G5338,G5339,G5340,
       G5341,G5342,G5343,G5344,G5345,G5346,G5347,G5348,G5349,G5350,G5351,G5352,G5353,G5354,G5355,G5356,G5357,G5358,G5359,G5360,
       G5361,G5362,G5363,G5364,G5365,G5366,G5367,G5368,G5369,G5370,G5371,G5372,G5373,G5374,G5375,G5376,G5377,G5378,G5379,G5380,
       G5381,G5382,G5383,G5384,G5385,G5386,G5387,G5388,G5389,G5390,G5391,G5392,G5393,G5394,G5395,G5396,G5397,G5398,G5399,G5400,
       G5401,G5402,G5403,G5404,G5405,G5406,G5407,G5408,G5409,G5410,G5411,G5412,G5413,G5414,G5415,G5416,G5417,G5418,G5419,G5420,
       G5421,G5422,G5423,G5424,G5425,G5426,G5427,G5428,G5429,G5430,G5431,G5432,G5433,G5434,G5435,G5436,G5437,G5438,G5439,G5440,
       G5441,G5442,G5443,G5444,G5445,G5446,G5447,G5448,G5449,G5450,G5451,G5452,G5453,G5454,G5455,G5456,G5457,G5458,G5459,G5460,
       G5461,G5462,G5463,G5464,G5465,G5466,G5467,G5468,G5469,G5470,G5471,G5472,G5473,G5474,G5475,G5476,G5477,G5478,G5479,G5480,
       G5481,G5482,G5483,G5484,G5485,G5486,G5487,G5488,G5489,G5490,G5491,G5492,G5493,G5494,G5495,G5496,G5497,G5498,G5499,G5500,
       G5501,G5502,G5503,G5504,G5505,G5506,G5507,G5508,G5509,G5510,G5511,G5512,G5513,G5514,G5515,G5516,G5517,G5518,G5519,G5520,
       G5521,G5522,G5523,G5524,G5525,G5526,G5527,G5528,G5529,G5530,G5531,G5532,G5533,G5534,G5535,G5536,G5537,G5538,G5539,G5540,
       G5541,G5542,G5543,G5544,G5545,G5546,G5547,G5548,G5549,G5550,G5551,G5552,G5553,G5554,G5555,G5556,G5557,G5558,G5559,G5560,
       G5561,G5562,G5563,G5564,G5565,G5566,G5567,G5568,G5569,G5570,G5571,G5572,G5573,G5574,G5575,G5576,G5577,G5578,G5579,G5580,
       G5581,G5582,G5583,G5584,G5585,G5586,G5587,G5588,G5589,G5590,G5591,G5592,G5593,G5594,G5595,G5596,G5597,G5598,G5599,G5600,
       G5601,G5602,G5603,G5604,G5605,G5606,G5607,G5608,G5609,G5610,G5611,G5612,G5613,G5614,G5615,G5616,G5617,G5618,G5619,G5620,
       G5621,G5622,G5623,G5624,G5625,G5626,G5627,G5628,G5629,G5630,G5631,G5632,G5633,G5634,G5635,G5636,G5637,G5638,G5639,G5640,
       G5641,G5642,G5643,G5644,G5645,G5646,G5647,G5648,G5649,G5650,G5651,G5652,G5653,G5654,G5655,G5656,G5657,G5658,G5659,G5660,
       G5661,G5662,G5663,G5664,G5665,G5666,G5667,G5668,G5669,G5670,G5671,G5672,G5673,G5674,G5675,G5676,G5677,G5678,G5679,G5680,
       G5681,G5682,G5683,G5684,G5685,G5686,G5687,G5688,G5689,G5690,G5691,G5692,G5693,G5694,G5695,G5696,G5697,G5698,G5699,G5700,
       G5701,G5702,G5703,G5704,G5705,G5706,G5707,G5708,G5709,G5710,G5711,G5712,G5713,G5714,G5715,G5716,G5717,G5718,G5719,G5720,
       G5721,G5722,G5723,G5724,G5725,G5726,G5727,G5728,G5729,G5730,G5731,G5732,G5733,G5734,G5735,G5736,G5737,G5738,G5739,G5740,
       G5741,G5742,G5743,G5744,G5745,G5746,G5747,G5748,G5749,G5750,G5751,G5752,G5753,G5754,G5755,G5756,G5757,G5758,G5759,G5760,
       G5761,G5762,G5763,G5764,G5765,G5766,G5767,G5768,G5769,G5770,G5771,G5772,G5773,G5774,G5775,G5776,G5777,G5778,G5779,G5780,
       G5781,G5782,G5783,G5784,G5785,G5786,G5787,G5788,G5789,G5790,G5791,G5792,G5793,G5794,G5795,G5796,G5797,G5798,G5799,G5800,
       G5801,G5802,G5803,G5804,G5805,G5806,G5807,G5808,G5809,G5810,G5811,G5812,G5813,G5814,G5815,G5816,G5817,G5818,G5819,G5820,
       G5821,G5822,G5823,G5824,G5825,G5826,G5827,G5828,G5829,G5830,G5831,G5832,G5833,G5834,G5835,G5836,G5837,G5838,G5839,G5840,
       G5841,G5842,G5843,G5844,G5845,G5846,G5847,G5848,G5849,G5850,G5851,G5852,G5853,G5854,G5855,G5856,G5857,G5858,G5859,G5860,
       G5861,G5862,G5863,G5864,G5865,G5866,G5867,G5868,G5869,G5870,G5871,G5872,G5873,G5874,G5875,G5876,G5877,G5878,G5879,G5880,
       G5881,G5882,G5883,G5884,G5885,G5886,G5887,G5888,G5889,G5890,G5891,G5892,G5893,G5894,G5895,G5896,G5897,G5898,G5899,G5900,
       G5901,G5902,G5903,G5904,G5905,G5906,G5907,G5908,G5909,G5910,G5911,G5912,G5913,G5914,G5915,G5916,G5917,G5918,G5919,G5920,
       G5921,G5922,G5923,G5924,G5925,G5926,G5927,G5928,G5929,G5930,G5931,G5932,G5933,G5934,G5935,G5936,G5937,G5938,G5939,G5940,
       G5941,G5942,G5943,G5944,G5945,G5946,G5947,G5948,G5949,G5950,G5951,G5952,G5953,G5954,G5955,G5956,G5957,G5958,G5959,G5960,
       G5961,G5962,G5963,G5964,G5965,G5966,G5967,G5968,G5969,G5970,G5971,G5972,G5973,G5974,G5975,G5976,G5977,G5978,G5979,G5980,
       G5981,G5982,G5983,G5984,G5985,G5986,G5987,G5988,G5989,G5990,G5991,G5992,G5993,G5994,G5995,G5996,G5997,G5998,G5999,G6000,
       G6001,G6002,G6003,G6004,G6005,G6006,G6007,G6008,G6009,G6010,G6011,G6012,G6013,G6014,G6015,G6016,G6017,G6018,G6019,G6020,
       G6021,G6022,G6023,G6024,G6025,G6026,G6027,G6028,G6029,G6030,G6031,G6032,G6033,G6034,G6035,G6036,G6037,G6038,G6039,G6040,
       G6041,G6042,G6043,G6044,G6045,G6046,G6047,G6048,G6049,G6050,G6051,G6052,G6053,G6054,G6055,G6056,G6057,G6058,G6059,G6060,
       G6061,G6062,G6063,G6064,G6065,G6066,G6067,G6068,G6069,G6070,G6071,G6072,G6073,G6074,G6075,G6076,G6077,G6078,G6079,G6080,
       G6081,G6082,G6083,G6084,G6085,G6086,G6087,G6088,G6089,G6090,G6091,G6092,G6093,G6094,G6095,G6096,G6097,G6098,G6099,G6100,
       G6101,G6102,G6103,G6104,G6105,G6106,G6107,G6108,G6109,G6110,G6111,G6112,G6113,G6114,G6115,G6116,G6117,G6118,G6119,G6120,
       G6121,G6122,G6123,G6124,G6125,G6126,G6127,G6128,G6129,G6130,G6131,G6132,G6133,G6134,G6135,G6136,G6137,G6138,G6139,G6140,
       G6141,G6142,G6143,G6144,G6145,G6146,G6147,G6148,G6149,G6150,G6151,G6152,G6153,G6154,G6155,G6156,G6157,G6158,G6159,G6160,
       G6161,G6162,G6163,G6164,G6165,G6166,G6167,G6168,G6169,G6170,G6171,G6172,G6173,G6174,G6175,G6176,G6177,G6178,G6179,G6180,
       G6181,G6182,G6183,G6184,G6185,G6186,G6187,G6188,G6189,G6190,G6191,G6192,G6193,G6194,G6195,G6196,G6197,G6198,G6199,G6200,
       G6201,G6202,G6203,G6204,G6205,G6206,G6207,G6208,G6209,G6210,G6211,G6212,G6213,G6214,G6215,G6216,G6217,G6218,G6219,G6220,
       G6221,G6222,G6223,G6224,G6225,G6226,G6227,G6228,G6229,G6230,G6231,G6232,G6233,G6234,G6235,G6236,G6237,G6238,G6239,G6240,
       G6241,G6242,G6243,G6244,G6245,G6246,G6247,G6248,G6249,G6250,G6251,G6252,G6253,G6254,G6255,G6256,G6257,G6258,G6259,G6260,
       G6261,G6262,G6263,G6264,G6265,G6266,G6267,G6268,G6269,G6270,G6271,G6272,G6273,G6274,G6275,G6276,G6277,G6278,G6279,G6280,
       G6281,G6282,G6283,G6284,G6285,G6286,G6287,G6288,G6289,G6290,G6291,G6292,G6293,G6294,G6295,G6296,G6297,G6298,G6299,G6300,
       G6301,G6302,G6303,G6304,G6305,G6306,G6307,G6308,G6309,G6310,G6311,G6312,G6313,G6314,G6315,G6316,G6317,G6318,G6319,G6320,
       G6321,G6322,G6323,G6324,G6325,G6326,G6327,G6328,G6329,G6330,G6331,G6332,G6333,G6334,G6335,G6336,G6337,G6338,G6339,G6340,
       G6341,G6342,G6343,G6344,G6345,G6346,G6347,G6348,G6349,G6350,G6351,G6352,G6353,G6354,G6355,G6356,G6357,G6358,G6359,G6360,
       G6361,G6362,G6363,G6364,G6365,G6366,G6367,G6368,G6369,G6370,G6371,G6372,G6373,G6374,G6375,G6376,G6377,G6378,G6379,G6380,
       G6381,G6382,G6383,G6384,G6385,G6386,G6387,G6388,G6389,G6390,G6391,G6392,G6393,G6394,G6395,G6396,G6397,G6398,G6399,G6400,
       G6401,G6402,G6403,G6404,G6405,G6406,G6407,G6408,G6409,G6410,G6411,G6412,G6413,G6414,G6415,G6416,G6417,G6418,G6419,G6420,
       G6421,G6422,G6423,G6424,G6425,G6426,G6427,G6428,G6429,G6430,G6431,G6432,G6433,G6434,G6435,G6436,G6437,G6438,G6439,G6440,
       G6441,G6442,G6443,G6444,G6445,G6446,G6447,G6448,G6449,G6450,G6451,G6452,G6453,G6454,G6455,G6456,G6457,G6458,G6459,G6460,
       G6461,G6462,G6463,G6464,G6465,G6466,G6467,G6468,G6469,G6470,G6471,G6472,G6473,G6474,G6475,G6476,G6477,G6478,G6479,G6480,
       G6481,G6482,G6483,G6484,G6485,G6486,G6487,G6488,G6489,G6490,G6491,G6492,G6493,G6494,G6495,G6496,G6497,G6498,G6499,G6500,
       G6501,G6502,G6503,G6504,G6505,G6506,G6507,G6508,G6509,G6510,G6511,G6512,G6513,G6514,G6515,G6516,G6517,G6518,G6519,G6520,
       G6521,G6522,G6523,G6524,G6525,G6526,G6527,G6528,G6529,G6530,G6531,G6532,G6533,G6534,G6535,G6536,G6537,G6538,G6539,G6540,
       G6541,G6542,G6543,G6544,G6545,G6546,G6547,G6548,G6549,G6550,G6551,G6552,G6553,G6554,G6555,G6556,G6557,G6558,G6559,G6560,
       G6561,G6562,G6563,G6564,G6565,G6566,G6567,G6568,G6569,G6570,G6571,G6572,G6573,G6574,G6575,G6576,G6577,G6578,G6579,G6580,
       G6581,G6582,G6583,G6584,G6585,G6586,G6587,G6588,G6589,G6590,G6591,G6592,G6593,G6594,G6595,G6596,G6597,G6598,G6599,G6600,
       G6601,G6602,G6603,G6604,G6605,G6606,G6607,G6608,G6609,G6610,G6611,G6612,G6613,G6614,G6615,G6616,G6617,G6618,G6619,G6620,
       G6621,G6622,G6623,G6624,G6625,G6626,G6627,G6628,G6629,G6630,G6631,G6632,G6633,G6634,G6635,G6636,G6637,G6638,G6639,G6640,
       G6641,G6642,G6643,G6644,G6645,G6646,G6647,G6648,G6649,G6650,G6651,G6652,G6653,G6654,G6655,G6656,G6657,G6658,G6659,G6660,
       G6661,G6662,G6663,G6664,G6665,G6666,G6667,G6668,G6669,G6670,G6671,G6672,G6673,G6674,G6675,G6676,G6677,G6678,G6679,G6680,
       G6681,G6682,G6683,G6684,G6685,G6686,G6687,G6688,G6689,G6690,G6691,G6692,G6693,G6694,G6695,G6696,G6697,G6698,G6699,G6700,
       G6701,G6702,G6703,G6704,G6705,G6706,G6707,G6708,G6709,G6710,G6711,G6712,G6713,G6714,G6715,G6716,G6717,G6718,G6719,G6720,
       G6721,G6722,G6723,G6724,G6725,G6726,G6727,G6728,G6729,G6730,G6731,G6732,G6733,G6734,G6735,G6736,G6737,G6738,G6739,G6740,
       G6741,G6742,G6743,G6744,G6745,G6746,G6747,G6748,G6749,G6750,G6751,G6752,G6753,G6754,G6755,G6756,G6757,G6758,G6759,G6760,
       G6761,G6762,G6763,G6764,G6765,G6766,G6767,G6768,G6769,G6770,G6771,G6772,G6773,G6774,G6775,G6776,G6777,G6778,G6779,G6780,
       G6781,G6782,G6783,G6784,G6785,G6786,G6787,G6788,G6789,G6790,G6791,G6792,G6793,G6794,G6795,G6796,G6797,G6798,G6799,G6800,
       G6801,G6802,G6803,G6804,G6805,G6806,G6807,G6808,G6809,G6810,G6811,G6812,G6813,G6814,G6815,G6816,G6817,G6818,G6819,G6820,
       G6821,G6822,G6823,G6824,G6825,G6826,G6827,G6828,G6829,G6830,G6831,G6832,G6833,G6834,G6835,G6836,G6837,G6838,G6839,G6840,
       G6841,G6842,G6843,G6844,G6845,G6846,G6847,G6848,G6849,G6850,G6851,G6852,G6853,G6854,G6855,G6856,G6857,G6858,G6859,G6860,
       G6861,G6862,G6863,G6864,G6865,G6866,G6867,G6868,G6869,G6870,G6871,G6872,G6873,G6874,G6875,G6876,G6877,G6878,G6879,G6880,
       G6881,G6882,G6883,G6884,G6885,G6886,G6887,G6888,G6889,G6890,G6891,G6892,G6893,G6894,G6895,G6896,G6897,G6898,G6899,G6900,
       G6901,G6902,G6903,G6904,G6905,G6906,G6907,G6908,G6909,G6910,G6911,G6912,G6913,G6914,G6915,G6916,G6917,G6918,G6919,G6920,
       G6921,G6922,G6923,G6924,G6925,G6926,G6927,G6928,G6929,G6930,G6931,G6932,G6933,G6934,G6935,G6936,G6937,G6938,G6939,G6940,
       G6941,G6942,G6943,G6944,G6945,G6946,G6947,G6948,G6949,G6950,G6951,G6952,G6953,G6954,G6955,G6956,G6957,G6958,G6959,G6960,
       G6961,G6962,G6963,G6964,G6965,G6966,G6967,G6968,G6969,G6970,G6971,G6972,G6973,G6974,G6975,G6976,G6977,G6978,G6979,G6980,
       G6981,G6982,G6983,G6984,G6985,G6986,G6987,G6988,G6989,G6990,G6991,G6992,G6993,G6994,G6995,G6996,G6997,G6998,G6999,G7000,
       G7001,G7002,G7003,G7004,G7005,G7006,G7007,G7008,G7009,G7010,G7011,G7012,G7013,G7014,G7015,G7016,G7017,G7018,G7019,G7020,
       G7021,G7022,G7023,G7024,G7025,G7026,G7027,G7028,G7029,G7030,G7031,G7032,G7033,G7034,G7035,G7036,G7037,G7038,G7039,G7040,
       G7041,G7042,G7043,G7044,G7045,G7046,G7047,G7048,G7049,G7050,G7051,G7052,G7053,G7054,G7055,G7056,G7057,G7058,G7059,G7060,
       G7061,G7062,G7063,G7064,G7065,G7066,G7067,G7068,G7069,G7070,G7071,G7072,G7073,G7074,G7075,G7076,G7077,G7078,G7079,G7080,
       G7081,G7082,G7083,G7084,G7085,G7086,G7087,G7088,G7089,G7090,G7091,G7092,G7093,G7094,G7095,G7096,G7097,G7098,G7099,G7100,
       G7101,G7102,G7103,G7104,G7105,G7106,G7107,G7108,G7109,G7110,G7111,G7112,G7113,G7114,G7115,G7116,G7117,G7118,G7119,G7120,
       G7121,G7122,G7123,G7124,G7125,G7126,G7127,G7128,G7129,G7130,G7131,G7132,G7133,G7134,G7135,G7136,G7137,G7138,G7139,G7140,
       G7141,G7142,G7143,G7144,G7145,G7146,G7147,G7148,G7149,G7150,G7151,G7152,G7153,G7154,G7155,G7156,G7157,G7158,G7159,G7160,
       G7161,G7162,G7163,G7164,G7165,G7166,G7167,G7168,G7169,G7170,G7171,G7172,G7173,G7174,G7175,G7176,G7177,G7178,G7179,G7180,
       G7181,G7182,G7183,G7184,G7185,G7186,G7187,G7188,G7189,G7190,G7191,G7192,G7193,G7194,G7195,G7196,G7197,G7198,G7199,G7200,
       G7201,G7202,G7203,G7204,G7205,G7206,G7207,G7208,G7209,G7210,G7211,G7212,G7213,G7214,G7215,G7216,G7217,G7218,G7219,G7220,
       G7221,G7222,G7223,G7224,G7225,G7226,G7227,G7228,G7229,G7230,G7231,G7232,G7233,G7234,G7235,G7236,G7237,G7238,G7239,G7240,
       G7241,G7242,G7243,G7244,G7245,G7246,G7247,G7248,G7249,G7250,G7251,G7252,G7253,G7254,G7255,G7256,G7257,G7258,G7259,G7260,
       G7261,G7262,G7263,G7264,G7265,G7266,G7267,G7268,G7269,G7270,G7271,G7272,G7273,G7274,G7275,G7276,G7277,G7278,G7279,G7280,
       G7281,G7282,G7283,G7284,G7285,G7286,G7287,G7288,G7289,G7290,G7291,G7292,G7293,G7294,G7295,G7296,G7297,G7298,G7299,G7300,
       G7301,G7302,G7303,G7304,G7305,G7306,G7307,G7308,G7309,G7310,G7311,G7312,G7313,G7314,G7315,G7316,G7317,G7318,G7319,G7320,
       G7321,G7322,G7323,G7324,G7325,G7326,G7327,G7328,G7329,G7330,G7331,G7332,G7333,G7334,G7335,G7336,G7337,G7338,G7339,G7340,
       G7341,G7342,G7343,G7344,G7345,G7346,G7347,G7348,G7349,G7350,G7351,G7352,G7353,G7354,G7355,G7356,G7357,G7358,G7359,G7360,
       G7361,G7362,G7363,G7364,G7365,G7366,G7367,G7368,G7369,G7370,G7371,G7372,G7373,G7374,G7375,G7376,G7377,G7378,G7379,G7380,
       G7381,G7382,G7383,G7384,G7385,G7386,G7387,G7388,G7389,G7390,G7391,G7392,G7393,G7394,G7395,G7396,G7397,G7398,G7399,G7400,
       G7401,G7402,G7403,G7404,G7405,G7406,G7407,G7408,G7409,G7410,G7411,G7412,G7413,G7414,G7415,G7416,G7417,G7418,G7419,G7420,
       G7421,G7422,G7423,G7424,G7425,G7426,G7427,G7428,G7429,G7430,G7431,G7432,G7433,G7434,G7435,G7436,G7437,G7438,G7439,G7440,
       G7441,G7442,G7443,G7444,G7445,G7446,G7447,G7448,G7449,G7450,G7451,G7452,G7453,G7454,G7455,G7456,G7457,G7458,G7459,G7460,
       G7461,G7462,G7463,G7464,G7465,G7466,G7467,G7468,G7469,G7470,G7471,G7472,G7473,G7474,G7475,G7476,G7477,G7478,G7479,G7480,
       G7481,G7482,G7483,G7484,G7485,G7486,G7487,G7488,G7489,G7490,G7491,G7492,G7493,G7494,G7495,G7496,G7497,G7498,G7499,G7500,
       G7501,G7502,G7503,G7504,G7505,G7506,G7507,G7508,G7509,G7510,G7511,G7512,G7513,G7514,G7515,G7516,G7517,G7518,G7519,G7520,
       G7521,G7522,G7523,G7524,G7525,G7526,G7527,G7528,G7529,G7530,G7531,G7532,G7533,G7534,G7535,G7536,G7537,G7538,G7539,G7540,
       G7541,G7542,G7543,G7544,G7545,G7546,G7547,G7548,G7549,G7550,G7551,G7552,G7553,G7554,G7555,G7556,G7557,G7558,G7559,G7560,
       G7561,G7562,G7563,G7564,G7565,G7566,G7567,G7568,G7569,G7570,G7571,G7572,G7573,G7574,G7575,G7576,G7577,G7578,G7579,G7580,
       G7581,G7582,G7583,G7584,G7585,G7586,G7587,G7588,G7589,G7590,G7591,G7592,G7593,G7594,G7595,G7596,G7597,G7598,G7599,G7600,
       G7601,G7602,G7603,G7604,G7605,G7606,G7607,G7608,G7609,G7610,G7611,G7612,G7613,G7614,G7615,G7616,G7617,G7618,G7619,G7620,
       G7621,G7622,G7623,G7624,G7625,G7626,G7627,G7628,G7629,G7630,G7631,G7632,G7633,G7634,G7635,G7636,G7637,G7638,G7639,G7640,
       G7641,G7642,G7643,G7644,G7645,G7646,G7647,G7648,G7649,G7650,G7651,G7652,G7653,G7654,G7655,G7656,G7657,G7658,G7659,G7660,
       G7661,G7662,G7663,G7664,G7665,G7666,G7667,G7668,G7669,G7670,G7671,G7672,G7673,G7674,G7675,G7676,G7677,G7678,G7679,G7680,
       G7681,G7682,G7683,G7684,G7685,G7686,G7687,G7688,G7689,G7690,G7691,G7692,G7693,G7694,G7695,G7696,G7697,G7698,G7699,G7700,
       G7701,G7702,G7703,G7704,G7705,G7706,G7707,G7708,G7709,G7710,G7711,G7712,G7713,G7714,G7715,G7716,G7717,G7718,G7719,G7720,
       G7721,G7722,G7723,G7724,G7725,G7726,G7727,G7728,G7729,G7730,G7731,G7732,G7733,G7734,G7735,G7736,G7737,G7738,G7739,G7740,
       G7741,G7742,G7743,G7744,G7745,G7746,G7747,G7748,G7749,G7750,G7751,G7752,G7753,G7754,G7755,G7756,G7757,G7758,G7759,G7760,
       G7761,G7762,G7763,G7764,G7765,G7766,G7767,G7768,G7769,G7770,G7771,G7772,G7773,G7774,G7775,G7776,G7777,G7778,G7779,G7780,
       G7781,G7782,G7783,G7784,G7785,G7786,G7787,G7788,G7789,G7790,G7791,G7792,G7793,G7794,G7795,G7796,G7797,G7798,G7799,G7800,
       G7801,G7802,G7803,G7804,G7805,G7806,G7807,G7808,G7809,G7810,G7811,G7812,G7813,G7814,G7815,G7816,G7817,G7818,G7819,G7820,
       G7821,G7822,G7823,G7824,G7825,G7826,G7827,G7828,G7829,G7830,G7831,G7832,G7833,G7834,G7835,G7836,G7837,G7838,G7839,G7840,
       G7841,G7842,G7843,G7844,G7845,G7846,G7847,G7848,G7849,G7850,G7851,G7852,G7853,G7854,G7855,G7856,G7857,G7858,G7859,G7860,
       G7861,G7862,G7863,G7864,G7865,G7866,G7867,G7868,G7869,G7870,G7871,G7872,G7873,G7874,G7875,G7876,G7877,G7878,G7879,G7880,
       G7881,G7882,G7883,G7884,G7885,G7886,G7887,G7888,G7889,G7890,G7891,G7892,G7893,G7894,G7895,G7896,G7897,G7898,G7899,G7900,
       G7901,G7902,G7903,G7904,G7905,G7906,G7907,G7908,G7909,G7910,G7911,G7912,G7913,G7914,G7915,G7916,G7917,G7918,G7919,G7920,
       G7921,G7922,G7923,G7924,G7925,G7926,G7927,G7928,G7929,G7930,G7931,G7932,G7933,G7934,G7935,G7936,G7937,G7938,G7939,G7940,
       G7941,G7942,G7943,G7944,G7945,G7946,G7947,G7948,G7949,G7950,G7951,G7952,G7953,G7954,G7955,G7956,G7957,G7958,G7959,G7960,
       G7961,G7962,G7963,G7964,G7965,G7966,G7967,G7968,G7969,G7970,G7971,G7972,G7973,G7974,G7975,G7976,G7977,G7978,G7979,G7980,
       G7981,G7982,G7983,G7984,G7985,G7986,G7987,G7988,G7989,G7990,G7991,G7992,G7993,G7994,G7995,G7996,G7997,G7998,G7999,G8000,
       G8001,G8002,G8003,G8004,G8005,G8006,G8007,G8008,G8009,G8010,G8011,G8012,G8013,G8014,G8015,G8016,G8017,G8018,G8019,G8020,
       G8021,G8022,G8023,G8024,G8025,G8026,G8027,G8028,G8029,G8030,G8031,G8032,G8033,G8034,G8035,G8036,G8037,G8038,G8039,G8040,
       G8041,G8042,G8043,G8044,G8045,G8046,G8047,G8048,G8049,G8050,G8051,G8052,G8053,G8054,G8055,G8056,G8057,G8058,G8059,G8060,
       G8061,G8062,G8063,G8064,G8065,G8066,G8067,G8068,G8069,G8070,G8071,G8072,G8073,G8074,G8075,G8076,G8077,G8078,G8079,G8080,
       G8081,G8082,G8083,G8084,G8085,G8086,G8087,G8088,G8089,G8090,G8091,G8092,G8093,G8094,G8095,G8096,G8097,G8098,G8099,G8100,
       G8101,G8102,G8103,G8104,G8105,G8106,G8107,G8108,G8109,G8110,G8111,G8112,G8113,G8114,G8115,G8116,G8117,G8118,G8119,G8120,
       G8121,G8122,G8123,G8124,G8125,G8126,G8127,G8128,G8129,G8130,G8131,G8132,G8133,G8134,G8135,G8136,G8137,G8138,G8139,G8140,
       G8141,G8142,G8143,G8144,G8145,G8146,G8147,G8148,G8149,G8150,G8151,G8152,G8153,G8154,G8155,G8156,G8157,G8158,G8159,G8160,
       G8161,G8162,G8163,G8164,G8165,G8166,G8167,G8168,G8169,G8170,G8171,G8172,G8173,G8174,G8175,G8176,G8177,G8178,G8179,G8180,
       G8181,G8182,G8183,G8184,G8185,G8186,G8187,G8188,G8189,G8190,G8191,G8192,G8193,G8194,G8195,G8196,G8197,G8198,G8199,G8200,
       G8201,G8202,G8203,G8204,G8205,G8206,G8207,G8208,G8209,G8210,G8211,G8212,G8213,G8214,G8215,G8216,G8217,G8218,G8219,G8220,
       G8221,G8222,G8223,G8224,G8225,G8226,G8227,G8228,G8229,G8230,G8231,G8232,G8233,G8234,G8235,G8236,G8237,G8238,G8239,G8240,
       G8241,G8242,G8243,G8244,G8245,G8246,G8247,G8248,G8249,G8250,G8251,G8252,G8253,G8254,G8255,G8256,G8257,G8258,G8259,G8260,
       G8261,G8262,G8263,G8264,G8265,G8266,G8267,G8268,G8269,G8270,G8271,G8272,G8273,G8274,G8275,G8276,G8277,G8278,G8279,G8280,
       G8281,G8282,G8283,G8284,G8285,G8286,G8287,G8288,G8289,G8290,G8291,G8292,G8293,G8294,G8295,G8296,G8297,G8298,G8299,G8300,
       G8301,G8302,G8303,G8304,G8305,G8306,G8307,G8308,G8309,G8310,G8311,G8312,G8313,G8314,G8315,G8316,G8317,G8318,G8319,G8320,
       G8321,G8322,G8323,G8324,G8325,G8326,G8327,G8328,G8329,G8330,G8331,G8332,G8333,G8334,G8335,G8336,G8337,G8338,G8339,G8340,
       G8341,G8342,G8343,G8344,G8345,G8346,G8347,G8348,G8349,G8350,G8351,G8352,G8353,G8354,G8355,G8356,G8357,G8358,G8359,G8360,
       G8361,G8362,G8363,G8364,G8365,G8366,G8367,G8368,G8369,G8370,G8371,G8372,G8373,G8374,G8375,G8376,G8377,G8378,G8379,G8380,
       G8381,G8382,G8383,G8384,G8385,G8386,G8387,G8388,G8389,G8390,G8391,G8392,G8393,G8394,G8395,G8396,G8397,G8398,G8399,G8400,
       G8401,G8402,G8403,G8404,G8405,G8406,G8407,G8408,G8409,G8410,G8411,G8412,G8413,G8414,G8415,G8416,G8417,G8418,G8419,G8420,
       G8421,G8422,G8423,G8424,G8425,G8426,G8427,G8428,G8429,G8430,G8431,G8432,G8433,G8434,G8435,G8436,G8437,G8438,G8439,G8440,
       G8441,G8442,G8443,G8444,G8445,G8446,G8447,G8448,G8449,G8450,G8451,G8452,G8453,G8454,G8455,G8456,G8457,G8458,G8459,G8460,
       G8461,G8462,G8463,G8464,G8465,G8466,G8467,G8468,G8469,G8470,G8471,G8472,G8473,G8474,G8475,G8476,G8477,G8478,G8479,G8480,
       G8481,G8482,G8483,G8484,G8485,G8486,G8487,G8488,G8489,G8490,G8491,G8492,G8493,G8494,G8495,G8496,G8497,G8498,G8499,G8500,
       G8501,G8502,G8503,G8504,G8505,G8506,G8507,G8508,G8509,G8510,G8511,G8512,G8513,G8514,G8515,G8516,G8517,G8518,G8519,G8520,
       G8521,G8522,G8523,G8524,G8525,G8526,G8527,G8528,G8529,G8530,G8531,G8532,G8533,G8534,G8535,G8536,G8537,G8538,G8539,G8540,
       G8541,G8542,G8543,G8544,G8545,G8546,G8547,G8548,G8549,G8550,G8551,G8552,G8553,G8554,G8555,G8556,G8557,G8558,G8559,G8560,
       G8561,G8562,G8563,G8564,G8565,G8566,G8567,G8568,G8569,G8570,G8571,G8572,G8573,G8574,G8575,G8576,G8577,G8578,G8579,G8580,
       G8581,G8582,G8583,G8584,G8585,G8586,G8587,G8588,G8589,G8590,G8591,G8592,G8593,G8594,G8595,G8596,G8597,G8598,G8599,G8600,
       G8601,G8602,G8603,G8604,G8605,G8606,G8607,G8608,G8609,G8610,G8611,G8612,G8613,G8614,G8615,G8616,G8617,G8618,G8619,G8620,
       G8621,G8622,G8623,G8624,G8625,G8626,G8627,G8628,G8629,G8630,G8631,G8632,G8633,G8634,G8635,G8636,G8637,G8638,G8639,G8640,
       G8641,G8642,G8643,G8644,G8645,G8646,G8647,G8648,G8649,G8650,G8651,G8652,G8653,G8654,G8655,G8656,G8657,G8658,G8659,G8660,
       G8661,G8662,G8663,G8664,G8665,G8666,G8667,G8668,G8669,G8670,G8671,G8672,G8673,G8674,G8675,G8676,G8677,G8678,G8679,G8680,
       G8681,G8682,G8683,G8684,G8685,G8686,G8687,G8688,G8689,G8690,G8691,G8692,G8693,G8694,G8695,G8696,G8697,G8698,G8699,G8700,
       G8701,G8702,G8703,G8704,G8705,G8706,G8707,G8708,G8709,G8710,G8711,G8712,G8713,G8714,G8715,G8716,G8717,G8718,G8719,G8720,
       G8721,G8722,G8723,G8724,G8725,G8726,G8727,G8728,G8729,G8730,G8731,G8732,G8733,G8734,G8735,G8736,G8737,G8738,G8739,G8740,
       G8741,G8742,G8743,G8744,G8745,G8746,G8747,G8748,G8749,G8750,G8751,G8752,G8753,G8754,G8755,G8756,G8757,G8758,G8759,G8760,
       G8761,G8762,G8763,G8764,G8765,G8766,G8767,G8768,G8769,G8770,G8771,G8772,G8773,G8774,G8775,G8776,G8777,G8778,G8779,G8780,
       G8781,G8782,G8783,G8784,G8785,G8786,G8787,G8788,G8789,G8790,G8791,G8792,G8793,G8794,G8795,G8796,G8797,G8798,G8799,G8800,
       G8801,G8802,G8803,G8804,G8805,G8806,G8807,G8808,G8809,G8810,G8811,G8812,G8813,G8814,G8815,G8816,G8817,G8818,G8819,G8820,
       G8821,G8822,G8823,G8824,G8825,G8826,G8827,G8828,G8829,G8830,G8831,G8832,G8833,G8834,G8835,G8836,G8837,G8838,G8839,G8840,
       G8841,G8842,G8843,G8844,G8845,G8846,G8847,G8848,G8849,G8850,G8851,G8852,G8853,G8854,G8855,G8856,G8857,G8858,G8859,G8860,
       G8861,G8862,G8863,G8864,G8865,G8866,G8867,G8868,G8869,G8870,G8871,G8872,G8873,G8874,G8875,G8876,G8877,G8878,G8879,G8880,
       G8881,G8882,G8883,G8884,G8885,G8886,G8887,G8888,G8889,G8890,G8891,G8892,G8893,G8894,G8895,G8896,G8897,G8898,G8899,G8900,
       G8901,G8902,G8903,G8904,G8905,G8906,G8907,G8908,G8909,G8910,G8911,G8912,G8913,G8914,G8915,G8916,G8917,G8918,G8919,G8920,
       G8921,G8922,G8923,G8924,G8925,G8926,G8927,G8928,G8929,G8930,G8931,G8932,G8933,G8934,G8935,G8936,G8937,G8938,G8939,G8940,
       G8941,G8942,G8943,G8944,G8945,G8946,G8947,G8948,G8949,G8950,G8951,G8952,G8953,G8954,G8955,G8956,G8957,G8958,G8959,G8960,
       G8961,G8962,G8963,G8964,G8965,G8966,G8967,G8968,G8969,G8970,G8971,G8972,G8973,G8974,G8975,G8976,G8977,G8978,G8979,G8980,
       G8981,G8982,G8983,G8984,G8985,G8986,G8987,G8988,G8989,G8990,G8991,G8992,G8993,G8994,G8995,G8996,G8997,G8998,G8999,G9000,
       G9001,G9002,G9003,G9004,G9005,G9006,G9007,G9008,G9009,G9010,G9011,G9012,G9013,G9014,G9015,G9016,G9017,G9018,G9019,G9020,
       G9021,G9022,G9023,G9024,G9025,G9026,G9027,G9028,G9029,G9030,G9031,G9032,G9033,G9034,G9035,G9036,G9037,G9038,G9039,G9040,
       G9041,G9042,G9043,G9044,G9045,G9046,G9047,G9048,G9049,G9050,G9051,G9052,G9053,G9054,G9055,G9056,G9057,G9058,G9059,G9060,
       G9061,G9062,G9063,G9064,G9065,G9066,G9067,G9068,G9069,G9070,G9071,G9072,G9073,G9074,G9075,G9076,G9077,G9078,G9079,G9080,
       G9081,G9082,G9083,G9084,G9085,G9086,G9087,G9088,G9089,G9090,G9091,G9092,G9093,G9094,G9095,G9096,G9097,G9098,G9099,G9100,
       G9101,G9102,G9103,G9104,G9105,G9106,G9107,G9108,G9109,G9110,G9111,G9112,G9113,G9114,G9115,G9116,G9117,G9118,G9119,G9120,
       G9121,G9122,G9123,G9124,G9125,G9126,G9127,G9128,G9129,G9130,G9131,G9132,G9133,G9134,G9135,G9136,G9137,G9138,G9139,G9140,
       G9141,G9142,G9143,G9144,G9145,G9146,G9147,G9148,G9149,G9150,G9151,G9152,G9153,G9154,G9155,G9156,G9157,G9158,G9159,G9160,
       G9161,G9162,G9163,G9164,G9165,G9166,G9167,G9168,G9169,G9170,G9171,G9172,G9173,G9174,G9175,G9176,G9177,G9178,G9179,G9180,
       G9181,G9182,G9183,G9184,G9185,G9186,G9187,G9188,G9189,G9190,G9191,G9192,G9193,G9194,G9195,G9196,G9197,G9198,G9199,G9200,
       G9201,G9202,G9203,G9204,G9205,G9206,G9207,G9208,G9209,G9210,G9211,G9212,G9213,G9214,G9215,G9216,G9217,G9218,G9219,G9220,
       G9221,G9222,G9223,G9224,G9225,G9226,G9227,G9228,G9229,G9230,G9231,G9232,G9233,G9234,G9235,G9236,G9237,G9238,G9239,G9240,
       G9241,G9242,G9243,G9244,G9245,G9246,G9247,G9248,G9249,G9250,G9251,G9252,G9253,G9254,G9255,G9256,G9257,G9258,G9259,G9260,
       G9261,G9262,G9263,G9264,G9265,G9266,G9267,G9268,G9269,G9270,G9271,G9272,G9273,G9274,G9275,G9276,G9277,G9278,G9279,G9280,
       G9281,G9282,G9283,G9284,G9285,G9286,G9287,G9288,G9289,G9290,G9291,G9292,G9293,G9294,G9295,G9296,G9297,G9298,G9299,G9300,
       G9301,G9302,G9303,G9304,G9305,G9306,G9307,G9308,G9309,G9310,G9311,G9312,G9313,G9314,G9315,G9316,G9317,G9318,G9319,G9320,
       G9321,G9322,G9323,G9324,G9325,G9326,G9327,G9328,G9329,G9330,G9331,G9332,G9333,G9334,G9335,G9336,G9337,G9338,G9339,G9340,
       G9341,G9342,G9343,G9344,G9345,G9346,G9347,G9348,G9349,G9350,G9351,G9352,G9353,G9354,G9355,G9356,G9357,G9358,G9359,G9360,
       G9361,G9362,G9363,G9364,G9365,G9366,G9367,G9368,G9369,G9370,G9371,G9372,G9373,G9374,G9375,G9376,G9377,G9378,G9379,G9380,
       G9381,G9382,G9383,G9384,G9385,G9386,G9387,G9388,G9389,G9390,G9391,G9392,G9393,G9394,G9395,G9396,G9397,G9398,G9399,G9400,
       G9401,G9402,G9403,G9404,G9405,G9406,G9407,G9408,G9409,G9410,G9411,G9412,G9413,G9414,G9415,G9416,G9417,G9418,G9419,G9420,
       G9421,G9422,G9423,G9424,G9425,G9426,G9427,G9428,G9429,G9430,G9431,G9432,G9433,G9434,G9435,G9436,G9437,G9438,G9439,G9440,
       G9441,G9442,G9443,G9444,G9445,G9446,G9447,G9448,G9449,G9450,G9451,G9452,G9453,G9454,G9455,G9456,G9457,G9458,G9459,G9460,
       G9461,G9462,G9463,G9464,G9465,G9466,G9467,G9468,G9469,G9470,G9471,G9472,G9473,G9474,G9475,G9476,G9477,G9478,G9479,G9480,
       G9481,G9482,G9483,G9484,G9485,G9486,G9487,G9488,G9489,G9490,G9491,G9492,G9493,G9494,G9495,G9496,G9497,G9498,G9499,G9500,
       G9501,G9502,G9503,G9504,G9505,G9506,G9507,G9508,G9509,G9510,G9511,G9512,G9513,G9514,G9515,G9516,G9517,G9518,G9519,G9520,
       G9521,G9522,G9523,G9524,G9525,G9526,G9527,G9528,G9529,G9530,G9531,G9532,G9533,G9534,G9535,G9536,G9537,G9538,G9539,G9540,
       G9541,G9542,G9543,G9544,G9545,G9546,G9547,G9548,G9549,G9550,G9551,G9552,G9553,G9554,G9555,G9556,G9557,G9558,G9559,G9560,
       G9561,G9562,G9563,G9564,G9565,G9566,G9567,G9568,G9569,G9570,G9571,G9572,G9573,G9574,G9575,G9576,G9577,G9578,G9579,G9580,
       G9581,G9582,G9583,G9584,G9585,G9586,G9587,G9588,G9589,G9590,G9591,G9592,G9593,G9594,G9595,G9596,G9597,G9598,G9599,G9600,
       G9601,G9602,G9603,G9604,G9605,G9606,G9607,G9608,G9609,G9610,G9611,G9612,G9613,G9614,G9615,G9616,G9617,G9618,G9619,G9620,
       G9621,G9622,G9623,G9624,G9625,G9626,G9627,G9628,G9629,G9630,G9631,G9632,G9633,G9634,G9635,G9636,G9637,G9638,G9639,G9640,
       G9641,G9642,G9643,G9644,G9645,G9646,G9647,G9648,G9649,G9650,G9651,G9652,G9653,G9654,G9655,G9656,G9657,G9658,G9659,G9660,
       G9661,G9662,G9663,G9664,G9665,G9666,G9667,G9668,G9669,G9670,G9671,G9672,G9673,G9674,G9675,G9676,G9677,G9678,G9679,G9680,
       G9681,G9682,G9683,G9684,G9685,G9686,G9687,G9688,G9689,G9690,G9691,G9692,G9693,G9694,G9695,G9696,G9697,G9698,G9699,G9700,
       G9701,G9702,G9703,G9704,G9705,G9706,G9707,G9708,G9709,G9710,G9711,G9712,G9713,G9714,G9715,G9716,G9717,G9718,G9719,G9720,
       G9721,G9722,G9723,G9724,G9725,G9726,G9727,G9728,G9729,G9730,G9731,G9732,G9733,G9734,G9735,G9736,G9737,G9738,G9739,G9740,
       G9741,G9742,G9743,G9744,G9745,G9746,G9747,G9748,G9749,G9750,G9751,G9752,G9753,G9754,G9755,G9756,G9757,G9758,G9759,G9760,
       G9761,G9762,G9763,G9764,G9765,G9766,G9767,G9768,G9769,G9770,G9771,G9772,G9773,G9774,G9775,G9776,G9777,G9778,G9779,G9780,
       G9781,G9782,G9783,G9784,G9785,G9786,G9787,G9788,G9789,G9790,G9791,G9792,G9793,G9794,G9795,G9796,G9797,G9798,G9799,G9800,
       G9801,G9802,G9803,G9804,G9805,G9806,G9807,G9808,G9809,G9810,G9811,G9812,G9813,G9814,G9815,G9816,G9817,G9818,G9819,G9820,
       G9821,G9822,G9823,G9824,G9825,G9826,G9827,G9828,G9829,G9830,G9831,G9832,G9833,G9834,G9835,G9836,G9837,G9838,G9839,G9840,
       G9841,G9842,G9843,G9844,G9845,G9846,G9847,G9848,G9849,G9850,G9851,G9852,G9853,G9854,G9855,G9856,G9857,G9858,G9859,G9860,
       G9861,G9862,G9863,G9864,G9865,G9866,G9867,G9868,G9869,G9870,G9871,G9872,G9873,G9874,G9875,G9876,G9877,G9878,G9879,G9880,
       G9881,G9882,G9883,G9884,G9885,G9886,G9887,G9888,G9889,G9890,G9891,G9892,G9893,G9894,G9895,G9896,G9897,G9898,G9899,G9900,
       G9901,G9902,G9903,G9904,G9905,G9906,G9907,G9908,G9909,G9910,G9911,G9912,G9913,G9914,G9915,G9916,G9917,G9918,G9919,G9920,
       G9921,G9922,G9923,G9924,G9925,G9926,G9927,G9928,G9929,G9930,G9931,G9932,G9933,G9934,G9935,G9936,G9937,G9938,G9939,G9940,
       G9941,G9942,G9943,G9944,G9945,G9946,G9947,G9948,G9949,G9950,G9951,G9952,G9953,G9954,G9955,G9956,G9957,G9958,G9959,G9960,
       G9961,G9962,G9963,G9964,G9965,G9966,G9967,G9968,G9969,G9970,G9971,G9972,G9973,G9974,G9975,G9976,G9977,G9978,G9979,G9980,
       G9981,G9982,G9983,G9984,G9985,G9986,G9987,G9988,G9989,G9990,G9991,G9992,G9993,G9994,G9995,G9996,G9997,G9998,G9999,G10000,
       G10001,G10002,G10003,G10004,G10005,G10006,G10007,G10008,G10009,G10010,G10011,G10012,G10013,G10014,G10015,G10016,G10017,G10018,G10019,G10020,
       G10021,G10022,G10023,G10024,G10025,G10026,G10027,G10028,G10029,G10030,G10031,G10032,G10033,G10034,G10035,G10036,G10037,G10038,G10039,G10040,
       G10041,G10042,G10043,G10044,G10045,G10046,G10047,G10048,G10049,G10050,G10051,G10052,G10053,G10054,G10055,G10056,G10057,G10058,G10059,G10060,
       G10061,G10062,G10063,G10064,G10065,G10066,G10067,G10068,G10069,G10070,G10071,G10072,G10073,G10074,G10075,G10076,G10077,G10078,G10079,G10080,
       G10081,G10082,G10083,G10084,G10085,G10086,G10087,G10088,G10089,G10090,G10091,G10092,G10093,G10094,G10095,G10096,G10097,G10098,G10099,G10100,
       G10101,G10102,G10103,G10104,G10105,G10106,G10107,G10108,G10109,G10110,G10111,G10112,G10113,G10114,G10115,G10116,G10117,G10118,G10119,G10120,
       G10121,G10122,G10123,G10124,G10125,G10126,G10127,G10128,G10129,G10130,G10131,G10132,G10133,G10134,G10135,G10136,G10137,G10138,G10139,G10140,
       G10141,G10142,G10143,G10144,G10145,G10146,G10147,G10148,G10149,G10150,G10151,G10152,G10153,G10154,G10155,G10156,G10157,G10158,G10159,G10160,
       G10161,G10162,G10163,G10164,G10165,G10166,G10167,G10168,G10169,G10170,G10171,G10172,G10173,G10174,G10175,G10176,G10177,G10178,G10179,G10180,
       G10181,G10182,G10183,G10184,G10185,G10186,G10187,G10188,G10189,G10190,G10191,G10192,G10193,G10194,G10195,G10196,G10197,G10198,G10199,G10200,
       G10201,G10202,G10203,G10204,G10205,G10206,G10207,G10208,G10209,G10210,G10211,G10212,G10213,G10214,G10215,G10216,G10217,G10218,G10219,G10220,
       G10221,G10222,G10223,G10224,G10225,G10226,G10227,G10228,G10229,G10230,G10231,G10232,G10233,G10234,G10235,G10236,G10237,G10238,G10239,G10240,
       G10241,G10242,G10243,G10244,G10245,G10246,G10247,G10248,G10249,G10250,G10251,G10252,G10253,G10254,G10255,G10256,G10257,G10258,G10259,G10260,
       G10261,G10262,G10263,G10264,G10265,G10266,G10267,G10268,G10269,G10270,G10271,G10272,G10273,G10274,G10275,G10276,G10277,G10278,G10279,G10280,
       G10281,G10282,G10283,G10284,G10285,G10286,G10287,G10288,G10289,G10290,G10291,G10292,G10293,G10294,G10295,G10296,G10297,G10298,G10299,G10300,
       G10301,G10302,G10303,G10304,G10305,G10306,G10307,G10308,G10309,G10310,G10311,G10312,G10313,G10314,G10315,G10316,G10317,G10318,G10319,G10320,
       G10321,G10322,G10323,G10324,G10325,G10326,G10327,G10328,G10329,G10330,G10331,G10332,G10333,G10334,G10335,G10336,G10337,G10338,G10339,G10340,
       G10341,G10342,G10343,G10344,G10345,G10346,G10347,G10348,G10349,G10350,G10351,G10352,G10353,G10354,G10355,G10356,G10357,G10358,G10359,G10360,
       G10361,G10362,G10363,G10364,G10365,G10366,G10367,G10368,G10369,G10370,G10371,G10372,G10373,G10374,G10375,G10376,G10377,G10378,G10379,G10380,
       G10381,G10382,G10383,G10384,G10385,G10386,G10387,G10388,G10389,G10390,G10391,G10392,G10393,G10394,G10395,G10396,G10397,G10398,G10399,G10400,
       G10401,G10402,G10403,G10404,G10405,G10406,G10407,G10408,G10409,G10410,G10411,G10412,G10413,G10414,G10415,G10416,G10417,G10418,G10419,G10420,
       G10421,G10422,G10423,G10424,G10425,G10426,G10427,G10428,G10429,G10430,G10431,G10432,G10433,G10434,G10435,G10436,G10437,G10438,G10439,G10440,
       G10441,G10442,G10443,G10444,G10445,G10446,G10447,G10448,G10449,G10450,G10451,G10452,G10453,G10454,G10455,G10456,G10457,G10458,G10459,G10460,
       G10461,G10462,G10463,G10464,G10465,G10466,G10467,G10468,G10469,G10470,G10471,G10472,G10473,G10474,G10475,G10476,G10477,G10478,G10479,G10480,
       G10481,G10482,G10483,G10484,G10485,G10486,G10487,G10488,G10489,G10490,G10491,G10492,G10493,G10494,G10495,G10496,G10497,G10498,G10499,G10500,
       G10501,G10502,G10503,G10504,G10505,G10506,G10507,G10508,G10509,G10510,G10511,G10512,G10513,G10514,G10515,G10516,G10517,G10518,G10519,G10520,
       G10521,G10522,G10523,G10524,G10525,G10526,G10527,G10528,G10529,G10530,G10531,G10532,G10533,G10534,G10535,G10536,G10537,G10538,G10539,G10540,
       G10541,G10542,G10543,G10544,G10545,G10546,G10547,G10548,G10549,G10550,G10551,G10552,G10553,G10554,G10555,G10556,G10557,G10558,G10559,G10560,
       G10561,G10562,G10563,G10564,G10565,G10566,G10567,G10568,G10569,G10570,G10571,G10572,G10573,G10574,G10575,G10576,G10577,G10578,G10579,G10580,
       G10581,G10582,G10583,G10584,G10585,G10586,G10587,G10588,G10589,G10590,G10591,G10592,G10593,G10594,G10595,G10596,G10597,G10598,G10599,G10600,
       G10601,G10602,G10603,G10604,G10605,G10606,G10607,G10608,G10609,G10610,G10611,G10612,G10613,G10614,G10615,G10616,G10617,G10618,G10619,G10620,
       G10621,G10622,G10623,G10624,G10625,G10626,G10627,G10628,G10629,G10630,G10631,G10632,G10633,G10634,G10635,G10636,G10637,G10638,G10639,G10640,
       G10641,G10642,G10643,G10644,G10645,G10646,G10647,G10648,G10649,G10650,G10651,G10652,G10653,G10654,G10655,G10656,G10657,G10658,G10659,G10660,
       G10661,G10662,G10663,G10664,G10665,G10666,G10667,G10668,G10669,G10670,G10671,G10672,G10673,G10674,G10675,G10676,G10677,G10678,G10679,G10680,
       G10681,G10682,G10683,G10684,G10685,G10686,G10687,G10688,G10689,G10690,G10691,G10692,G10693,G10694,G10695,G10696,G10697,G10698,G10699,G10700,
       G10701,G10702,G10703,G10704,G10705,G10706,G10707,G10708,G10709,G10710,G10711,G10712,G10713,G10714,G10715,G10716,G10717,G10718,G10719,G10720,
       G10721,G10722,G10723,G10724,G10725,G10726,G10727,G10728,G10729,G10730,G10731,G10732,G10733,G10734,G10735,G10736,G10737,G10738,G10739,G10740,
       G10741,G10742,G10743,G10744,G10745,G10746,G10747,G10748,G10749,G10750,G10751,G10752,G10753,G10754,G10755,G10756,G10757,G10758,G10759,G10760,
       G10761,G10762,G10763,G10764,G10765,G10766,G10767,G10768,G10769,G10770,G10771,G10772,G10773,G10774,G10775,G10776,G10777,G10778,G10779,G10780,
       G10781,G10782,G10783,G10784,G10785,G10786,G10787,G10788,G10789,G10790,G10791,G10792,G10793,G10794,G10795,G10796,G10797,G10798,G10799,G10800,
       G10801,G10802,G10803,G10804,G10805,G10806,G10807,G10808,G10809,G10810,G10811,G10812,G10813,G10814,G10815,G10816,G10817,G10818,G10819,G10820,
       G10821,G10822,G10823,G10824,G10825,G10826,G10827,G10828,G10829,G10830,G10831,G10832,G10833,G10834,G10835,G10836,G10837,G10838,G10839,G10840,
       G10841,G10842,G10843,G10844,G10845,G10846,G10847,G10848,G10849,G10850,G10851,G10852,G10853,G10854,G10855,G10856,G10857,G10858,G10859,G10860,
       G10861,G10862,G10863,G10864,G10865,G10866,G10867,G10868,G10869,G10870,G10871,G10872,G10873,G10874,G10875,G10876,G10877,G10878,G10879,G10880,
       G10881,G10882,G10883,G10884,G10885,G10886,G10887,G10888,G10889,G10890,G10891,G10892,G10893,G10894,G10895,G10896,G10897,G10898,G10899,G10900,
       G10901,G10902,G10903,G10904,G10905,G10906,G10907,G10908,G10909,G10910,G10911,G10912,G10913,G10914,G10915,G10916,G10917,G10918,G10919,G10920,
       G10921,G10922,G10923,G10924,G10925,G10926,G10927,G10928,G10929,G10930,G10931,G10932,G10933,G10934,G10935,G10936,G10937,G10938,G10939,G10940,
       G10941,G10942,G10943,G10944,G10945,G10946,G10947,G10948,G10949,G10950,G10951,G10952,G10953,G10954,G10955,G10956,G10957,G10958,G10959,G10960,
       G10961,G10962,G10963,G10964,G10965,G10966,G10967,G10968,G10969,G10970,G10971,G10972,G10973,G10974,G10975,G10976,G10977,G10978,G10979,G10980,
       G10981,G10982,G10983,G10984,G10985,G10986,G10987,G10988,G10989,G10990,G10991,G10992,G10993,G10994,G10995,G10996,G10997,G10998,G10999,G11000,
       G11001,G11002,G11003,G11004,G11005,G11006,G11007,G11008,G11009,G11010,G11011,G11012,G11013,G11014,G11015,G11016,G11017,G11018,G11019,G11020,
       G11021,G11022,G11023,G11024,G11025,G11026,G11027,G11028,G11029,G11030,G11031,G11032,G11033,G11034,G11035,G11036,G11037,G11038,G11039,G11040,
       G11041,G11042,G11043,G11044,G11045,G11046,G11047,G11048,G11049,G11050,G11051,G11052,G11053,G11054,G11055,G11056,G11057,G11058,G11059,G11060,
       G11061,G11062,G11063,G11064,G11065,G11066,G11067,G11068,G11069,G11070,G11071,G11072,G11073,G11074,G11075,G11076,G11077,G11078,G11079,G11080,
       G11081,G11082,G11083,G11084,G11085,G11086,G11087,G11088,G11089,G11090,G11091,G11092,G11093,G11094,G11095,G11096,G11097,G11098,G11099,G11100,
       G11101,G11102,G11103,G11104,G11105,G11106,G11107,G11108,G11109,G11110,G11111,G11112,G11113,G11114,G11115,G11116,G11117,G11118,G11119,G11120,
       G11121,G11122,G11123,G11124,G11125,G11126,G11127,G11128,G11129,G11130,G11131,G11132,G11133,G11134,G11135,G11136,G11137,G11138,G11139,G11140,
       G11141,G11142,G11143,G11144,G11145,G11146,G11147,G11148,G11149,G11150,G11151,G11152,G11153,G11154,G11155,G11156,G11157,G11158,G11159,G11160,
       G11161,G11162,G11163,G11164,G11165,G11166,G11167,G11168,G11169,G11170,G11171,G11172,G11173,G11174,G11175,G11176,G11177,G11178,G11179,G11180,
       G11181,G11182,G11183,G11184,G11185,G11186,G11187,G11188,G11189,G11190,G11191,G11192,G11193,G11194,G11195,G11196,G11197,G11198,G11199,G11200,
       G11201,G11202,G11203,G11204,G11205,G11206,G11207,G11208,G11209,G11210,G11211,G11212,G11213,G11214,G11215,G11216,G11217,G11218,G11219,G11220,
       G11221,G11222,G11223,G11224,G11225,G11226,G11227,G11228,G11229,G11230,G11231,G11232,G11233,G11234,G11235,G11236,G11237,G11238,G11239,G11240,
       G11241,G11242,G11243,G11244,G11245,G11246,G11247,G11248,G11249,G11250,G11251,G11252,G11253,G11254,G11255,G11256,G11257,G11258,G11259,G11260,
       G11261,G11262,G11263,G11264,G11265,G11266,G11267,G11268,G11269,G11270,G11271,G11272,G11273,G11274,G11275,G11276,G11277,G11278,G11279,G11280,
       G11281,G11282,G11283,G11284,G11285,G11286,G11287,G11288,G11289,G11290,G11291,G11292,G11293,G11294,G11295,G11296,G11297,G11298,G11299,G11300,
       G11301,G11302,G11303,G11304,G11305,G11306,G11307,G11308,G11309,G11310,G11311,G11312,G11313,G11314,G11315,G11316,G11317,G11318,G11319,G11320,
       G11321,G11322,G11323,G11324,G11325,G11326,G11327,G11328,G11329,G11330,G11331,G11332,G11333,G11334,G11335,G11336,G11337,G11338,G11339,G11340,
       G11341,G11342,G11343,G11344,G11345,G11346,G11347,G11348,G11349,G11350,G11351,G11352,G11353,G11354,G11355,G11356,G11357,G11358,G11359,G11360,
       G11361,G11362,G11363,G11364,G11365,G11366,G11367,G11368,G11369,G11370,G11371,G11372,G11373,G11374,G11375,G11376,G11377,G11378,G11379,G11380,
       G11381,G11382,G11383,G11384,G11385,G11386,G11387,G11388,G11389,G11390,G11391,G11392,G11393,G11394,G11395,G11396,G11397,G11398,G11399,G11400,
       G11401,G11402,G11403,G11404,G11405,G11406,G11407,G11408,G11409,G11410,G11411,G11412,G11413,G11414,G11415,G11416,G11417,G11418,G11419,G11420,
       G11421,G11422,G11423,G11424,G11425,G11426,G11427,G11428,G11429,G11430,G11431,G11432,G11433,G11434,G11435,G11436,G11437,G11438,G11439,G11440,
       G11441,G11442,G11443,G11444,G11445,G11446,G11447,G11448,G11449,G11450,G11451,G11452,G11453,G11454,G11455,G11456,G11457,G11458,G11459,G11460,
       G11461,G11462,G11463,G11464,G11465,G11466,G11467,G11468,G11469,G11470,G11471,G11472,G11473,G11474,G11475,G11476,G11477,G11478,G11479,G11480,
       G11481,G11482,G11483,G11484,G11485,G11486,G11487,G11488,G11489,G11490,G11491,G11492,G11493,G11494,G11495,G11496,G11497,G11498,G11499,G11500,
       G11501,G11502,G11503,G11504,G11505,G11506,G11507,G11508,G11509,G11510,G11511,G11512,G11513,G11514,G11515,G11516,G11517,G11518,G11519,G11520,
       G11521,G11522,G11523,G11524,G11525,G11526,G11527,G11528,G11529,G11530,G11531,G11532,G11533,G11534,G11535,G11536,G11537,G11538,G11539,G11540,
       G11541,G11542,G11543,G11544,G11545,G11546,G11547,G11548,G11549,G11550,G11551,G11552,G11553,G11554,G11555,G11556,G11557,G11558,G11559,G11560,
       G11561,G11562,G11563,G11564,G11565,G11566,G11567,G11568,G11569,G11570,G11571,G11572,G11573,G11574,G11575,G11576,G11577,G11578,G11579,G11580,
       G11581,G11582,G11583,G11584,G11585,G11586,G11587,G11588,G11589,G11590,G11591,G11592,G11593,G11594,G11595,G11596,G11597,G11598,G11599,G11600,
       G11601,G11602,G11603,G11604,G11605,G11606,G11607,G11608,G11609,G11610,G11611,G11612,G11613,G11614,G11615,G11616,G11617,G11618,G11619,G11620,
       G11621,G11622,G11623,G11624,G11625,G11626,G11627,G11628,G11629,G11630,G11631,G11632,G11633,G11634,G11635,G11636,G11637,G11638,G11639,G11640,
       G11641,G11642,G11643,G11644,G11645,G11646,G11647,G11648,G11649,G11650,G11651,G11652,G11653,G11654,G11655,G11656,G11657,G11658,G11659,G11660,
       G11661,G11662,G11663,G11664,G11665,G11666,G11667,G11668,G11669,G11670,G11671,G11672,G11673,G11674,G11675,G11676,G11677,G11678,G11679,G11680,
       G11681,G11682,G11683,G11684,G11685,G11686,G11687,G11688,G11689,G11690,G11691,G11692,G11693,G11694,G11695,G11696,G11697,G11698,G11699,G11700,
       G11701,G11702,G11703,G11704,G11705,G11706,G11707,G11708,G11709,G11710,G11711,G11712,G11713,G11714,G11715,G11716,G11717,G11718,G11719,G11720,
       G11721,G11722,G11723,G11724,G11725,G11726,G11727,G11728,G11729,G11730,G11731,G11732,G11733,G11734,G11735,G11736,G11737,G11738,G11739,G11740,
       G11741,G11742,G11743,G11744,G11745,G11746,G11747,G11748,G11749,G11750,G11751,G11752,G11753,G11754,G11755,G11756,G11757,G11758,G11759,G11760,
       G11761,G11762,G11763,G11764,G11765,G11766,G11767,G11768,G11769,G11770,G11771,G11772,G11773,G11774,G11775,G11776,G11777,G11778,G11779,G11780,
       G11781,G11782,G11783,G11784,G11785,G11786,G11787,G11788,G11789,G11790,G11791,G11792,G11793,G11794,G11795,G11796,G11797,G11798,G11799,G11800,
       G11801,G11802,G11803,G11804,G11805,G11806,G11807,G11808,G11809,G11810,G11811,G11812,G11813,G11814,G11815,G11816,G11817,G11818,G11819,G11820,
       G11821,G11822,G11823,G11824,G11825,G11826,G11827,G11828,G11829,G11830,G11831,G11832,G11833,G11834,G11835,G11836,G11837,G11838,G11839,G11840,
       G11841,G11842,G11843,G11844,G11845,G11846,G11847,G11848,G11849,G11850,G11851,G11852,G11853,G11854,G11855,G11856,G11857,G11858,G11859,G11860,
       G11861,G11862,G11863,G11864,G11865,G11866,G11867,G11868,G11869,G11870,G11871,G11872,G11873,G11874,G11875,G11876,G11877,G11878,G11879,G11880,
       G11881,G11882,G11883,G11884,G11885,G11886,G11887,G11888,G11889,G11890,G11891,G11892,G11893,G11894,G11895,G11896,G11897,G11898,G11899,G11900,
       G11901,G11902,G11903,G11904,G11905,G11906,G11907,G11908,G11909,G11910,G11911,G11912,G11913,G11914,G11915,G11916,G11917,G11918,G11919,G11920,
       G11921,G11922,G11923,G11924,G11925,G11926,G11927,G11928,G11929,G11930,G11931,G11932,G11933,G11934,G11935,G11936,G11937,G11938,G11939,G11940,
       G11941,G11942,G11943,G11944,G11945,G11946,G11947,G11948,G11949,G11950,G11951,G11952,G11953,G11954,G11955,G11956,G11957,G11958,G11959,G11960,
       G11961,G11962,G11963,G11964,G11965,G11966,G11967,G11968,G11969,G11970,G11971,G11972,G11973,G11974,G11975,G11976,G11977,G11978,G11979,G11980,
       G11981,G11982,G11983,G11984,G11985,G11986,G11987,G11988,G11989,G11990,G11991,G11992,G11993,G11994,G11995,G11996,G11997,G11998,G11999,G12000,
       G12001,G12002,G12003,G12004,G12005,G12006,G12007,G12008,G12009,G12010,G12011,G12012,G12013,G12014,G12015,G12016,G12017,G12018,G12019,G12020,
       G12021,G12022,G12023,G12024,G12025,G12026,G12027,G12028,G12029,G12030,G12031,G12032,G12033,G12034,G12035,G12036,G12037,G12038,G12039,G12040,
       G12041,G12042,G12043,G12044,G12045,G12046,G12047,G12048,G12049,G12050,G12051,G12052,G12053,G12054,G12055,G12056,G12057,G12058,G12059,G12060,
       G12061,G12062,G12063,G12064,G12065,G12066,G12067,G12068,G12069,G12070,G12071,G12072,G12073,G12074,G12075,G12076,G12077,G12078,G12079,G12080,
       G12081,G12082,G12083,G12084,G12085,G12086,G12087,G12088,G12089,G12090,G12091,G12092,G12093,G12094,G12095,G12096,G12097,G12098,G12099,G12100,
       G12101,G12102,G12103,G12104,G12105,G12106,G12107,G12108,G12109,G12110,G12111,G12112,G12113,G12114,G12115,G12116,G12117,G12118,G12119,G12120,
       G12121,G12122,G12123,G12124,G12125,G12126,G12127,G12128,G12129,G12130,G12131,G12132,G12133,G12134,G12135,G12136,G12137,G12138,G12139,G12140,
       G12141,G12142,G12143,G12144,G12145,G12146,G12147,G12148,G12149,G12150,G12151,G12152,G12153,G12154,G12155,G12156,G12157,G12158,G12159,G12160,
       G12161,G12162,G12163,G12164,G12165,G12166,G12167,G12168,G12169,G12170,G12171,G12172,G12173,G12174,G12175,G12176,G12177,G12178,G12179,G12180,
       G12181,G12182,G12183,G12184,G12185,G12186,G12187,G12188,G12189,G12190,G12191,G12192,G12193,G12194,G12195,G12196,G12197,G12198,G12199,G12200,
       G12201,G12202,G12203,G12204,G12205,G12206,G12207,G12208,G12209,G12210,G12211,G12212,G12213,G12214,G12215,G12216,G12217,G12218,G12219,G12220,
       G12221,G12222,G12223,G12224,G12225,G12226,G12227,G12228,G12229,G12230,G12231,G12232,G12233,G12234,G12235,G12236,G12237,G12238,G12239,G12240,
       G12241,G12242,G12243,G12244,G12245,G12246,G12247,G12248,G12249,G12250,G12251,G12252,G12253,G12254,G12255,G12256,G12257,G12258,G12259,G12260,
       G12261,G12262,G12263,G12264,G12265,G12266,G12267,G12268,G12269,G12270,G12271,G12272,G12273,G12274,G12275,G12276,G12277,G12278,G12279,G12280,
       G12281,G12282,G12283,G12284,G12285,G12286,G12287,G12288,G12289,G12290,G12291,G12292,G12293,G12294,G12295,G12296,G12297,G12298,G12299,G12300,
       G12301,G12302,G12303,G12304,G12305,G12306,G12307,G12308,G12309,G12310,G12311,G12312,G12313,G12314,G12315,G12316,G12317,G12318,G12319,G12320,
       G12321,G12322,G12323,G12324,G12325,G12326,G12327,G12328,G12329,G12330,G12331,G12332,G12333,G12334,G12335,G12336,G12337,G12338,G12339,G12340,
       G12341,G12342,G12343,G12344,G12345,G12346,G12347,G12348,G12349,G12350,G12351,G12352,G12353,G12354,G12355,G12356,G12357,G12358,G12359,G12360,
       G12361,G12362,G12363,G12364,G12365,G12366,G12367,G12368,G12369,G12370,G12371,G12372,G12373,G12374,G12375,G12376,G12377,G12378,G12379,G12380,
       G12381,G12382,G12383,G12384,G12385,G12386,G12387,G12388,G12389,G12390,G12391,G12392,G12393,G12394,G12395,G12396,G12397,G12398,G12399,G12400,
       G12401,G12402,G12403,G12404,G12405,G12406,G12407,G12408,G12409,G12410,G12411,G12412,G12413,G12414,G12415,G12416,G12417,G12418,G12419,G12420,
       G12421,G12422,G12423,G12424,G12425,G12426,G12427,G12428,G12429,G12430,G12431,G12432,G12433,G12434,G12435,G12436,G12437,G12438,G12439,G12440,
       G12441,G12442,G12443,G12444,G12445,G12446,G12447,G12448,G12449,G12450,G12451,G12452,G12453,G12454,G12455,G12456,G12457,G12458,G12459,G12460,
       G12461,G12462,G12463,G12464,G12465,G12466,G12467,G12468,G12469,G12470,G12471,G12472,G12473,G12474,G12475,G12476,G12477,G12478,G12479,G12480,
       G12481,G12482,G12483,G12484,G12485,G12486,G12487,G12488,G12489,G12490,G12491,G12492,G12493,G12494,G12495,G12496,G12497,G12498,G12499,G12500,
       G12501,G12502,G12503,G12504,G12505,G12506,G12507,G12508,G12509,G12510,G12511,G12512,G12513,G12514,G12515,G12516,G12517,G12518,G12519,G12520,
       G12521,G12522,G12523,G12524,G12525,G12526,G12527,G12528,G12529,G12530,G12531,G12532,G12533,G12534,G12535,G12536,G12537,G12538,G12539,G12540,
       G12541,G12542,G12543,G12544,G12545,G12546,G12547,G12548,G12549,G12550,G12551,G12552,G12553,G12554,G12555,G12556,G12557,G12558,G12559,G12560,
       G12561,G12562,G12563,G12564,G12565,G12566,G12567,G12568,G12569,G12570,G12571,G12572,G12573,G12574,G12575,G12576,G12577,G12578,G12579,G12580,
       G12581,G12582,G12583,G12584,G12585,G12586,G12587,G12588,G12589,G12590,G12591,G12592,G12593,G12594,G12595,G12596,G12597,G12598,G12599,G12600,
       G12601,G12602,G12603,G12604,G12605,G12606,G12607,G12608,G12609,G12610,G12611,G12612,G12613,G12614,G12615,G12616,G12617,G12618,G12619,G12620,
       G12621,G12622,G12623,G12624,G12625,G12626,G12627,G12628,G12629,G12630,G12631,G12632,G12633,G12634,G12635,G12636,G12637,G12638,G12639,G12640,
       G12641,G12642,G12643,G12644,G12645,G12646,G12647,G12648,G12649,G12650,G12651,G12652,G12653,G12654,G12655,G12656,G12657,G12658,G12659,G12660,
       G12661,G12662,G12663,G12664,G12665,G12666,G12667,G12668,G12669,G12670,G12671,G12672,G12673,G12674,G12675,G12676,G12677,G12678,G12679,G12680,
       G12681,G12682,G12683,G12684,G12685,G12686,G12687,G12688,G12689,G12690,G12691,G12692,G12693,G12694,G12695,G12696,G12697,G12698,G12699,G12700,
       G12701,G12702,G12703,G12704,G12705,G12706,G12707,G12708,G12709,G12710,G12711,G12712,G12713,G12714,G12715,G12716,G12717,G12718,G12719,G12720,
       G12721,G12722,G12723,G12724,G12725,G12726,G12727,G12728,G12729,G12730,G12731,G12732,G12733,G12734,G12735,G12736,G12737,G12738,G12739,G12740,
       G12741,G12742,G12743,G12744,G12745,G12746,G12747,G12748,G12749,G12750,G12751,G12752,G12753,G12754,G12755,G12756,G12757,G12758,G12759,G12760,
       G12761,G12762,G12763,G12764,G12765,G12766,G12767,G12768,G12769,G12770,G12771,G12772,G12773,G12774,G12775,G12776,G12777,G12778,G12779,G12780,
       G12781,G12782,G12783,G12784,G12785,G12786,G12787,G12788,G12789,G12790,G12791,G12792,G12793,G12794,G12795,G12796,G12797,G12798,G12799,G12800,
       G12801,G12802,G12803,G12804,G12805,G12806,G12807,G12808,G12809,G12810,G12811,G12812,G12813,G12814,G12815,G12816,G12817,G12818,G12819,G12820,
       G12821,G12822,G12823,G12824,G12825,G12826,G12827,G12828,G12829,G12830,G12831,G12832,G12833,G12834,G12835,G12836,G12837,G12838,G12839,G12840,
       G12841,G12842,G12843,G12844,G12845,G12846,G12847,G12848,G12849,G12850,G12851,G12852,G12853,G12854,G12855,G12856,G12857,G12858,G12859,G12860,
       G12861,G12862,G12863,G12864,G12865,G12866,G12867,G12868,G12869,G12870,G12871,G12872,G12873,G12874,G12875,G12876,G12877,G12878,G12879,G12880,
       G12881,G12882,G12883,G12884,G12885,G12886,G12887,G12888,G12889,G12890,G12891,G12892,G12893,G12894,G12895,G12896,G12897,G12898,G12899,G12900,
       G12901,G12902,G12903,G12904,G12905,G12906,G12907,G12908,G12909,G12910,G12911,G12912,G12913,G12914,G12915,G12916,G12917,G12918,G12919,G12920,
       G12921,G12922,G12923,G12924,G12925,G12926,G12927,G12928,G12929,G12930,G12931,G12932,G12933,G12934,G12935,G12936,G12937,G12938,G12939,G12940,
       G12941,G12942,G12943,G12944,G12945,G12946,G12947,G12948,G12949,G12950,G12951,G12952,G12953,G12954,G12955,G12956,G12957,G12958,G12959,G12960,
       G12961,G12962,G12963,G12964,G12965,G12966,G12967,G12968,G12969,G12970,G12971,G12972,G12973,G12974,G12975,G12976,G12977,G12978,G12979,G12980,
       G12981,G12982,G12983,G12984,G12985,G12986,G12987,G12988,G12989,G12990,G12991,G12992,G12993,G12994,G12995,G12996,G12997,G12998,G12999,G13000,
       G13001,G13002,G13003,G13004,G13005,G13006,G13007,G13008,G13009,G13010,G13011,G13012,G13013,G13014,G13015,G13016,G13017,G13018,G13019,G13020,
       G13021,G13022,G13023,G13024,G13025,G13026,G13027,G13028,G13029,G13030,G13031,G13032,G13033,G13034,G13035,G13036,G13037,G13038,G13039,G13040,
       G13041,G13042,G13043,G13044,G13045,G13046,G13047,G13048,G13049,G13050,G13051,G13052,G13053,G13054,G13055,G13056,G13057,G13058,G13059,G13060,
       G13061,G13062,G13063,G13064,G13065,G13066,G13067,G13068,G13069,G13070,G13071,G13072,G13073,G13074,G13075,G13076,G13077,G13078,G13079,G13080,
       G13081,G13082,G13083,G13084,G13085,G13086,G13087,G13088,G13089,G13090,G13091,G13092,G13093,G13094,G13095,G13096,G13097,G13098,G13099,G13100,
       G13101,G13102,G13103,G13104,G13105,G13106,G13107,G13108,G13109,G13110,G13111,G13112,G13113,G13114,G13115,G13116,G13117,G13118,G13119,G13120,
       G13121,G13122,G13123,G13124,G13125,G13126,G13127,G13128,G13129,G13130,G13131,G13132,G13133,G13134,G13135,G13136,G13137,G13138,G13139,G13140,
       G13141,G13142,G13143,G13144,G13145,G13146,G13147,G13148,G13149,G13150,G13151,G13152,G13153,G13154,G13155,G13156,G13157,G13158,G13159,G13160,
       G13161,G13162,G13163,G13164,G13165,G13166,G13167,G13168,G13169,G13170,G13171,G13172,G13173,G13174,G13175,G13176,G13177,G13178,G13179,G13180,
       G13181,G13182,G13183,G13184,G13185,G13186,G13187,G13188,G13189,G13190,G13191,G13192,G13193,G13194,G13195,G13196,G13197,G13198,G13199,G13200,
       G13201,G13202,G13203,G13204,G13205,G13206,G13207,G13208,G13209,G13210,G13211,G13212,G13213,G13214,G13215,G13216,G13217,G13218,G13219,G13220,
       G13221,G13222,G13223,G13224,G13225,G13226,G13227,G13228,G13229,G13230,G13231,G13232,G13233,G13234,G13235,G13236,G13237,G13238,G13239,G13240,
       G13241,G13242,G13243,G13244,G13245,G13246,G13247,G13248,G13249,G13250,G13251,G13252,G13253,G13254,G13255,G13256,G13257,G13258,G13259,G13260,
       G13261,G13262,G13263,G13264,G13265,G13266,G13267,G13268,G13269,G13270,G13271,G13272,G13273,G13274,G13275,G13276,G13277,G13278,G13279,G13280,
       G13281,G13282,G13283,G13284,G13285,G13286,G13287,G13288,G13289,G13290,G13291,G13292,G13293,G13294,G13295,G13296,G13297,G13298,G13299,G13300,
       G13301,G13302,G13303,G13304,G13305,G13306,G13307,G13308,G13309,G13310,G13311,G13312,G13313,G13314,G13315,G13316,G13317,G13318,G13319,G13320,
       G13321,G13322,G13323,G13324,G13325,G13326,G13327,G13328,G13329,G13330,G13331,G13332,G13333,G13334,G13335,G13336,G13337,G13338,G13339,G13340,
       G13341,G13342,G13343,G13344,G13345,G13346,G13347,G13348,G13349,G13350,G13351,G13352,G13353,G13354,G13355,G13356,G13357,G13358,G13359,G13360,
       G13361,G13362,G13363,G13364,G13365,G13366,G13367,G13368,G13369,G13370,G13371,G13372,G13373,G13374,G13375,G13376,G13377,G13378,G13379,G13380,
       G13381,G13382,G13383,G13384,G13385,G13386,G13387,G13388,G13389,G13390,G13391,G13392,G13393,G13394,G13395,G13396,G13397,G13398,G13399,G13400,
       G13401,G13402,G13403,G13404,G13405,G13406,G13407,G13408,G13409,G13410,G13411,G13412,G13413,G13414,G13415,G13416,G13417,G13418,G13419,G13420,
       G13421,G13422,G13423,G13424,G13425,G13426,G13427,G13428,G13429,G13430,G13431,G13432,G13433,G13434,G13435,G13436,G13437,G13438,G13439,G13440,
       G13441,G13442,G13443,G13444,G13445,G13446,G13447,G13448,G13449,G13450,G13451,G13452,G13453,G13454,G13455,G13456,G13457,G13458,G13459,G13460,
       G13461,G13462,G13463,G13464,G13465,G13466,G13467,G13468,G13469,G13470,G13471,G13472,G13473,G13474,G13475,G13476,G13477,G13478,G13479,G13480,
       G13481,G13482,G13483,G13484,G13485,G13486,G13487,G13488,G13489,G13490,G13491,G13492,G13493,G13494,G13495,G13496,G13497,G13498,G13499,G13500,
       G13501,G13502,G13503,G13504,G13505,G13506,G13507,G13508,G13509,G13510,G13511,G13512,G13513,G13514,G13515,G13516,G13517,G13518,G13519,G13520,
       G13521,G13522,G13523,G13524,G13525,G13526,G13527,G13528,G13529,G13530,G13531,G13532,G13533,G13534,G13535,G13536,G13537,G13538,G13539,G13540,
       G13541,G13542,G13543,G13544,G13545,G13546,G13547,G13548,G13549,G13550,G13551,G13552,G13553,G13554,G13555,G13556,G13557,G13558,G13559,G13560,
       G13561,G13562,G13563,G13564,G13565,G13566,G13567,G13568,G13569,G13570,G13571,G13572,G13573,G13574,G13575,G13576,G13577,G13578,G13579,G13580,
       G13581,G13582,G13583,G13584,G13585,G13586,G13587,G13588,G13589,G13590,G13591,G13592,G13593,G13594,G13595,G13596,G13597,G13598,G13599,G13600,
       G13601,G13602,G13603,G13604,G13605,G13606,G13607,G13608,G13609,G13610,G13611,G13612,G13613,G13614,G13615,G13616,G13617,G13618,G13619,G13620,
       G13621,G13622,G13623,G13624,G13625,G13626,G13627,G13628,G13629,G13630,G13631,G13632,G13633,G13634,G13635,G13636,G13637,G13638,G13639,G13640,
       G13641,G13642,G13643,G13644,G13645,G13646,G13647,G13648,G13649,G13650,G13651,G13652,G13653,G13654,G13655,G13656,G13657,G13658,G13659,G13660,
       G13661,G13662,G13663,G13664,G13665,G13666,G13667,G13668,G13669,G13670,G13671,G13672,G13673,G13674,G13675,G13676,G13677,G13678,G13679,G13680,
       G13681,G13682,G13683,G13684,G13685,G13686,G13687,G13688,G13689,G13690,G13691,G13692,G13693,G13694,G13695,G13696,G13697,G13698,G13699,G13700,
       G13701,G13702,G13703,G13704,G13705,G13706,G13707,G13708,G13709,G13710,G13711,G13712,G13713,G13714,G13715,G13716,G13717,G13718,G13719,G13720,
       G13721,G13722,G13723,G13724,G13725,G13726,G13727,G13728,G13729,G13730,G13731,G13732,G13733,G13734,G13735,G13736,G13737,G13738,G13739,G13740,
       G13741,G13742,G13743,G13744,G13745,G13746,G13747,G13748,G13749,G13750,G13751,G13752,G13753,G13754,G13755,G13756,G13757,G13758,G13759,G13760,
       G13761,G13762,G13763,G13764,G13765,G13766,G13767,G13768,G13769,G13770,G13771,G13772,G13773,G13774,G13775,G13776,G13777,G13778,G13779,G13780,
       G13781,G13782,G13783,G13784,G13785,G13786,G13787,G13788,G13789,G13790,G13791,G13792,G13793,G13794,G13795,G13796,G13797,G13798,G13799,G13800,
       G13801,G13802,G13803,G13804,G13805,G13806,G13807,G13808,G13809,G13810,G13811,G13812,G13813,G13814,G13815,G13816,G13817,G13818,G13819,G13820,
       G13821,G13822,G13823,G13824,G13825,G13826,G13827,G13828,G13829,G13830,G13831,G13832,G13833,G13834,G13835,G13836,G13837,G13838,G13839,G13840,
       G13841,G13842,G13843,G13844,G13845,G13846,G13847,G13848,G13849,G13850,G13851,G13852,G13853,G13854,G13855,G13856,G13857,G13858,G13859,G13860,
       G13861,G13862,G13863,G13864,G13865,G13866,G13867,G13868,G13869,G13870,G13871,G13872,G13873,G13874,G13875,G13876,G13877,G13878,G13879,G13880,
       G13881,G13882,G13883,G13884,G13885,G13886,G13887,G13888,G13889,G13890,G13891,G13892,G13893,G13894,G13895,G13896,G13897,G13898,G13899,G13900,
       G13901,G13902,G13903,G13904,G13905,G13906,G13907,G13908,G13909,G13910,G13911,G13912,G13913,G13914,G13915,G13916,G13917,G13918,G13919,G13920,
       G13921,G13922,G13923,G13924,G13925,G13926,G13927,G13928,G13929,G13930,G13931,G13932,G13933,G13934,G13935,G13936,G13937,G13938,G13939,G13940,
       G13941,G13942,G13943,G13944,G13945,G13946,G13947,G13948,G13949,G13950,G13951,G13952,G13953,G13954,G13955,G13956,G13957,G13958,G13959,G13960,
       G13961,G13962,G13963,G13964,G13965,G13966,G13967,G13968,G13969,G13970,G13971,G13972,G13973,G13974,G13975,G13976,G13977,G13978,G13979,G13980,
       G13981,G13982,G13983,G13984,G13985,G13986,G13987,G13988,G13989,G13990,G13991,G13992,G13993,G13994,G13995,G13996,G13997,G13998,G13999,G14000,
       G14001,G14002,G14003,G14004,G14005,G14006,G14007,G14008,G14009,G14010,G14011,G14012,G14013,G14014,G14015,G14016,G14017,G14018,G14019,G14020,
       G14021,G14022,G14023,G14024,G14025,G14026,G14027,G14028,G14029,G14030,G14031,G14032,G14033,G14034,G14035,G14036,G14037,G14038,G14039,G14040,
       G14041,G14042,G14043,G14044,G14045,G14046,G14047,G14048,G14049,G14050,G14051,G14052,G14053,G14054,G14055,G14056,G14057,G14058,G14059,G14060,
       G14061,G14062,G14063,G14064,G14065,G14066,G14067,G14068,G14069,G14070,G14071,G14072,G14073,G14074,G14075,G14076,G14077,G14078,G14079,G14080,
       G14081,G14082,G14083,G14084,G14085,G14086,G14087,G14088,G14089,G14090,G14091,G14092,G14093,G14094,G14095,G14096,G14097,G14098,G14099,G14100,
       G14101,G14102,G14103,G14104,G14105,G14106,G14107,G14108,G14109,G14110,G14111,G14112,G14113,G14114,G14115,G14116,G14117,G14118,G14119,G14120,
       G14121,G14122,G14123,G14124,G14125,G14126,G14127,G14128,G14129,G14130,G14131,G14132,G14133,G14134,G14135,G14136,G14137,G14138,G14139,G14140,
       G14141,G14142,G14143,G14144,G14145,G14146,G14147,G14148,G14149,G14150,G14151,G14152,G14153,G14154,G14155,G14156,G14157,G14158,G14159,G14160,
       G14161,G14162,G14163,G14164,G14165,G14166,G14167,G14168,G14169,G14170,G14171,G14172,G14173,G14174,G14175,G14176,G14177,G14178,G14179,G14180,
       G14181,G14182,G14183,G14184,G14185,G14186,G14187,G14188,G14189,G14190,G14191,G14192,G14193,G14194,G14195,G14196,G14197,G14198,G14199,G14200,
       G14201,G14202,G14203,G14204,G14205,G14206,G14207,G14208,G14209,G14210,G14211,G14212,G14213,G14214,G14215,G14216,G14217,G14218,G14219,G14220,
       G14221,G14222,G14223,G14224,G14225,G14226,G14227,G14228,G14229,G14230,G14231,G14232,G14233,G14234,G14235,G14236,G14237,G14238,G14239,G14240,
       G14241,G14242,G14243,G14244,G14245,G14246,G14247,G14248,G14249,G14250,G14251,G14252,G14253,G14254,G14255,G14256,G14257,G14258,G14259,G14260,
       G14261,G14262,G14263,G14264,G14265,G14266,G14267,G14268,G14269,G14270,G14271,G14272,G14273,G14274,G14275,G14276,G14277,G14278,G14279,G14280,
       G14281,G14282,G14283,G14284,G14285,G14286,G14287,G14288,G14289,G14290,G14291,G14292,G14293,G14294,G14295,G14296,G14297,G14298,G14299,G14300,
       G14301,G14302,G14303,G14304,G14305,G14306,G14307,G14308,G14309,G14310,G14311,G14312,G14313,G14314,G14315,G14316,G14317,G14318,G14319,G14320,
       G14321,G14322,G14323,G14324,G14325,G14326,G14327,G14328,G14329,G14330,G14331,G14332,G14333,G14334,G14335,G14336,G14337,G14338,G14339,G14340,
       G14341,G14342,G14343,G14344,G14345,G14346,G14347,G14348,G14349,G14350,G14351,G14352,G14353,G14354,G14355,G14356,G14357,G14358,G14359,G14360,
       G14361,G14362,G14363,G14364,G14365,G14366,G14367,G14368,G14369,G14370,G14371,G14372,G14373,G14374,G14375,G14376,G14377,G14378,G14379,G14380,
       G14381,G14382,G14383,G14384,G14385,G14386,G14387,G14388,G14389,G14390,G14391,G14392,G14393,G14394,G14395,G14396,G14397,G14398,G14399,G14400,
       G14401,G14402,G14403,G14404,G14405,G14406,G14407,G14408,G14409,G14410,G14411,G14412,G14413,G14414,G14415,G14416,G14417,G14418,G14419,G14420,
       G14421,G14422,G14423,G14424,G14425,G14426,G14427,G14428,G14429,G14430,G14431,G14432,G14433,G14434,G14435,G14436,G14437,G14438,G14439,G14440,
       G14441,G14442,G14443,G14444,G14445,G14446,G14447,G14448,G14449,G14450,G14451,G14452,G14453,G14454,G14455,G14456,G14457,G14458,G14459,G14460,
       G14461,G14462,G14463,G14464,G14465,G14466,G14467,G14468,G14469,G14470,G14471,G14472,G14473,G14474,G14475,G14476,G14477,G14478,G14479,G14480,
       G14481,G14482,G14483,G14484,G14485,G14486,G14487,G14488,G14489,G14490,G14491,G14492,G14493,G14494,G14495,G14496,G14497,G14498,G14499,G14500,
       G14501,G14502,G14503,G14504,G14505,G14506,G14507,G14508,G14509,G14510,G14511,G14512,G14513,G14514,G14515,G14516,G14517,G14518,G14519,G14520,
       G14521,G14522,G14523,G14524,G14525,G14526,G14527,G14528,G14529,G14530,G14531,G14532,G14533,G14534,G14535,G14536,G14537,G14538,G14539,G14540,
       G14541,G14542,G14543,G14544,G14545,G14546,G14547,G14548,G14549,G14550,G14551,G14552,G14553,G14554,G14555,G14556,G14557,G14558,G14559,G14560,
       G14561,G14562,G14563,G14564,G14565,G14566,G14567,G14568,G14569,G14570,G14571,G14572,G14573,G14574,G14575,G14576,G14577,G14578,G14579,G14580,
       G14581,G14582,G14583,G14584,G14585,G14586,G14587,G14588,G14589,G14590,G14591,G14592,G14593,G14594,G14595,G14596,G14597,G14598,G14599,G14600,
       G14601,G14602,G14603,G14604,G14605,G14606,G14607,G14608,G14609,G14610,G14611,G14612,G14613,G14614,G14615,G14616,G14617,G14618,G14619,G14620,
       G14621,G14622,G14623,G14624,G14625,G14626,G14627,G14628,G14629,G14630,G14631,G14632,G14633,G14634,G14635,G14636,G14637,G14638,G14639,G14640,
       G14641,G14642,G14643,G14644,G14645,G14646,G14647,G14648,G14649,G14650,G14651,G14652,G14653,G14654,G14655,G14656,G14657,G14658,G14659,G14660,
       G14661,G14662,G14663,G14664,G14665,G14666,G14667,G14668,G14669,G14670,G14671,G14672,G14673,G14674,G14675,G14676,G14677,G14678,G14679,G14680,
       G14681,G14682,G14683,G14684,G14685,G14686,G14687,G14688,G14689,G14690,G14691,G14692,G14693,G14694,G14695,G14696,G14697,G14698,G14699,G14700,
       G14701,G14702,G14703,G14704,G14705,G14706,G14707,G14708,G14709,G14710,G14711,G14712,G14713,G14714,G14715,G14716,G14717,G14718,G14719,G14720,
       G14721,G14722,G14723,G14724,G14725,G14726,G14727,G14728,G14729,G14730,G14731,G14732,G14733,G14734,G14735,G14736,G14737,G14738,G14739,G14740,
       G14741,G14742,G14743,G14744,G14745,G14746,G14747,G14748,G14749,G14750,G14751,G14752,G14753,G14754,G14755,G14756,G14757,G14758,G14759,G14760,
       G14761,G14762,G14763,G14764,G14765,G14766,G14767,G14768,G14769,G14770,G14771,G14772,G14773,G14774,G14775,G14776,G14777,G14778,G14779,G14780,
       G14781,G14782,G14783,G14784,G14785,G14786,G14787,G14788,G14789,G14790,G14791,G14792,G14793,G14794,G14795,G14796,G14797,G14798,G14799,G14800,
       G14801,G14802,G14803,G14804,G14805,G14806,G14807,G14808,G14809,G14810,G14811,G14812,G14813,G14814,G14815,G14816,G14817,G14818,G14819,G14820,
       G14821,G14822,G14823,G14824,G14825,G14826,G14827,G14828,G14829,G14830,G14831,G14832,G14833,G14834,G14835,G14836,G14837,G14838,G14839,G14840,
       G14841,G14842,G14843,G14844,G14845,G14846,G14847,G14848,G14849,G14850,G14851,G14852,G14853,G14854,G14855,G14856,G14857,G14858,G14859,G14860,
       G14861,G14862,G14863,G14864,G14865,G14866,G14867,G14868,G14869,G14870,G14871,G14872,G14873,G14874,G14875,G14876,G14877,G14878,G14879,G14880,
       G14881,G14882,G14883,G14884,G14885,G14886,G14887,G14888,G14889,G14890,G14891,G14892,G14893,G14894,G14895,G14896,G14897,G14898,G14899,G14900,
       G14901,G14902,G14903,G14904,G14905,G14906,G14907,G14908,G14909,G14910,G14911,G14912,G14913,G14914,G14915,G14916,G14917,G14918,G14919,G14920,
       G14921,G14922,G14923,G14924,G14925,G14926,G14927,G14928,G14929,G14930,G14931,G14932,G14933,G14934,G14935,G14936,G14937,G14938,G14939,G14940,
       G14941,G14942,G14943,G14944,G14945,G14946,G14947,G14948,G14949,G14950,G14951,G14952,G14953,G14954,G14955,G14956,G14957,G14958,G14959,G14960,
       G14961,G14962,G14963,G14964,G14965,G14966,G14967,G14968,G14969,G14970,G14971,G14972,G14973,G14974,G14975,G14976,G14977,G14978,G14979,G14980,
       G14981,G14982,G14983,G14984,G14985,G14986,G14987,G14988,G14989,G14990,G14991,G14992,G14993,G14994,G14995,G14996,G14997,G14998,G14999,G15000,
       G15001,G15002,G15003,G15004,G15005,G15006,G15007,G15008,G15009,G15010,G15011,G15012,G15013,G15014,G15015,G15016,G15017,G15018,G15019,G15020,
       G15021,G15022,G15023,G15024,G15025,G15026,G15027,G15028,G15029,G15030,G15031,G15032,G15033,G15034,G15035,G15036,G15037,G15038,G15039,G15040,
       G15041,G15042,G15043,G15044,G15045,G15046,G15047,G15048,G15049,G15050,G15051,G15052,G15053,G15054,G15055,G15056,G15057,G15058,G15059,G15060,
       G15061,G15062,G15063,G15064,G15065,G15066,G15067,G15068,G15069,G15070,G15071,G15072,G15073,G15074,G15075,G15076,G15077,G15078,G15079,G15080,
       G15081,G15082,G15083,G15084,G15085,G15086,G15087,G15088,G15089,G15090,G15091,G15092,G15093,G15094,G15095,G15096,G15097,G15098,G15099,G15100,
       G15101,G15102,G15103,G15104,G15105,G15106,G15107,G15108,G15109,G15110,G15111,G15112,G15113,G15114,G15115,G15116,G15117,G15118,G15119,G15120,
       G15121,G15122,G15123,G15124,G15125,G15126,G15127,G15128,G15129,G15130,G15131,G15132,G15133,G15134,G15135,G15136,G15137,G15138,G15139,G15140,
       G15141,G15142,G15143,G15144,G15145,G15146,G15147,G15148,G15149,G15150,G15151,G15152,G15153,G15154,G15155,G15156,G15157,G15158,G15159,G15160,
       G15161,G15162,G15163,G15164,G15165,G15166,G15167,G15168,G15169,G15170,G15171,G15172,G15173,G15174,G15175,G15176,G15177,G15178,G15179,G15180,
       G15181,G15182,G15183,G15184,G15185,G15186,G15187,G15188,G15189,G15190,G15191,G15192,G15193,G15194,G15195,G15196,G15197,G15198,G15199,G15200,
       G15201,G15202,G15203,G15204,G15205,G15206,G15207,G15208,G15209,G15210,G15211,G15212,G15213,G15214,G15215,G15216,G15217,G15218,G15219,G15220,
       G15221,G15222,G15223,G15224,G15225,G15226,G15227,G15228,G15229,G15230,G15231,G15232,G15233,G15234,G15235,G15236,G15237,G15238,G15239,G15240,
       G15241,G15242,G15243,G15244,G15245,G15246,G15247,G15248,G15249,G15250,G15251,G15252,G15253,G15254,G15255,G15256,G15257,G15258,G15259,G15260,
       G15261,G15262,G15263,G15264,G15265,G15266,G15267,G15268,G15269,G15270,G15271,G15272,G15273,G15274,G15275,G15276,G15277,G15278,G15279,G15280,
       G15281,G15282,G15283,G15284,G15285,G15286,G15287,G15288,G15289,G15290,G15291,G15292,G15293,G15294,G15295,G15296,G15297,G15298,G15299,G15300,
       G15301,G15302,G15303,G15304,G15305,G15306,G15307,G15308,G15309,G15310,G15311,G15312,G15313,G15314,G15315,G15316,G15317,G15318,G15319,G15320,
       G15321,G15322,G15323,G15324,G15325,G15326,G15327,G15328,G15329,G15330,G15331,G15332,G15333,G15334,G15335,G15336,G15337,G15338,G15339,G15340,
       G15341,G15342,G15343,G15344,G15345,G15346,G15347,G15348,G15349,G15350,G15351,G15352,G15353,G15354,G15355,G15356,G15357,G15358,G15359,G15360,
       G15361,G15362,G15363,G15364,G15365,G15366,G15367,G15368,G15369,G15370,G15371,G15372,G15373,G15374,G15375,G15376,G15377,G15378,G15379,G15380,
       G15381,G15382,G15383,G15384,G15385,G15386,G15387,G15388,G15389,G15390,G15391,G15392,G15393,G15394,G15395,G15396,G15397,G15398,G15399,G15400,
       G15401,G15402,G15403,G15404,G15405,G15406,G15407,G15408,G15409,G15410,G15411,G15412,G15413,G15414,G15415,G15416,G15417,G15418,G15419,G15420,
       G15421,G15422,G15423,G15424,G15425,G15426,G15427,G15428,G15429,G15430,G15431,G15432,G15433,G15434,G15435,G15436,G15437,G15438,G15439,G15440,
       G15441,G15442,G15443,G15444,G15445,G15446,G15447,G15448,G15449,G15450,G15451,G15452,G15453,G15454,G15455,G15456,G15457,G15458,G15459,G15460,
       G15461,G15462,G15463,G15464,G15465,G15466,G15467,G15468,G15469,G15470,G15471,G15472,G15473,G15474,G15475,G15476,G15477,G15478,G15479,G15480,
       G15481,G15482,G15483,G15484,G15485,G15486,G15487,G15488,G15489,G15490,G15491,G15492,G15493,G15494,G15495,G15496,G15497,G15498,G15499,G15500,
       G15501,G15502,G15503,G15504,G15505,G15506,G15507,G15508,G15509,G15510,G15511,G15512,G15513,G15514,G15515,G15516,G15517,G15518,G15519,G15520,
       G15521,G15522,G15523,G15524,G15525,G15526,G15527,G15528,G15529,G15530,G15531,G15532,G15533,G15534,G15535,G15536,G15537,G15538,G15539,G15540,
       G15541,G15542,G15543,G15544,G15545,G15546,G15547,G15548,G15549,G15550,G15551,G15552,G15553,G15554,G15555,G15556,G15557,G15558,G15559,G15560,
       G15561,G15562,G15563,G15564,G15565,G15566,G15567,G15568,G15569,G15570,G15571,G15572,G15573,G15574,G15575,G15576,G15577,G15578,G15579,G15580,
       G15581,G15582,G15583,G15584,G15585,G15586,G15587,G15588,G15589,G15590,G15591,G15592,G15593,G15594,G15595,G15596,G15597,G15598,G15599,G15600,
       G15601,G15602,G15603,G15604,G15605,G15606,G15607,G15608,G15609,G15610,G15611,G15612,G15613,G15614,G15615,G15616,G15617,G15618,G15619,G15620,
       G15621,G15622,G15623,G15624,G15625,G15626,G15627,G15628,G15629,G15630,G15631,G15632,G15633,G15634,G15635,G15636,G15637,G15638,G15639,G15640,
       G15641,G15642,G15643,G15644,G15645,G15646,G15647,G15648,G15649,G15650,G15651,G15652,G15653,G15654,G15655,G15656,G15657,G15658,G15659,G15660,
       G15661,G15662,G15663,G15664,G15665,G15666,G15667,G15668,G15669,G15670,G15671,G15672,G15673,G15674,G15675,G15676,G15677,G15678,G15679,G15680,
       G15681,G15682,G15683,G15684,G15685,G15686,G15687,G15688,G15689,G15690,G15691,G15692,G15693,G15694,G15695,G15696,G15697,G15698,G15699,G15700,
       G15701,G15702,G15703,G15704,G15705,G15706,G15707,G15708,G15709,G15710,G15711,G15712,G15713,G15714,G15715,G15716,G15717,G15718,G15719,G15720,
       G15721,G15722,G15723,G15724,G15725,G15726,G15727,G15728,G15729,G15730,G15731,G15732,G15733,G15734,G15735,G15736,G15737,G15738,G15739,G15740,
       G15741,G15742,G15743,G15744,G15745,G15746,G15747,G15748,G15749,G15750,G15751,G15752,G15753,G15754,G15755,G15756,G15757,G15758,G15759,G15760,
       G15761,G15762,G15763,G15764,G15765,G15766,G15767,G15768,G15769,G15770,G15771,G15772,G15773,G15774,G15775,G15776,G15777,G15778,G15779,G15780,
       G15781,G15782,G15783,G15784,G15785,G15786,G15787,G15788,G15789,G15790,G15791,G15792,G15793,G15794,G15795,G15796,G15797,G15798,G15799,G15800,
       G15801,G15802,G15803,G15804,G15805,G15806,G15807,G15808,G15809,G15810,G15811,G15812,G15813,G15814,G15815,G15816,G15817,G15818,G15819,G15820,
       G15821,G15822,G15823,G15824,G15825,G15826,G15827,G15828,G15829,G15830,G15831,G15832,G15833,G15834,G15835,G15836,G15837,G15838,G15839,G15840,
       G15841,G15842,G15843,G15844,G15845,G15846,G15847,G15848,G15849,G15850,G15851,G15852,G15853,G15854,G15855,G15856,G15857,G15858,G15859,G15860,
       G15861,G15862,G15863,G15864,G15865,G15866,G15867,G15868,G15869,G15870,G15871,G15872,G15873,G15874,G15875,G15876,G15877,G15878,G15879,G15880,
       G15881,G15882,G15883,G15884,G15885,G15886,G15887,G15888,G15889,G15890,G15891,G15892,G15893,G15894,G15895,G15896,G15897,G15898,G15899,G15900,
       G15901,G15902,G15903,G15904,G15905,G15906,G15907,G15908,G15909,G15910,G15911,G15912,G15913,G15914,G15915,G15916,G15917,G15918,G15919,G15920,
       G15921,G15922,G15923,G15924,G15925,G15926,G15927,G15928,G15929,G15930,G15931,G15932,G15933,G15934,G15935,G15936,G15937,G15938,G15939,G15940,
       G15941,G15942,G15943,G15944,G15945,G15946,G15947,G15948,G15949,G15950,G15951,G15952,G15953,G15954,G15955,G15956,G15957,G15958,G15959,G15960,
       G15961,G15962,G15963,G15964,G15965,G15966,G15967,G15968,G15969,G15970,G15971,G15972,G15973,G15974,G15975,G15976,G15977,G15978,G15979,G15980,
       G15981,G15982,G15983,G15984,G15985,G15986,G15987,G15988,G15989,G15990,G15991,G15992,G15993,G15994,G15995,G15996,G15997,G15998,G15999,G16000,
       G16001,G16002,G16003,G16004,G16005,G16006,G16007,G16008,G16009,G16010,G16011,G16012,G16013,G16014,G16015,G16016,G16017,G16018,G16019,G16020,
       G16021,G16022,G16023,G16024,G16025,G16026,G16027,G16028,G16029,G16030,G16031,G16032,G16033,G16034,G16035,G16036,G16037,G16038,G16039,G16040,
       G16041,G16042,G16043,G16044,G16045,G16046,G16047,G16048,G16049,G16050,G16051,G16052,G16053,G16054,G16055,G16056,G16057,G16058,G16059,G16060,
       G16061,G16062,G16063,G16064,G16065,G16066,G16067,G16068,G16069,G16070,G16071,G16072,G16073,G16074,G16075,G16076,G16077,G16078,G16079,G16080,
       G16081,G16082,G16083,G16084,G16085,G16086,G16087,G16088,G16089,G16090,G16091,G16092,G16093,G16094,G16095,G16096,G16097,G16098,G16099,G16100,
       G16101,G16102,G16103,G16104,G16105,G16106,G16107,G16108,G16109,G16110,G16111,G16112,G16113,G16114,G16115,G16116,G16117,G16118,G16119,G16120,
       G16121,G16122,G16123,G16124,G16125,G16126,G16127,G16128,G16129,G16130,G16131,G16132,G16133,G16134,G16135,G16136,G16137,G16138,G16139,G16140,
       G16141,G16142,G16143,G16144,G16145,G16146,G16147,G16148,G16149,G16150,G16151,G16152,G16153,G16154,G16155,G16156,G16157,G16158,G16159,G16160,
       G16161,G16162,G16163,G16164,G16165,G16166,G16167,G16168,G16169,G16170,G16171,G16172,G16173,G16174,G16175,G16176,G16177,G16178,G16179,G16180,
       G16181,G16182,G16183,G16184,G16185,G16186,G16187,G16188,G16189,G16190,G16191,G16192,G16193,G16194,G16195,G16196,G16197,G16198,G16199,G16200,
       G16201,G16202,G16203,G16204,G16205,G16206,G16207,G16208,G16209,G16210,G16211,G16212,G16213,G16214,G16215,G16216,G16217,G16218,G16219,G16220,
       G16221,G16222,G16223,G16224,G16225,G16226,G16227,G16228,G16229,G16230,G16231,G16232,G16233,G16234,G16235,G16236,G16237,G16238,G16239,G16240,
       G16241,G16242,G16243,G16244,G16245,G16246,G16247,G16248,G16249,G16250,G16251,G16252,G16253,G16254,G16255,G16256,G16257,G16258,G16259,G16260,
       G16261,G16262,G16263,G16264,G16265,G16266,G16267,G16268,G16269,G16270,G16271,G16272,G16273,G16274,G16275,G16276,G16277,G16278,G16279,G16280,
       G16281,G16282,G16283,G16284,G16285,G16286,G16287,G16288,G16289,G16290,G16291,G16292,G16293,G16294,G16295,G16296,G16297,G16298,G16299,G16300,
       G16301,G16302,G16303,G16304,G16305,G16306,G16307,G16308,G16309,G16310,G16311,G16312,G16313,G16314,G16315,G16316,G16317,G16318,G16319,G16320,
       G16321,G16322,G16323,G16324,G16325,G16326,G16327,G16328,G16329,G16330,G16331,G16332,G16333,G16334,G16335,G16336,G16337,G16338,G16339,G16340,
       G16341,G16342,G16343,G16344,G16345,G16346,G16347,G16348,G16349,G16350,G16351,G16352,G16353,G16354,G16355,G16356,G16357,G16358,G16359,G16360,
       G16361,G16362,G16363,G16364,G16365,G16366,G16367,G16368,G16369,G16370,G16371,G16372,G16373,G16374,G16375,G16376,G16377,G16378,G16379,G16380,
       G16381,G16382,G16383,G16384,G16385,G16386,G16387,G16388,G16389,G16390,G16391,G16392,G16393,G16394,G16395,G16396,G16397,G16398,G16399,G16400,
       G16401,G16402,G16403,G16404,G16405,G16406,G16407,G16408,G16409,G16410,G16411,G16412,G16413,G16414,G16415,G16416,G16417,G16418,G16419,G16420,
       G16421,G16422,G16423,G16424,G16425,G16426,G16427,G16428,G16429,G16430,G16431,G16432,G16433,G16434,G16435,G16436,G16437,G16438,G16439,G16440,
       G16441,G16442,G16443,G16444,G16445,G16446,G16447,G16448,G16449,G16450,G16451,G16452,G16453,G16454,G16455,G16456,G16457,G16458,G16459,G16460,
       G16461,G16462,G16463,G16464,G16465,G16466,G16467,G16468,G16469,G16470,G16471,G16472,G16473,G16474,G16475,G16476,G16477,G16478,G16479,G16480,
       G16481,G16482,G16483,G16484,G16485,G16486,G16487,G16488,G16489,G16490,G16491,G16492,G16493,G16494,G16495,G16496,G16497,G16498,G16499,G16500,
       G16501,G16502,G16503,G16504,G16505,G16506,G16507,G16508,G16509,G16510,G16511,G16512,G16513,G16514,G16515,G16516,G16517,G16518,G16519,G16520,
       G16521,G16522,G16523,G16524,G16525,G16526,G16527,G16528,G16529,G16530,G16531,G16532,G16533,G16534,G16535,G16536,G16537,G16538,G16539,G16540,
       G16541,G16542,G16543,G16544,G16545,G16546,G16547,G16548,G16549,G16550,G16551,G16552,G16553,G16554,G16555,G16556,G16557,G16558,G16559,G16560,
       G16561,G16562,G16563,G16564,G16565,G16566,G16567,G16568,G16569,G16570,G16571,G16572,G16573,G16574,G16575,G16576,G16577,G16578,G16579,G16580,
       G16581,G16582,G16583,G16584,G16585,G16586,G16587,G16588,G16589,G16590,G16591,G16592,G16593,G16594,G16595,G16596,G16597,G16598,G16599,G16600,
       G16601,G16602,G16603,G16604,G16605,G16606,G16607,G16608,G16609,G16610,G16611,G16612,G16613,G16614,G16615,G16616,G16617,G16618,G16619,G16620,
       G16621,G16622,G16623,G16624,G16625,G16626,G16627,G16628,G16629,G16630,G16631,G16632,G16633,G16634,G16635,G16636,G16637,G16638,G16639,G16640,
       G16641,G16642,G16643,G16644,G16645,G16646,G16647,G16648,G16649,G16650,G16651,G16652,G16653,G16654,G16655,G16656,G16657,G16658,G16659,G16660,
       G16661,G16662,G16663,G16664,G16665,G16666,G16667,G16668,G16669,G16670,G16671,G16672,G16673,G16674,G16675,G16676,G16677,G16678,G16679,G16680,
       G16681,G16682,G16683,G16684,G16685,G16686,G16687,G16688,G16689,G16690,G16691,G16692,G16693,G16694,G16695,G16696,G16697,G16698,G16699,G16700,
       G16701,G16702,G16703,G16704,G16705,G16706,G16707,G16708,G16709,G16710,G16711,G16712,G16713,G16714,G16715,G16716,G16717,G16718,G16719,G16720,
       G16721,G16722,G16723,G16724,G16725,G16726,G16727,G16728,G16729,G16730,G16731,G16732,G16733,G16734,G16735,G16736,G16737,G16738,G16739,G16740,
       G16741,G16742,G16743,G16744,G16745,G16746,G16747,G16748,G16749,G16750,G16751,G16752,G16753,G16754,G16755,G16756,G16757,G16758,G16759,G16760,
       G16761,G16762,G16763,G16764,G16765,G16766,G16767,G16768,G16769,G16770,G16771,G16772,G16773,G16774,G16775,G16776,G16777,G16778,G16779,G16780,
       G16781,G16782,G16783,G16784,G16785,G16786,G16787,G16788,G16789,G16790,G16791,G16792,G16793,G16794,G16795,G16796,G16797,G16798,G16799,G16800,
       G16801,G16802,G16803,G16804,G16805,G16806,G16807,G16808,G16809,G16810,G16811,G16812,G16813,G16814,G16815,G16816,G16817,G16818,G16819,G16820,
       G16821,G16822,G16823,G16824,G16825,G16826,G16827,G16828,G16829,G16830,G16831,G16832,G16833,G16834,G16835,G16836,G16837,G16838,G16839,G16840,
       G16841,G16842,G16843,G16844,G16845,G16846,G16847,G16848,G16849,G16850,G16851,G16852,G16853,G16854,G16855,G16856,G16857,G16858,G16859,G16860,
       G16861,G16862,G16863,G16864,G16865,G16866,G16867,G16868,G16869,G16870,G16871,G16872,G16873,G16874,G16875,G16876,G16877,G16878,G16879,G16880,
       G16881,G16882,G16883,G16884,G16885,G16886,G16887,G16888,G16889,G16890,G16891,G16892,G16893,G16894,G16895,G16896,G16897,G16898,G16899,G16900,
       G16901,G16902,G16903,G16904,G16905,G16906,G16907,G16908,G16909,G16910,G16911,G16912,G16913,G16914,G16915,G16916,G16917,G16918,G16919,G16920,
       G16921,G16922,G16923,G16924,G16925,G16926,G16927,G16928,G16929,G16930,G16931,G16932,G16933,G16934,G16935,G16936,G16937,G16938,G16939,G16940,
       G16941,G16942,G16943,G16944,G16945,G16946,G16947,G16948,G16949,G16950,G16951,G16952,G16953,G16954,G16955,G16956,G16957,G16958,G16959,G16960,
       G16961,G16962,G16963,G16964,G16965,G16966,G16967,G16968,G16969,G16970,G16971,G16972,G16973,G16974,G16975,G16976,G16977,G16978,G16979,G16980,
       G16981,G16982,G16983,G16984,G16985,G16986,G16987,G16988,G16989,G16990,G16991,G16992,G16993,G16994,G16995,G16996,G16997,G16998,G16999,G17000,
       G17001,G17002,G17003,G17004,G17005,G17006,G17007,G17008,G17009,G17010,G17011,G17012,G17013,G17014,G17015,G17016,G17017,G17018,G17019,G17020,
       G17021,G17022,G17023,G17024,G17025,G17026,G17027,G17028,G17029,G17030,G17031,G17032,G17033,G17034,G17035,G17036,G17037,G17038,G17039,G17040,
       G17041,G17042,G17043,G17044,G17045,G17046,G17047,G17048,G17049,G17050,G17051,G17052,G17053,G17054,G17055,G17056,G17057,G17058,G17059,G17060,
       G17061,G17062,G17063,G17064,G17065,G17066,G17067,G17068,G17069,G17070,G17071,G17072,G17073,G17074,G17075,G17076,G17077,G17078,G17079,G17080,
       G17081,G17082,G17083,G17084,G17085,G17086,G17087,G17088,G17089,G17090,G17091,G17092,G17093,G17094,G17095,G17096,G17097,G17098,G17099,G17100,
       G17101,G17102,G17103,G17104,G17105,G17106,G17107,G17108,G17109,G17110,G17111,G17112,G17113,G17114,G17115,G17116,G17117,G17118,G17119,G17120,
       G17121,G17122,G17123,G17124,G17125,G17126,G17127,G17128,G17129,G17130,G17131,G17132,G17133,G17134,G17135,G17136,G17137,G17138,G17139,G17140,
       G17141,G17142,G17143,G17144,G17145,G17146,G17147,G17148,G17149,G17150,G17151,G17152,G17153,G17154,G17155,G17156,G17157,G17158,G17159,G17160,
       G17161,G17162,G17163,G17164,G17165,G17166,G17167,G17168,G17169,G17170,G17171,G17172,G17173,G17174,G17175,G17176,G17177,G17178,G17179,G17180,
       G17181,G17182,G17183,G17184,G17185,G17186,G17187,G17188,G17189,G17190,G17191,G17192,G17193,G17194,G17195,G17196,G17197,G17198,G17199,G17200,
       G17201,G17202,G17203,G17204,G17205,G17206,G17207,G17208,G17209,G17210,G17211,G17212,G17213,G17214,G17215,G17216,G17217,G17218,G17219,G17220,
       G17221,G17222,G17223,G17224,G17225,G17226,G17227,G17228,G17229,G17230,G17231,G17232,G17233,G17234,G17235,G17236,G17237,G17238,G17239,G17240,
       G17241,G17242,G17243,G17244,G17245,G17246,G17247,G17248,G17249,G17250,G17251,G17252,G17253,G17254,G17255,G17256,G17257,G17258,G17259,G17260,
       G17261,G17262,G17263,G17264,G17265,G17266,G17267,G17268,G17269,G17270,G17271,G17272,G17273,G17274,G17275,G17276,G17277,G17278,G17279,G17280,
       G17281,G17282,G17283,G17284,G17285,G17286,G17287,G17288,G17289,G17290,G17291,G17292,G17293,G17294,G17295,G17296,G17297,G17298,G17299,G17300,
       G17301,G17302,G17303,G17304,G17305,G17306,G17307,G17308,G17309,G17310,G17311,G17312,G17313,G17314,G17315,G17316,G17317,G17318,G17319,G17320,
       G17321,G17322,G17323,G17324,G17325,G17326,G17327,G17328,G17329,G17330,G17331,G17332,G17333,G17334,G17335,G17336,G17337,G17338,G17339,G17340,
       G17341,G17342,G17343,G17344,G17345,G17346,G17347,G17348,G17349,G17350,G17351,G17352,G17353,G17354,G17355,G17356,G17357,G17358,G17359,G17360,
       G17361,G17362,G17363,G17364,G17365,G17366,G17367,G17368,G17369,G17370,G17371,G17372,G17373,G17374,G17375,G17376,G17377,G17378,G17379,G17380,
       G17381,G17382,G17383,G17384,G17385,G17386,G17387,G17388,G17389,G17390,G17391,G17392,G17393,G17394,G17395,G17396,G17397,G17398,G17399,G17400,
       G17401,G17402,G17403,G17404,G17405,G17406,G17407,G17408,G17409,G17410,G17411,G17412,G17413,G17414,G17415,G17416,G17417,G17418,G17419,G17420,
       G17421,G17422,G17423,G17424,G17425,G17426,G17427,G17428,G17429,G17430,G17431,G17432,G17433,G17434,G17435,G17436,G17437,G17438,G17439,G17440,
       G17441,G17442,G17443,G17444,G17445,G17446,G17447,G17448,G17449,G17450,G17451,G17452,G17453,G17454,G17455,G17456,G17457,G17458,G17459,G17460,
       G17461,G17462,G17463,G17464,G17465,G17466,G17467,G17468,G17469,G17470,G17471,G17472,G17473,G17474,G17475,G17476,G17477,G17478,G17479,G17480,
       G17481,G17482,G17483,G17484,G17485,G17486,G17487,G17488,G17489,G17490,G17491,G17492,G17493,G17494,G17495,G17496,G17497,G17498,G17499,G17500,
       G17501,G17502,G17503,G17504,G17505,G17506,G17507,G17508,G17509,G17510,G17511,G17512,G17513,G17514,G17515,G17516,G17517,G17518,G17519,G17520,
       G17521,G17522,G17523,G17524,G17525,G17526,G17527,G17528,G17529,G17530,G17531,G17532,G17533,G17534,G17535,G17536,G17537,G17538,G17539,G17540,
       G17541,G17542,G17543,G17544,G17545,G17546,G17547,G17548,G17549,G17550,G17551,G17552,G17553,G17554,G17555,G17556,G17557,G17558,G17559,G17560,
       G17561,G17562,G17563,G17564,G17565,G17566,G17567,G17568,G17569,G17570,G17571,G17572,G17573,G17574,G17575,G17576,G17577,G17578,G17579,G17580,
       G17581,G17582,G17583,G17584,G17585,G17586,G17587,G17588,G17589,G17590,G17591,G17592,G17593,G17594,G17595,G17596,G17597,G17598,G17599,G17600,
       G17601,G17602,G17603,G17604,G17605,G17606,G17607,G17608,G17609,G17610,G17611,G17612,G17613,G17614,G17615,G17616,G17617,G17618,G17619,G17620,
       G17621,G17622,G17623,G17624,G17625,G17626,G17627,G17628,G17629,G17630,G17631,G17632,G17633,G17634,G17635,G17636,G17637,G17638,G17639,G17640,
       G17641,G17642,G17643,G17644,G17645,G17646,G17647,G17648,G17649,G17650,G17651,G17652,G17653,G17654,G17655,G17656,G17657,G17658,G17659,G17660,
       G17661,G17662,G17663,G17664,G17665,G17666,G17667,G17668,G17669,G17670,G17671,G17672,G17673,G17674,G17675,G17676,G17677,G17678,G17679,G17680,
       G17681,G17682,G17683,G17684,G17685,G17686,G17687,G17688,G17689,G17690,G17691,G17692,G17693,G17694,G17695,G17696,G17697,G17698,G17699,G17700,
       G17701,G17702,G17703,G17704,G17705,G17706,G17707,G17708,G17709,G17710,G17711,G17712,G17713,G17714,G17715,G17716,G17717,G17718,G17719,G17720,
       G17721,G17722,G17723,G17724,G17725,G17726,G17727,G17728,G17729,G17730,G17731,G17732,G17733,G17734,G17735,G17736,G17737,G17738,G17739,G17740,
       G17741,G17742,G17743,G17744,G17745,G17746,G17747,G17748,G17749,G17750,G17751,G17752,G17753,G17754,G17755,G17756,G17757,G17758,G17759,G17760,
       G17761,G17762,G17763,G17764,G17765,G17766,G17767,G17768,G17769,G17770,G17771,G17772,G17773,G17774,G17775,G17776,G17777,G17778,G17779,G17780,
       G17781,G17782,G17783,G17784,G17785,G17786,G17787,G17788,G17789,G17790,G17791,G17792,G17793,G17794,G17795,G17796,G17797,G17798,G17799,G17800,
       G17801,G17802,G17803,G17804,G17805,G17806,G17807,G17808,G17809,G17810,G17811,G17812,G17813,G17814,G17815,G17816,G17817,G17818,G17819,G17820,
       G17821,G17822,G17823,G17824,G17825,G17826,G17827,G17828,G17829,G17830,G17831,G17832,G17833,G17834,G17835,G17836,G17837,G17838,G17839,G17840,
       G17841,G17842,G17843,G17844,G17845,G17846,G17847,G17848,G17849,G17850,G17851,G17852,G17853,G17854,G17855,G17856,G17857,G17858,G17859,G17860,
       G17861,G17862,G17863,G17864,G17865,G17866,G17867,G17868,G17869,G17870,G17871,G17872,G17873,G17874,G17875,G17876,G17877,G17878,G17879,G17880,
       G17881,G17882,G17883,G17884,G17885,G17886,G17887,G17888,G17889,G17890,G17891,G17892,G17893,G17894,G17895,G17896,G17897,G17898,G17899,G17900,
       G17901,G17902,G17903,G17904,G17905,G17906,G17907,G17908,G17909,G17910,G17911,G17912,G17913,G17914,G17915,G17916,G17917,G17918,G17919,G17920,
       G17921,G17922,G17923,G17924,G17925,G17926,G17927,G17928,G17929,G17930,G17931,G17932,G17933,G17934,G17935,G17936,G17937,G17938,G17939,G17940,
       G17941,G17942,G17943,G17944,G17945,G17946,G17947,G17948,G17949,G17950,G17951,G17952,G17953,G17954,G17955,G17956,G17957,G17958,G17959,G17960,
       G17961,G17962,G17963,G17964,G17965,G17966,G17967,G17968,G17969,G17970,G17971,G17972,G17973,G17974,G17975,G17976,G17977,G17978,G17979,G17980,
       G17981,G17982,G17983,G17984,G17985,G17986,G17987,G17988,G17989,G17990,G17991,G17992,G17993,G17994,G17995,G17996,G17997,G17998,G17999,G18000,
       G18001,G18002,G18003,G18004,G18005,G18006,G18007,G18008,G18009,G18010,G18011,G18012,G18013,G18014,G18015,G18016,G18017,G18018,G18019,G18020,
       G18021,G18022,G18023,G18024,G18025,G18026,G18027,G18028,G18029,G18030,G18031,G18032,G18033,G18034,G18035,G18036,G18037,G18038,G18039,G18040,
       G18041,G18042,G18043,G18044,G18045,G18046,G18047,G18048,G18049,G18050,G18051,G18052,G18053,G18054,G18055,G18056,G18057,G18058,G18059,G18060,
       G18061,G18062,G18063,G18064,G18065,G18066,G18067,G18068,G18069,G18070,G18071,G18072,G18073,G18074,G18075,G18076,G18077,G18078,G18079,G18080,
       G18081,G18082,G18083,G18084,G18085,G18086,G18087,G18088,G18089,G18090,G18091,G18092,G18093,G18094,G18095,G18096,G18097,G18098,G18099,G18100,
       G18101,G18102,G18103,G18104,G18105,G18106,G18107,G18108,G18109,G18110,G18111,G18112,G18113,G18114,G18115,G18116,G18117,G18118,G18119,G18120,
       G18121,G18122,G18123,G18124,G18125,G18126,G18127,G18128,G18129,G18130,G18131,G18132,G18133,G18134,G18135,G18136,G18137,G18138,G18139,G18140,
       G18141,G18142,G18143,G18144,G18145,G18146,G18147,G18148,G18149,G18150,G18151,G18152,G18153,G18154,G18155,G18156,G18157,G18158,G18159,G18160,
       G18161,G18162,G18163,G18164,G18165,G18166,G18167,G18168,G18169,G18170,G18171,G18172,G18173,G18174,G18175,G18176,G18177,G18178,G18179,G18180,
       G18181,G18182,G18183,G18184,G18185,G18186,G18187,G18188,G18189,G18190,G18191,G18192,G18193,G18194,G18195,G18196,G18197,G18198,G18199,G18200,
       G18201,G18202,G18203,G18204,G18205,G18206,G18207,G18208,G18209,G18210,G18211,G18212,G18213,G18214,G18215,G18216,G18217,G18218,G18219,G18220,
       G18221,G18222,G18223,G18224,G18225,G18226,G18227,G18228,G18229,G18230,G18231,G18232,G18233,G18234,G18235,G18236,G18237,G18238,G18239,G18240,
       G18241,G18242,G18243,G18244,G18245,G18246,G18247,G18248,G18249,G18250,G18251,G18252,G18253,G18254,G18255,G18256,G18257,G18258,G18259,G18260,
       G18261,G18262,G18263,G18264,G18265,G18266,G18267,G18268,G18269,G18270,G18271,G18272,G18273,G18274,G18275,G18276,G18277,G18278,G18279,G18280,
       G18281,G18282,G18283,G18284,G18285,G18286,G18287,G18288,G18289,G18290,G18291,G18292,G18293,G18294,G18295,G18296,G18297,G18298,G18299,G18300,
       G18301,G18302,G18303,G18304,G18305,G18306,G18307,G18308,G18309,G18310,G18311,G18312,G18313,G18314,G18315,G18316,G18317,G18318,G18319,G18320,
       G18321,G18322,G18323,G18324,G18325,G18326,G18327,G18328,G18329,G18330,G18331,G18332,G18333,G18334,G18335,G18336,G18337,G18338,G18339,G18340,
       G18341,G18342,G18343,G18344,G18345,G18346,G18347,G18348,G18349,G18350,G18351,G18352,G18353,G18354,G18355,G18356,G18357,G18358,G18359,G18360,
       G18361,G18362,G18363,G18364,G18365,G18366,G18367,G18368,G18369,G18370,G18371,G18372,G18373,G18374,G18375,G18376,G18377,G18378,G18379,G18380,
       G18381,G18382,G18383,G18384,G18385,G18386,G18387,G18388,G18389,G18390,G18391,G18392,G18393,G18394,G18395,G18396,G18397,G18398,G18399,G18400,
       G18401,G18402,G18403,G18404,G18405,G18406,G18407,G18408,G18409,G18410,G18411,G18412,G18413,G18414,G18415,G18416,G18417,G18418,G18419,G18420,
       G18421,G18422,G18423,G18424,G18425,G18426,G18427,G18428,G18429,G18430,G18431,G18432,G18433,G18434,G18435,G18436,G18437,G18438,G18439,G18440,
       G18441,G18442,G18443,G18444,G18445,G18446,G18447,G18448,G18449,G18450,G18451,G18452,G18453,G18454,G18455,G18456,G18457,G18458,G18459,G18460,
       G18461,G18462,G18463,G18464,G18465,G18466,G18467,G18468,G18469,G18470,G18471,G18472,G18473,G18474,G18475,G18476,G18477,G18478,G18479,G18480,
       G18481,G18482,G18483,G18484,G18485,G18486,G18487,G18488,G18489,G18490,G18491,G18492,G18493,G18494,G18495,G18496,G18497,G18498,G18499,G18500,
       G18501,G18502,G18503,G18504,G18505,G18506,G18507,G18508,G18509,G18510,G18511,G18512,G18513,G18514,G18515,G18516,G18517,G18518,G18519,G18520,
       G18521,G18522,G18523,G18524,G18525,G18526,G18527,G18528,G18529,G18530,G18531,G18532,G18533,G18534,G18535,G18536,G18537,G18538,G18539,G18540,
       G18541,G18542,G18543,G18544,G18545,G18546,G18547,G18548,G18549,G18550,G18551,G18552,G18553,G18554,G18555,G18556,G18557,G18558,G18559,G18560,
       G18561,G18562,G18563,G18564,G18565,G18566,G18567,G18568,G18569,G18570,G18571,G18572,G18573,G18574,G18575,G18576,G18577,G18578,G18579,G18580,
       G18581,G18582,G18583,G18584,G18585,G18586,G18587,G18588,G18589,G18590,G18591,G18592,G18593,G18594,G18595,G18596,G18597,G18598,G18599,G18600,
       G18601,G18602,G18603,G18604,G18605,G18606,G18607,G18608,G18609,G18610,G18611,G18612,G18613,G18614,G18615,G18616,G18617,G18618,G18619,G18620,
       G18621,G18622,G18623,G18624,G18625,G18626,G18627,G18628,G18629,G18630,G18631,G18632,G18633,G18634,G18635,G18636,G18637,G18638,G18639,G18640,
       G18641,G18642,G18643,G18644,G18645,G18646,G18647,G18648,G18649,G18650,G18651,G18652,G18653,G18654,G18655,G18656,G18657,G18658,G18659,G18660,
       G18661,G18662,G18663,G18664,G18665,G18666,G18667,G18668,G18669,G18670,G18671,G18672,G18673,G18674,G18675,G18676,G18677,G18678,G18679,G18680,
       G18681,G18682,G18683,G18684,G18685,G18686,G18687,G18688,G18689,G18690,G18691,G18692,G18693,G18694,G18695,G18696,G18697,G18698,G18699,G18700,
       G18701,G18702,G18703,G18704,G18705,G18706,G18707,G18708,G18709,G18710,G18711,G18712,G18713,G18714,G18715,G18716,G18717,G18718,G18719,G18720,
       G18721,G18722,G18723,G18724,G18725,G18726,G18727,G18728,G18729,G18730,G18731,G18732,G18733,G18734,G18735,G18736,G18737,G18738,G18739,G18740,
       G18741,G18742,G18743,G18744,G18745,G18746,G18747,G18748,G18749,G18750,G18751,G18752,G18753,G18754,G18755,G18756,G18757,G18758,G18759,G18760,
       G18761,G18762,G18763,G18764,G18765,G18766,G18767,G18768,G18769,G18770,G18771,G18772,G18773,G18774,G18775,G18776,G18777,G18778,G18779,G18780,
       G18781,G18782,G18783,G18784,G18785,G18786,G18787,G18788,G18789,G18790,G18791,G18792,G18793,G18794,G18795,G18796,G18797,G18798,G18799,G18800,
       G18801,G18802,G18803,G18804,G18805,G18806,G18807,G18808,G18809,G18810,G18811,G18812,G18813,G18814,G18815,G18816,G18817,G18818,G18819,G18820,
       G18821,G18822,G18823,G18824,G18825,G18826,G18827,G18828,G18829,G18830,G18831,G18832,G18833,G18834,G18835,G18836,G18837,G18838,G18839,G18840,
       G18841,G18842,G18843,G18844,G18845,G18846,G18847,G18848,G18849,G18850,G18851,G18852,G18853,G18854,G18855,G18856,G18857,G18858,G18859,G18860,
       G18861,G18862,G18863,G18864,G18865,G18866,G18867,G18868,G18869,G18870,G18871,G18872,G18873,G18874,G18875,G18876,G18877,G18878,G18879,G18880,
       G18881,G18882,G18883,G18884,G18885,G18886,G18887,G18888,G18889,G18890,G18891,G18892,G18893,G18894,G18895,G18896,G18897,G18898,G18899,G18900,
       G18901,G18902,G18903,G18904,G18905,G18906,G18907,G18908,G18909,G18910,G18911,G18912,G18913,G18914,G18915,G18916,G18917,G18918,G18919,G18920,
       G18921,G18922,G18923,G18924,G18925,G18926,G18927,G18928,G18929,G18930,G18931,G18932,G18933,G18934,G18935,G18936,G18937,G18938,G18939,G18940,
       G18941,G18942,G18943,G18944,G18945,G18946,G18947,G18948,G18949,G18950,G18951,G18952,G18953,G18954,G18955,G18956,G18957,G18958,G18959,G18960,
       G18961,G18962,G18963,G18964,G18965,G18966,G18967,G18968,G18969,G18970,G18971,G18972,G18973,G18974,G18975,G18976,G18977,G18978,G18979,G18980,
       G18981,G18982,G18983,G18984,G18985,G18986,G18987,G18988,G18989,G18990,G18991,G18992,G18993,G18994,G18995,G18996,G18997,G18998,G18999,G19000,
       G19001,G19002,G19003,G19004,G19005,G19006,G19007,G19008,G19009,G19010,G19011,G19012,G19013,G19014,G19015,G19016,G19017,G19018,G19019,G19020,
       G19021,G19022,G19023,G19024,G19025,G19026,G19027,G19028,G19029,G19030,G19031,G19032,G19033,G19034,G19035,G19036,G19037,G19038,G19039,G19040,
       G19041,G19042,G19043,G19044,G19045,G19046,G19047,G19048,G19049,G19050,G19051,G19052,G19053,G19054,G19055,G19056,G19057,G19058,G19059,G19060,
       G19061,G19062,G19063,G19064,G19065,G19066,G19067,G19068,G19069,G19070,G19071,G19072,G19073,G19074,G19075,G19076,G19077,G19078,G19079,G19080,
       G19081,G19082,G19083,G19084,G19085,G19086,G19087,G19088,G19089,G19090,G19091,G19092,G19093,G19094,G19095,G19096,G19097,G19098,G19099,G19100,
       G19101,G19102,G19103,G19104,G19105,G19106,G19107,G19108,G19109,G19110,G19111,G19112,G19113,G19114,G19115,G19116,G19117,G19118,G19119,G19120,
       G19121,G19122,G19123,G19124,G19125,G19126,G19127,G19128,G19129,G19130,G19131,G19132,G19133,G19134,G19135,G19136,G19137,G19138,G19139,G19140,
       G19141,G19142,G19143,G19144,G19145,G19146,G19147,G19148,G19149,G19150,G19151,G19152,G19153,G19154,G19155,G19156,G19157,G19158,G19159,G19160,
       G19161,G19162,G19163,G19164,G19165,G19166,G19167,G19168,G19169,G19170,G19171,G19172,G19173,G19174,G19175,G19176,G19177,G19178,G19179,G19180,
       G19181,G19182,G19183,G19184,G19185,G19186,G19187,G19188,G19189,G19190,G19191,G19192,G19193,G19194,G19195,G19196,G19197,G19198,G19199,G19200,
       G19201,G19202,G19203,G19204,G19205,G19206,G19207,G19208,G19209,G19210,G19211,G19212,G19213,G19214,G19215,G19216,G19217,G19218,G19219,G19220,
       G19221,G19222,G19223,G19224,G19225,G19226,G19227,G19228,G19229,G19230,G19231,G19232,G19233,G19234,G19235,G19236,G19237,G19238,G19239,G19240,
       G19241,G19242,G19243,G19244,G19245,G19246,G19247,G19248,G19249,G19250,G19251,G19252,G19253,G19254,G19255,G19256,G19257,G19258,G19259,G19260,
       G19261,G19262,G19263,G19264,G19265,G19266,G19267,G19268,G19269,G19270,G19271,G19272,G19273,G19274,G19275,G19276,G19277,G19278,G19279,G19280,
       G19281,G19282,G19283,G19284,G19285,G19286,G19287,G19288,G19289,G19290,G19291,G19292,G19293,G19294,G19295,G19296,G19297,G19298,G19299,G19300,
       G19301,G19302,G19303,G19304,G19305,G19306,G19307,G19308,G19309,G19310,G19311,G19312,G19313,G19314,G19315,G19316,G19317,G19318,G19319,G19320,
       G19321,G19322,G19323,G19324,G19325,G19326,G19327,G19328,G19329,G19330,G19331,G19332,G19333,G19334,G19335,G19336,G19337,G19338,G19339,G19340,
       G19341,G19342,G19343,G19344,G19345,G19346,G19347,G19348,G19349,G19350,G19351,G19352,G19353,G19354,G19355,G19356,G19357,G19358,G19359,G19360,
       G19361,G19362,G19363,G19364,G19365,G19366,G19367,G19368,G19369,G19370,G19371,G19372,G19373,G19374,G19375,G19376,G19377,G19378,G19379,G19380,
       G19381,G19382,G19383,G19384,G19385,G19386,G19387,G19388,G19389,G19390,G19391,G19392,G19393,G19394,G19395,G19396,G19397,G19398,G19399,G19400,
       G19401,G19402,G19403,G19404,G19405,G19406,G19407,G19408,G19409,G19410,G19411,G19412,G19413,G19414,G19415,G19416,G19417,G19418,G19419,G19420,
       G19421,G19422,G19423,G19424,G19425,G19426,G19427,G19428,G19429,G19430,G19431,G19432,G19433,G19434,G19435,G19436,G19437,G19438,G19439,G19440,
       G19441,G19442,G19443,G19444,G19445,G19446,G19447,G19448,G19449,G19450,G19451,G19452,G19453,G19454,G19455,G19456,G19457,G19458,G19459,G19460,
       G19461,G19462,G19463,G19464,G19465,G19466,G19467,G19468,G19469,G19470,G19471,G19472,G19473,G19474,G19475,G19476,G19477,G19478,G19479,G19480,
       G19481,G19482,G19483,G19484,G19485,G19486,G19487,G19488,G19489,G19490,G19491,G19492,G19493,G19494,G19495,G19496,G19497,G19498,G19499,G19500,
       G19501,G19502,G19503,G19504,G19505,G19506,G19507,G19508,G19509,G19510,G19511,G19512,G19513,G19514,G19515,G19516,G19517,G19518,G19519,G19520,
       G19521,G19522,G19523,G19524,G19525,G19526,G19527,G19528,G19529,G19530,G19531,G19532,G19533,G19534,G19535,G19536,G19537,G19538,G19539,G19540,
       G19541,G19542,G19543,G19544,G19545,G19546,G19547,G19548,G19549,G19550,G19551,G19552,G19553,G19554,G19555,G19556,G19557,G19558,G19559,G19560,
       G19561,G19562,G19563,G19564,G19565,G19566,G19567,G19568,G19569,G19570,G19571,G19572,G19573,G19574,G19575,G19576,G19577,G19578,G19579,G19580,
       G19581,G19582,G19583,G19584,G19585,G19586,G19587,G19588,G19589,G19590,G19591,G19592,G19593,G19594,G19595,G19596,G19597,G19598,G19599,G19600,
       G19601,G19602,G19603,G19604,G19605,G19606,G19607,G19608,G19609,G19610,G19611,G19612,G19613,G19614,G19615,G19616,G19617,G19618,G19619,G19620,
       G19621,G19622,G19623,G19624,G19625,G19626,G19627,G19628,G19629,G19630,G19631,G19632,G19633,G19634,G19635,G19636,G19637,G19638,G19639,G19640,
       G19641,G19642,G19643,G19644,G19645,G19646,G19647,G19648,G19649,G19650,G19651,G19652,G19653,G19654,G19655,G19656,G19657,G19658,G19659,G19660,
       G19661,G19662,G19663,G19664,G19665,G19666,G19667,G19668,G19669,G19670,G19671,G19672,G19673,G19674,G19675,G19676,G19677,G19678,G19679,G19680,
       G19681,G19682,G19683,G19684,G19685,G19686,G19687,G19688,G19689,G19690,G19691,G19692,G19693,G19694,G19695,G19696,G19697,G19698,G19699,G19700,
       G19701,G19702,G19703,G19704,G19705,G19706,G19707,G19708,G19709,G19710,G19711,G19712,G19713,G19714,G19715,G19716,G19717,G19718,G19719,G19720,
       G19721,G19722,G19723,G19724,G19725,G19726,G19727,G19728,G19729,G19730,G19731,G19732,G19733,G19734,G19735,G19736,G19737,G19738,G19739,G19740,
       G19741,G19742,G19743,G19744,G19745,G19746,G19747,G19748,G19749,G19750,G19751,G19752,G19753,G19754,G19755,G19756,G19757,G19758,G19759,G19760,
       G19761,G19762,G19763,G19764,G19765,G19766,G19767,G19768,G19769,G19770,G19771,G19772,G19773,G19774,G19775,G19776,G19777,G19778,G19779,G19780,
       G19781,G19782,G19783,G19784,G19785,G19786,G19787,G19788,G19789,G19790,G19791,G19792,G19793,G19794,G19795,G19796,G19797,G19798,G19799,G19800,
       G19801,G19802,G19803,G19804,G19805,G19806,G19807,G19808,G19809,G19810,G19811,G19812,G19813,G19814,G19815,G19816,G19817,G19818,G19819,G19820,
       G19821,G19822,G19823,G19824,G19825,G19826,G19827,G19828,G19829,G19830,G19831,G19832,G19833,G19834,G19835,G19836,G19837,G19838,G19839,G19840,
       G19841,G19842,G19843,G19844,G19845,G19846,G19847,G19848,G19849,G19850,G19851,G19852,G19853,G19854,G19855,G19856,G19857,G19858,G19859,G19860,
       G19861,G19862,G19863,G19864,G19865,G19866,G19867,G19868,G19869,G19870,G19871,G19872,G19873,G19874,G19875,G19876,G19877,G19878,G19879,G19880,
       G19881,G19882,G19883,G19884,G19885,G19886,G19887,G19888,G19889,G19890,G19891,G19892,G19893,G19894,G19895,G19896,G19897,G19898,G19899,G19900,
       G19901,G19902,G19903,G19904,G19905,G19906,G19907,G19908,G19909,G19910,G19911,G19912,G19913,G19914,G19915,G19916,G19917,G19918,G19919,G19920,
       G19921,G19922,G19923,G19924,G19925,G19926,G19927,G19928,G19929,G19930,G19931,G19932,G19933,G19934,G19935,G19936,G19937,G19938,G19939,G19940,
       G19941,G19942,G19943,G19944,G19945,G19946,G19947,G19948,G19949,G19950,G19951,G19952,G19953,G19954,G19955,G19956,G19957,G19958,G19959,G19960,
       G19961,G19962,G19963,G19964,G19965,G19966,G19967,G19968,G19969,G19970,G19971,G19972,G19973,G19974,G19975,G19976,G19977,G19978,G19979,G19980,
       G19981,G19982,G19983,G19984,G19985,G19986,G19987,G19988,G19989,G19990,G19991,G19992,G19993,G19994,G19995,G19996,G19997,G19998,G19999,G20000,
       G20001,G20002,G20003,G20004,G20005,G20006,G20007,G20008,G20009,G20010,G20011,G20012,G20013,G20014,G20015,G20016,G20017,G20018,G20019,G20020,
       G20021,G20022,G20023,G20024,G20025,G20026,G20027,G20028,G20029,G20030,G20031,G20032,G20033,G20034,G20035,G20036,G20037,G20038,G20039,G20040,
       G20041,G20042,G20043,G20044,G20045,G20046,G20047,G20048,G20049,G20050,G20051,G20052,G20053,G20054,G20055,G20056,G20057,G20058,G20059,G20060,
       G20061,G20062,G20063,G20064,G20065,G20066,G20067,G20068,G20069,G20070,G20071,G20072,G20073,G20074,G20075,G20076,G20077,G20078,G20079,G20080,
       G20081,G20082,G20083,G20084,G20085,G20086,G20087,G20088,G20089,G20090,G20091,G20092,G20093,G20094,G20095,G20096,G20097,G20098,G20099,G20100,
       G20101,G20102,G20103,G20104,G20105,G20106,G20107,G20108,G20109,G20110,G20111,G20112,G20113,G20114,G20115,G20116,G20117,G20118,G20119,G20120,
       G20121,G20122,G20123,G20124,G20125,G20126,G20127,G20128,G20129,G20130,G20131,G20132,G20133,G20134,G20135,G20136,G20137,G20138,G20139,G20140,
       G20141,G20142,G20143,G20144,G20145,G20146,G20147,G20148,G20149,G20150,G20151,G20152,G20153,G20154,G20155,G20156,G20157,G20158,G20159,G20160,
       G20161,G20162,G20163,G20164,G20165,G20166,G20167,G20168,G20169,G20170,G20171,G20172,G20173,G20174,G20175,G20176,G20177,G20178,G20179,G20180,
       G20181,G20182,G20183,G20184,G20185,G20186,G20187,G20188,G20189,G20190,G20191,G20192,G20193,G20194,G20195,G20196,G20197,G20198,G20199,G20200,
       G20201,G20202,G20203,G20204,G20205,G20206,G20207,G20208,G20209,G20210,G20211,G20212,G20213,G20214,G20215,G20216,G20217,G20218,G20219,G20220,
       G20221,G20222,G20223,G20224,G20225,G20226,G20227,G20228,G20229,G20230,G20231,G20232,G20233,G20234,G20235,G20236,G20237,G20238,G20239,G20240,
       G20241,G20242,G20243,G20244,G20245,G20246,G20247,G20248,G20249,G20250,G20251,G20252,G20253,G20254,G20255,G20256,G20257,G20258,G20259,G20260,
       G20261,G20262,G20263,G20264,G20265,G20266,G20267,G20268,G20269,G20270,G20271,G20272,G20273,G20274,G20275,G20276,G20277,G20278,G20279,G20280,
       G20281,G20282,G20283,G20284,G20285,G20286,G20287,G20288,G20289,G20290,G20291,G20292,G20293,G20294,G20295,G20296,G20297,G20298,G20299,G20300,
       G20301,G20302,G20303,G20304,G20305,G20306,G20307,G20308,G20309,G20310,G20311,G20312,G20313,G20314,G20315,G20316,G20317,G20318,G20319,G20320,
       G20321,G20322,G20323,G20324,G20325,G20326,G20327,G20328,G20329,G20330,G20331,G20332,G20333,G20334,G20335,G20336,G20337,G20338,G20339,G20340,
       G20341,G20342,G20343,G20344,G20345,G20346,G20347,G20348,G20349,G20350,G20351,G20352,G20353,G20354,G20355,G20356,G20357,G20358,G20359,G20360,
       G20361,G20362,G20363,G20364,G20365,G20366,G20367,G20368,G20369,G20370,G20371,G20372,G20373,G20374,G20375,G20376,G20377,G20378,G20379,G20380,
       G20381,G20382,G20383,G20384,G20385,G20386,G20387,G20388,G20389,G20390,G20391,G20392,G20393,G20394,G20395,G20396,G20397,G20398,G20399,G20400,
       G20401,G20402,G20403,G20404,G20405,G20406,G20407,G20408,G20409,G20410,G20411,G20412,G20413,G20414,G20415,G20416,G20417,G20418,G20419,G20420,
       G20421,G20422,G20423,G20424,G20425,G20426,G20427,G20428,G20429,G20430,G20431,G20432,G20433,G20434,G20435,G20436,G20437,G20438,G20439,G20440,
       G20441,G20442,G20443,G20444,G20445,G20446,G20447,G20448,G20449,G20450,G20451,G20452,G20453,G20454,G20455,G20456,G20457,G20458,G20459,G20460,
       G20461,G20462,G20463,G20464,G20465,G20466,G20467,G20468,G20469,G20470,G20471,G20472,G20473,G20474,G20475,G20476,G20477,G20478,G20479,G20480,
       G20481,G20482,G20483,G20484,G20485,G20486,G20487,G20488,G20489,G20490,G20491,G20492,G20493,G20494,G20495,G20496,G20497,G20498,G20499,G20500,
       G20501,G20502,G20503,G20504,G20505,G20506,G20507,G20508,G20509,G20510,G20511,G20512,G20513,G20514,G20515,G20516,G20517,G20518,G20519,G20520,
       G20521,G20522,G20523,G20524,G20525,G20526,G20527,G20528,G20529,G20530,G20531,G20532,G20533,G20534,G20535,G20536,G20537,G20538,G20539,G20540,
       G20541,G20542,G20543,G20544,G20545,G20546,G20547,G20548,G20549,G20550,G20551,G20552,G20553,G20554,G20555,G20556,G20557,G20558,G20559,G20560,
       G20561,G20562,G20563,G20564,G20565,G20566,G20567,G20568,G20569,G20570,G20571,G20572,G20573,G20574,G20575,G20576,G20577,G20578,G20579,G20580,
       G20581,G20582,G20583,G20584,G20585,G20586,G20587,G20588,G20589,G20590,G20591,G20592,G20593,G20594,G20595,G20596,G20597,G20598,G20599,G20600,
       G20601,G20602,G20603,G20604,G20605,G20606,G20607,G20608,G20609,G20610,G20611,G20612,G20613,G20614,G20615,G20616,G20617,G20618,G20619,G20620,
       G20621,G20622,G20623,G20624,G20625,G20626,G20627,G20628,G20629,G20630,G20631,G20632,G20633,G20634,G20635,G20636,G20637,G20638,G20639,G20640,
       G20641,G20642,G20643,G20644,G20645,G20646,G20647,G20648,G20649,G20650,G20651,G20652,G20653,G20654,G20655,G20656,G20657,G20658,G20659,G20660,
       G20661,G20662,G20663,G20664,G20665,G20666,G20667,G20668,G20669,G20670,G20671,G20672,G20673,G20674,G20675,G20676,G20677,G20678,G20679,G20680,
       G20681,G20682,G20683,G20684,G20685,G20686,G20687,G20688,G20689,G20690,G20691,G20692,G20693,G20694,G20695,G20696,G20697,G20698,G20699,G20700,
       G20701,G20702,G20703,G20704,G20705,G20706,G20707,G20708,G20709,G20710,G20711,G20712,G20713,G20714,G20715,G20716,G20717,G20718,G20719,G20720,
       G20721,G20722,G20723,G20724,G20725,G20726,G20727,G20728,G20729,G20730,G20731,G20732,G20733,G20734,G20735,G20736,G20737,G20738,G20739,G20740,
       G20741,G20742,G20743,G20744,G20745,G20746,G20747,G20748,G20749,G20750,G20751,G20752,G20753,G20754,G20755,G20756,G20757,G20758,G20759,G20760,
       G20761,G20762,G20763,G20764,G20765,G20766,G20767,G20768,G20769,G20770,G20771,G20772,G20773,G20774,G20775,G20776,G20777,G20778,G20779,G20780,
       G20781,G20782,G20783,G20784,G20785,G20786,G20787,G20788,G20789,G20790,G20791,G20792,G20793,G20794,G20795,G20796,G20797,G20798,G20799,G20800,
       G20801,G20802,G20803,G20804,G20805,G20806,G20807,G20808,G20809,G20810,G20811,G20812,G20813,G20814,G20815,G20816,G20817,G20818,G20819,G20820,
       G20821,G20822,G20823,G20824,G20825,G20826,G20827,G20828,G20829,G20830,G20831,G20832,G20833,G20834,G20835,G20836,G20837,G20838,G20839,G20840,
       G20841,G20842,G20843,G20844,G20845,G20846,G20847,G20848,G20849,G20850,G20851,G20852,G20853,G20854,G20855,G20856,G20857,G20858,G20859,G20860,
       G20861,G20862,G20863,G20864,G20865,G20866,G20867,G20868,G20869,G20870,G20871,G20872,G20873,G20874,G20875,G20876,G20877,G20878,G20879,G20880,
       G20881,G20882,G20883,G20884,G20885,G20886,G20887,G20888,G20889,G20890,G20891,G20892,G20893,G20894,G20895,G20896,G20897,G20898,G20899,G20900,
       G20901,G20902,G20903,G20904,G20905,G20906,G20907,G20908,G20909,G20910,G20911,G20912,G20913,G20914,G20915,G20916,G20917,G20918,G20919,G20920,
       G20921,G20922,G20923,G20924,G20925,G20926,G20927,G20928,G20929,G20930,G20931,G20932,G20933,G20934,G20935,G20936,G20937,G20938,G20939,G20940,
       G20941,G20942,G20943,G20944,G20945,G20946,G20947,G20948,G20949,G20950,G20951,G20952,G20953,G20954,G20955,G20956,G20957,G20958,G20959,G20960,
       G20961,G20962,G20963,G20964,G20965,G20966,G20967,G20968,G20969,G20970,G20971,G20972,G20973,G20974,G20975,G20976,G20977,G20978,G20979,G20980,
       G20981,G20982,G20983,G20984,G20985,G20986,G20987,G20988,G20989,G20990,G20991,G20992,G20993,G20994,G20995,G20996,G20997,G20998,G20999,G21000,
       G21001,G21002,G21003,G21004,G21005,G21006,G21007,G21008,G21009,G21010,G21011,G21012,G21013,G21014,G21015,G21016,G21017,G21018,G21019,G21020,
       G21021,G21022,G21023,G21024,G21025,G21026,G21027,G21028,G21029,G21030,G21031,G21032,G21033,G21034,G21035,G21036,G21037,G21038,G21039,G21040,
       G21041,G21042,G21043,G21044,G21045,G21046,G21047,G21048,G21049,G21050,G21051,G21052,G21053,G21054,G21055,G21056,G21057,G21058,G21059,G21060,
       G21061,G21062,G21063,G21064,G21065,G21066,G21067,G21068,G21069,G21070,G21071,G21072,G21073,G21074,G21075,G21076,G21077,G21078,G21079,G21080,
       G21081,G21082,G21083,G21084,G21085,G21086,G21087,G21088,G21089,G21090,G21091,G21092,G21093,G21094,G21095,G21096,G21097,G21098,G21099,G21100,
       G21101,G21102,G21103,G21104,G21105,G21106,G21107,G21108,G21109,G21110,G21111,G21112,G21113,G21114,G21115,G21116,G21117,G21118,G21119,G21120,
       G21121,G21122,G21123,G21124,G21125,G21126,G21127,G21128,G21129,G21130,G21131,G21132,G21133,G21134,G21135,G21136,G21137,G21138,G21139,G21140,
       G21141,G21142,G21143,G21144,G21145,G21146,G21147,G21148,G21149,G21150,G21151,G21152,G21153,G21154,G21155,G21156,G21157,G21158,G21159,G21160,
       G21161,G21162,G21163,G21164,G21165,G21166,G21167,G21168,G21169,G21170,G21171,G21172,G21173,G21174,G21175,G21176,G21177,G21178,G21179,G21180,
       G21181,G21182,G21183,G21184,G21185,G21186,G21187,G21188,G21189,G21190,G21191,G21192,G21193,G21194,G21195,G21196,G21197,G21198,G21199,G21200,
       G21201,G21202,G21203,G21204,G21205,G21206,G21207,G21208,G21209,G21210,G21211,G21212,G21213,G21214,G21215,G21216,G21217,G21218,G21219,G21220,
       G21221,G21222,G21223,G21224,G21225,G21226,G21227,G21228,G21229,G21230,G21231,G21232,G21233,G21234,G21235,G21236,G21237,G21238,G21239,G21240,
       G21241,G21242,G21243,G21244,G21245,G21246,G21247,G21248,G21249,G21250,G21251,G21252,G21253,G21254,G21255,G21256,G21257,G21258,G21259,G21260,
       G21261,G21262,G21263,G21264,G21265,G21266,G21267,G21268,G21269,G21270,G21271,G21272,G21273,G21274,G21275,G21276,G21277,G21278,G21279,G21280,
       G21281,G21282,G21283,G21284,G21285,G21286,G21287,G21288,G21289,G21290,G21291,G21292,G21293,G21294,G21295,G21296,G21297,G21298,G21299,G21300,
       G21301,G21302,G21303,G21304,G21305,G21306,G21307,G21308,G21309,G21310,G21311,G21312,G21313,G21314,G21315,G21316,G21317,G21318,G21319,G21320,
       G21321,G21322,G21323,G21324,G21325,G21326,G21327,G21328,G21329,G21330,G21331,G21332,G21333,G21334,G21335,G21336,G21337,G21338,G21339,G21340,
       G21341,G21342,G21343,G21344,G21345,G21346,G21347,G21348,G21349,G21350,G21351,G21352,G21353,G21354,G21355,G21356,G21357,G21358,G21359,G21360,
       G21361,G21362,G21363,G21364,G21365,G21366,G21367,G21368,G21369,G21370,G21371,G21372,G21373,G21374,G21375,G21376,G21377,G21378,G21379,G21380,
       G21381,G21382,G21383,G21384,G21385,G21386,G21387,G21388,G21389,G21390,G21391,G21392,G21393,G21394,G21395,G21396,G21397,G21398,G21399,G21400,
       G21401,G21402,G21403,G21404,G21405,G21406,G21407,G21408,G21409,G21410,G21411,G21412,G21413,G21414,G21415,G21416,G21417,G21418,G21419,G21420,
       G21421,G21422,G21423,G21424,G21425,G21426,G21427,G21428,G21429,G21430,G21431,G21432,G21433,G21434,G21435,G21436,G21437,G21438,G21439,G21440,
       G21441,G21442,G21443,G21444,G21445,G21446,G21447,G21448,G21449,G21450,G21451,G21452,G21453,G21454,G21455,G21456,G21457,G21458,G21459,G21460,
       G21461,G21462,G21463,G21464,G21465,G21466,G21467,G21468,G21469,G21470,G21471,G21472,G21473,G21474,G21475,G21476,G21477,G21478,G21479,G21480,
       G21481,G21482,G21483,G21484,G21485,G21486,G21487,G21488,G21489,G21490,G21491,G21492,G21493,G21494,G21495,G21496,G21497,G21498,G21499,G21500,
       G21501,G21502,G21503,G21504,G21505,G21506,G21507,G21508,G21509,G21510,G21511,G21512,G21513,G21514,G21515,G21516,G21517,G21518,G21519,G21520,
       G21521,G21522,G21523,G21524,G21525,G21526,G21527,G21528,G21529,G21530,G21531,G21532,G21533,G21534,G21535,G21536,G21537,G21538,G21539,G21540,
       G21541,G21542,G21543,G21544,G21545,G21546,G21547,G21548,G21549,G21550,G21551,G21552,G21553,G21554,G21555,G21556,G21557,G21558,G21559,G21560,
       G21561,G21562,G21563,G21564,G21565,G21566,G21567,G21568,G21569,G21570,G21571,G21572,G21573,G21574,G21575,G21576,G21577,G21578,G21579,G21580,
       G21581,G21582,G21583,G21584,G21585,G21586,G21587,G21588,G21589,G21590,G21591,G21592,G21593,G21594,G21595,G21596,G21597,G21598,G21599,G21600,
       G21601,G21602,G21603,G21604,G21605,G21606,G21607,G21608,G21609,G21610,G21611,G21612,G21613,G21614,G21615,G21616,G21617,G21618,G21619,G21620,
       G21621,G21622,G21623,G21624,G21625,G21626,G21627,G21628,G21629,G21630,G21631,G21632,G21633,G21634,G21635,G21636,G21637,G21638,G21639,G21640,
       G21641,G21642,G21643,G21644,G21645,G21646,G21647,G21648,G21649,G21650,G21651,G21652,G21653,G21654,G21655,G21656,G21657,G21658,G21659,G21660,
       G21661,G21662,G21663,G21664,G21665,G21666,G21667,G21668,G21669,G21670,G21671,G21672,G21673,G21674,G21675,G21676,G21677,G21678,G21679,G21680,
       G21681,G21682,G21683,G21684,G21685,G21686,G21687,G21688,G21689,G21690,G21691,G21692,G21693,G21694,G21695,G21696,G21697,G21698,G21699,G21700,
       G21701,G21702,G21703,G21704,G21705,G21706,G21707,G21708,G21709,G21710,G21711,G21712,G21713,G21714,G21715,G21716,G21717,G21718,G21719,G21720,
       G21721,G21722,G21723,G21724,G21725,G21726,G21727,G21728,G21729,G21730,G21731,G21732,G21733,G21734,G21735,G21736,G21737,G21738,G21739,G21740,
       G21741,G21742,G21743,G21744,G21745,G21746,G21747,G21748,G21749,G21750,G21751,G21752,G21753,G21754,G21755,G21756,G21757,G21758,G21759,G21760,
       G21761,G21762,G21763,G21764,G21765,G21766,G21767,G21768,G21769,G21770,G21771,G21772,G21773,G21774,G21775,G21776,G21777,G21778,G21779,G21780,
       G21781,G21782,G21783,G21784,G21785,G21786,G21787,G21788,G21789,G21790,G21791,G21792,G21793,G21794,G21795,G21796,G21797,G21798,G21799,G21800,
       G21801,G21802,G21803,G21804,G21805,G21806,G21807,G21808,G21809,G21810,G21811,G21812,G21813,G21814,G21815,G21816,G21817,G21818,G21819,G21820,
       G21821,G21822,G21823,G21824,G21825,G21826,G21827,G21828,G21829,G21830,G21831,G21832,G21833,G21834,G21835,G21836,G21837,G21838,G21839,G21840,
       G21841,G21842,G21843,G21844,G21845,G21846,G21847,G21848,G21849,G21850,G21851,G21852,G21853,G21854,G21855,G21856,G21857,G21858,G21859,G21860,
       G21861,G21862,G21863,G21864,G21865,G21866,G21867,G21868,G21869,G21870,G21871,G21872,G21873,G21874,G21875,G21876,G21877,G21878,G21879,G21880,
       G21881,G21882,G21883,G21884,G21885,G21886,G21887,G21888,G21889,G21890,G21891,G21892,G21893,G21894,G21895,G21896,G21897,G21898,G21899,G21900,
       G21901,G21902,G21903,G21904,G21905,G21906,G21907,G21908,G21909,G21910,G21911,G21912,G21913,G21914,G21915,G21916,G21917,G21918,G21919,G21920,
       G21921,G21922,G21923,G21924,G21925,G21926,G21927,G21928,G21929,G21930,G21931,G21932,G21933,G21934,G21935,G21936,G21937,G21938,G21939,G21940,
       G21941,G21942,G21943,G21944,G21945,G21946,G21947,G21948,G21949,G21950,G21951,G21952,G21953,G21954,G21955,G21956,G21957,G21958,G21959,G21960,
       G21961,G21962,G21963,G21964,G21965,G21966,G21967,G21968,G21969,G21970,G21971,G21972,G21973,G21974,G21975,G21976,G21977,G21978,G21979,G21980,
       G21981,G21982,G21983,G21984,G21985,G21986,G21987,G21988,G21989,G21990,G21991,G21992,G21993,G21994,G21995,G21996,G21997,G21998,G21999,G22000,
       G22001,G22002,G22003,G22004,G22005,G22006,G22007,G22008,G22009,G22010,G22011,G22012,G22013,G22014,G22015,G22016,G22017,G22018,G22019,G22020,
       G22021,G22022,G22023,G22024,G22025,G22026,G22027,G22028,G22029,G22030,G22031,G22032,G22033,G22034,G22035,G22036,G22037,G22038,G22039,G22040,
       G22041,G22042,G22043,G22044,G22045,G22046,G22047,G22048,G22049,G22050,G22051,G22052,G22053,G22054,G22055,G22056,G22057,G22058,G22059,G22060,
       G22061,G22062,G22063,G22064,G22065,G22066,G22067,G22068,G22069,G22070,G22071,G22072,G22073,G22074,G22075,G22076,G22077,G22078,G22079,G22080,
       G22081,G22082,G22083,G22084,G22085,G22086,G22087,G22088,G22089,G22090,G22091,G22092,G22093,G22094,G22095,G22096,G22097,G22098,G22099,G22100,
       G22101,G22102,G22103,G22104,G22105,G22106,G22107,G22108,G22109,G22110,G22111,G22112,G22113,G22114,G22115,G22116,G22117,G22118,G22119,G22120,
       G22121,G22122,G22123,G22124,G22125,G22126,G22127,G22128,G22129,G22130,G22131,G22132,G22133,G22134,G22135,G22136,G22137,G22138,G22139,G22140,
       G22141,G22142,G22143,G22144,G22145,G22146,G22147,G22148,G22149,G22150,G22151,G22152,G22153,G22154,G22155,G22156,G22157,G22158,G22159,G22160,
       G22161,G22162,G22163,G22164,G22165,G22166,G22167,G22168,G22169,G22170,G22171,G22172,G22173,G22174,G22175,G22176,G22177,G22178,G22179,G22180,
       G22181,G22182,G22183,G22184,G22185,G22186,G22187,G22188,G22189,G22190,G22191,G22192,G22193,G22194,G22195,G22196,G22197,G22198,G22199,G22200,
       G22201,G22202,G22203,G22204,G22205,G22206,G22207,G22208,G22209,G22210,G22211,G22212,G22213,G22214,G22215,G22216,G22217,G22218,G22219,G22220,
       G22221,G22222,G22223,G22224,G22225,G22226,G22227,G22228,G22229,G22230,G22231,G22232,G22233,G22234,G22235,G22236,G22237,G22238,G22239,G22240,
       G22241,G22242,G22243,G22244,G22245,G22246,G22247,G22248,G22249,G22250,G22251,G22252,G22253,G22254,G22255,G22256,G22257,G22258,G22259,G22260,
       G22261,G22262,G22263,G22264,G22265,G22266,G22267,G22268,G22269,G22270,G22271,G22272,G22273,G22274,G22275,G22276,G22277,G22278,G22279,G22280,
       G22281,G22282,G22283,G22284,G22285,G22286,G22287,G22288,G22289,G22290,G22291,G22292,G22293,G22294,G22295,G22296,G22297,G22298,G22299,G22300,
       G22301,G22302,G22303,G22304,G22305,G22306,G22307,G22308,G22309,G22310,G22311,G22312,G22313,G22314,G22315,G22316,G22317,G22318,G22319,G22320,
       G22321,G22322,G22323,G22324,G22325,G22326,G22327,G22328,G22329,G22330,G22331,G22332,G22333,G22334,G22335,G22336,G22337,G22338,G22339,G22340,
       G22341,G22342,G22343,G22344,G22345,G22346,G22347,G22348,G22349,G22350,G22351,G22352,G22353,G22354,G22355,G22356,G22357,G22358,G22359,G22360,
       G22361,G22362,G22363,G22364,G22365,G22366,G22367,G22368,G22369,G22370,G22371,G22372,G22373,G22374,G22375,G22376,G22377,G22378,G22379,G22380,
       G22381,G22382,G22383,G22384,G22385,G22386,G22387,G22388,G22389,G22390,G22391,G22392,G22393,G22394,G22395,G22396,G22397,G22398,G22399,G22400,
       G22401,G22402,G22403,G22404,G22405,G22406,G22407,G22408,G22409,G22410,G22411,G22412,G22413,G22414,G22415,G22416,G22417,G22418,G22419,G22420,
       G22421,G22422,G22423,G22424,G22425,G22426,G22427,G22428,G22429,G22430,G22431,G22432,G22433,G22434,G22435,G22436,G22437,G22438,G22439,G22440,
       G22441,G22442,G22443,G22444,G22445,G22446,G22447,G22448,G22449,G22450,G22451,G22452,G22453,G22454,G22455,G22456,G22457,G22458,G22459,G22460,
       G22461,G22462,G22463,G22464,G22465,G22466,G22467,G22468,G22469,G22470,G22471,G22472,G22473,G22474,G22475,G22476,G22477,G22478,G22479,G22480,
       G22481,G22482,G22483,G22484,G22485,G22486,G22487,G22488,G22489,G22490,G22491,G22492,G22493,G22494,G22495,G22496,G22497,G22498,G22499,G22500,
       G22501,G22502,G22503,G22504,G22505,G22506,G22507,G22508,G22509,G22510,G22511,G22512,G22513,G22514,G22515,G22516,G22517,G22518,G22519,G22520,
       G22521,G22522,G22523,G22524,G22525,G22526,G22527,G22528,G22529,G22530,G22531,G22532,G22533,G22534,G22535,G22536,G22537,G22538,G22539,G22540,
       G22541,G22542,G22543,G22544,G22545,G22546,G22547,G22548,G22549,G22550,G22551,G22552,G22553,G22554,G22555,G22556,G22557,G22558,G22559,G22560,
       G22561,G22562,G22563,G22564,G22565,G22566,G22567,G22568,G22569,G22570,G22571,G22572,G22573,G22574,G22575,G22576,G22577,G22578,G22579,G22580,
       G22581,G22582,G22583,G22584,G22585,G22586,G22587,G22588,G22589,G22590,G22591,G22592,G22593,G22594,G22595,G22596,G22597,G22598,G22599,G22600,
       G22601,G22602,G22603,G22604,G22605,G22606,G22607,G22608,G22609,G22610,G22611,G22612,G22613,G22614,G22615,G22616,G22617,G22618,G22619,G22620,
       G22621,G22622,G22623,G22624,G22625,G22626,G22627,G22628,G22629,G22630,G22631,G22632,G22633,G22634,G22635,G22636,G22637,G22638,G22639,G22640,
       G22641,G22642,G22643,G22644,G22645,G22646,G22647,G22648,G22649,G22650,G22651,G22652,G22653,G22654,G22655,G22656,G22657,G22658,G22659,G22660,
       G22661,G22662,G22663,G22664,G22665,G22666,G22667,G22668,G22669,G22670,G22671,G22672,G22673,G22674,G22675,G22676,G22677,G22678,G22679,G22680,
       G22681,G22682,G22683,G22684,G22685,G22686,G22687,G22688,G22689,G22690,G22691,G22692,G22693,G22694,G22695,G22696,G22697,G22698,G22699,G22700,
       G22701,G22702,G22703,G22704,G22705,G22706,G22707,G22708,G22709,G22710,G22711,G22712,G22713,G22714,G22715,G22716,G22717,G22718,G22719,G22720,
       G22721,G22722,G22723,G22724,G22725,G22726,G22727,G22728,G22729,G22730,G22731,G22732,G22733,G22734,G22735,G22736,G22737,G22738,G22739,G22740,
       G22741,G22742,G22743,G22744,G22745,G22746,G22747,G22748,G22749,G22750,G22751,G22752,G22753,G22754,G22755,G22756,G22757,G22758,G22759,G22760,
       G22761,G22762,G22763,G22764,G22765,G22766,G22767,G22768,G22769,G22770,G22771,G22772,G22773,G22774,G22775,G22776,G22777,G22778,G22779,G22780,
       G22781,G22782,G22783,G22784,G22785,G22786,G22787,G22788,G22789,G22790,G22791,G22792,G22793,G22794,G22795,G22796,G22797,G22798,G22799,G22800,
       G22801,G22802,G22803,G22804,G22805,G22806,G22807,G22808,G22809,G22810,G22811,G22812,G22813,G22814,G22815,G22816,G22817,G22818,G22819,G22820,
       G22821,G22822,G22823,G22824,G22825,G22826,G22827,G22828,G22829,G22830,G22831,G22832,G22833,G22834,G22835,G22836,G22837,G22838,G22839,G22840,
       G22841,G22842,G22843,G22844,G22845,G22846,G22847,G22848,G22849,G22850,G22851,G22852,G22853,G22854,G22855,G22856,G22857,G22858,G22859,G22860,
       G22861,G22862,G22863,G22864,G22865,G22866,G22867,G22868,G22869,G22870,G22871,G22872,G22873,G22874,G22875,G22876,G22877,G22878,G22879,G22880,
       G22881,G22882,G22883,G22884,G22885,G22886,G22887,G22888,G22889,G22890,G22891,G22892,G22893,G22894,G22895,G22896,G22897,G22898,G22899,G22900,
       G22901,G22902,G22903,G22904,G22905,G22906,G22907,G22908,G22909,G22910,G22911,G22912,G22913,G22914,G22915,G22916,G22917,G22918,G22919,G22920,
       G22921,G22922,G22923,G22924,G22925,G22926,G22927,G22928,G22929,G22930,G22931,G22932,G22933,G22934,G22935,G22936,G22937,G22938,G22939,G22940,
       G22941,G22942,G22943,G22944,G22945,G22946,G22947,G22948,G22949,G22950,G22951,G22952,G22953,G22954,G22955,G22956,G22957,G22958,G22959,G22960,
       G22961,G22962,G22963,G22964,G22965,G22966,G22967,G22968,G22969,G22970,G22971,G22972,G22973,G22974,G22975,G22976,G22977,G22978,G22979,G22980,
       G22981,G22982,G22983,G22984,G22985,G22986,G22987,G22988,G22989,G22990,G22991,G22992,G22993,G22994,G22995,G22996,G22997,G22998,G22999,G23000,
       G23001,G23002,G23003,G23004,G23005,G23006,G23007,G23008,G23009,G23010,G23011,G23012,G23013,G23014,G23015,G23016,G23017,G23018,G23019,G23020,
       G23021,G23022,G23023,G23024,G23025,G23026,G23027,G23028,G23029,G23030,G23031,G23032,G23033,G23034,G23035,G23036,G23037,G23038,G23039,G23040,
       G23041,G23042,G23043,G23044,G23045,G23046,G23047,G23048,G23049,G23050,G23051,G23052,G23053,G23054,G23055,G23056,G23057,G23058,G23059,G23060,
       G23061,G23062,G23063,G23064,G23065,G23066,G23067,G23068,G23069,G23070,G23071,G23072,G23073,G23074,G23075,G23076,G23077,G23078,G23079,G23080,
       G23081,G23082,G23083,G23084,G23085,G23086,G23087,G23088,G23089,G23090,G23091,G23092,G23093,G23094,G23095,G23096,G23097,G23098,G23099,G23100,
       G23101,G23102,G23103,G23104,G23105,G23106,G23107,G23108,G23109,G23110,G23111,G23112,G23113,G23114,G23115,G23116,G23117,G23118,G23119,G23120,
       G23121,G23122,G23123,G23124,G23125,G23126,G23127,G23128,G23129,G23130,G23131,G23132,G23133,G23134,G23135,G23136,G23137,G23138,G23139,G23140,
       G23141,G23142,G23143,G23144,G23145,G23146,G23147,G23148,G23149,G23150,G23151,G23152,G23153,G23154,G23155,G23156,G23157,G23158,G23159,G23160,
       G23161,G23162,G23163,G23164,G23165,G23166,G23167,G23168,G23169,G23170,G23171,G23172,G23173,G23174,G23175,G23176,G23177,G23178,G23179,G23180,
       G23181,G23182,G23183,G23184,G23185,G23186,G23187,G23188,G23189,G23190,G23191,G23192,G23193,G23194,G23195,G23196,G23197,G23198,G23199,G23200,
       G23201,G23202,G23203,G23204,G23205,G23206,G23207,G23208,G23209,G23210,G23211,G23212,G23213,G23214,G23215,G23216,G23217,G23218,G23219,G23220,
       G23221,G23222,G23223,G23224,G23225,G23226,G23227,G23228,G23229,G23230,G23231,G23232,G23233,G23234,G23235,G23236,G23237,G23238,G23239,G23240,
       G23241,G23242,G23243,G23244,G23245,G23246,G23247,G23248,G23249,G23250,G23251,G23252,G23253,G23254,G23255,G23256,G23257,G23258,G23259,G23260,
       G23261,G23262,G23263,G23264,G23265,G23266,G23267,G23268,G23269,G23270,G23271,G23272,G23273,G23274,G23275,G23276,G23277,G23278,G23279,G23280,
       G23281,G23282,G23283,G23284,G23285,G23286,G23287,G23288,G23289,G23290,G23291,G23292,G23293,G23294,G23295,G23296,G23297,G23298,G23299,G23300,
       G23301,G23302,G23303,G23304,G23305,G23306,G23307,G23308,G23309,G23310,G23311,G23312,G23313,G23314,G23315,G23316,G23317,G23318,G23319,G23320,
       G23321,G23322,G23323,G23324,G23325,G23326,G23327,G23328,G23329,G23330,G23331,G23332,G23333,G23334,G23335,G23336,G23337,G23338,G23339,G23340,
       G23341,G23342,G23343,G23344,G23345,G23346,G23347,G23348,G23349,G23350,G23351,G23352,G23353,G23354,G23355,G23356,G23357,G23358,G23359,G23360,
       G23361,G23362,G23363,G23364,G23365,G23366,G23367,G23368,G23369,G23370,G23371,G23372,G23373,G23374,G23375,G23376,G23377,G23378,G23379,G23380,
       G23381,G23382,G23383,G23384,G23385,G23386,G23387,G23388,G23389,G23390,G23391,G23392,G23393,G23394,G23395,G23396,G23397,G23398,G23399,G23400,
       G23401,G23402,G23403,G23404,G23405,G23406,G23407,G23408,G23409,G23410,G23411,G23412,G23413,G23414,G23415,G23416,G23417,G23418,G23419,G23420,
       G23421,G23422,G23423,G23424,G23425,G23426,G23427,G23428,G23429,G23430,G23431,G23432,G23433,G23434,G23435,G23436,G23437,G23438,G23439,G23440,
       G23441,G23442,G23443,G23444,G23445,G23446,G23447,G23448,G23449,G23450,G23451,G23452,G23453,G23454,G23455,G23456,G23457,G23458,G23459,G23460,
       G23461,G23462,G23463,G23464,G23465,G23466,G23467,G23468,G23469,G23470,G23471,G23472,G23473,G23474,G23475,G23476,G23477,G23478,G23479,G23480,
       G23481,G23482,G23483,G23484,G23485,G23486,G23487,G23488,G23489,G23490,G23491,G23492,G23493,G23494,G23495,G23496,G23497,G23498,G23499,G23500,
       G23501,G23502,G23503,G23504,G23505,G23506,G23507,G23508,G23509,G23510,G23511,G23512,G23513,G23514,G23515,G23516,G23517,G23518,G23519,G23520,
       G23521,G23522,G23523,G23524,G23525,G23526,G23527,G23528,G23529,G23530,G23531,G23532,G23533,G23534,G23535,G23536,G23537,G23538,G23539,G23540,
       G23541,G23542,G23543,G23544,G23545,G23546,G23547,G23548,G23549,G23550,G23551,G23552,G23553,G23554,G23555,G23556,G23557,G23558,G23559,G23560,
       G23561,G23562,G23563,G23564,G23565,G23566,G23567,G23568,G23569,G23570,G23571,G23572,G23573,G23574,G23575,G23576,G23577,G23578,G23579,G23580,
       G23581,G23582,G23583,G23584,G23585,G23586,G23587,G23588,G23589,G23590,G23591,G23592,G23593,G23594,G23595,G23596,G23597,G23598,G23599,G23600,
       G23601,G23602,G23603,G23604,G23605,G23606,G23607,G23608,G23609,G23610,G23611,G23612,G23613,G23614,G23615,G23616,G23617,G23618,G23619,G23620,
       G23621,G23622,G23623,G23624,G23625,G23626,G23627,G23628,G23629,G23630,G23631,G23632,G23633,G23634,G23635,G23636,G23637,G23638,G23639,G23640,
       G23641,G23642,G23643,G23644,G23645,G23646,G23647,G23648,G23649,G23650,G23651,G23652,G23653,G23654,G23655,G23656,G23657,G23658,G23659,G23660,
       G23661,G23662,G23663,G23664,G23665,G23666,G23667,G23668,G23669,G23670,G23671,G23672,G23673,G23674,G23675,G23676,G23677,G23678,G23679,G23680,
       G23681,G23682,G23683,G23684,G23685,G23686,G23687,G23688,G23689,G23690,G23691,G23692,G23693,G23694,G23695,G23696,G23697,G23698,G23699,G23700,
       G23701,G23702,G23703,G23704,G23705,G23706,G23707,G23708,G23709,G23710,G23711,G23712,G23713,G23714,G23715,G23716,G23717,G23718,G23719,G23720,
       G23721,G23722,G23723,G23724,G23725,G23726,G23727,G23728,G23729,G23730,G23731,G23732,G23733,G23734,G23735,G23736,G23737,G23738,G23739,G23740,
       G23741,G23742,G23743,G23744,G23745,G23746,G23747,G23748,G23749,G23750,G23751,G23752,G23753,G23754,G23755,G23756,G23757,G23758,G23759,G23760,
       G23761,G23762,G23763,G23764,G23765,G23766,G23767,G23768,G23769,G23770,G23771,G23772,G23773,G23774,G23775,G23776,G23777,G23778,G23779,G23780,
       G23781,G23782,G23783,G23784,G23785,G23786,G23787,G23788,G23789,G23790,G23791,G23792,G23793,G23794,G23795,G23796,G23797,G23798,G23799,G23800,
       G23801,G23802,G23803,G23804,G23805,G23806,G23807,G23808,G23809,G23810,G23811,G23812,G23813,G23814,G23815,G23816,G23817,G23818,G23819,G23820,
       G23821,G23822,G23823,G23824,G23825,G23826,G23827,G23828,G23829,G23830,G23831,G23832,G23833,G23834,G23835,G23836,G23837,G23838,G23839,G23840,
       G23841,G23842,G23843,G23844,G23845,G23846,G23847,G23848,G23849,G23850,G23851,G23852,G23853,G23854,G23855,G23856,G23857,G23858,G23859,G23860,
       G23861,G23862,G23863,G23864,G23865,G23866,G23867,G23868,G23869,G23870,G23871,G23872,G23873,G23874,G23875,G23876,G23877,G23878,G23879,G23880,
       G23881,G23882,G23883,G23884,G23885,G23886,G23887,G23888,G23889,G23890,G23891,G23892,G23893,G23894,G23895,G23896,G23897,G23898,G23899,G23900,
       G23901,G23902,G23903,G23904,G23905,G23906,G23907,G23908,G23909,G23910,G23911,G23912,G23913,G23914,G23915,G23916,G23917,G23918,G23919,G23920,
       G23921,G23922,G23923,G23924,G23925,G23926,G23927,G23928,G23929,G23930,G23931,G23932,G23933,G23934,G23935,G23936,G23937,G23938,G23939,G23940,
       G23941,G23942,G23943,G23944,G23945,G23946,G23947,G23948,G23949,G23950,G23951,G23952,G23953,G23954,G23955,G23956,G23957,G23958,G23959,G23960,
       G23961,G23962,G23963,G23964,G23965,G23966,G23967,G23968,G23969,G23970,G23971,G23972,G23973,G23974,G23975,G23976,G23977,G23978,G23979,G23980,
       G23981,G23982,G23983,G23984,G23985,G23986,G23987,G23988,G23989,G23990,G23991,G23992,G23993,G23994,G23995,G23996,G23997,G23998,G23999,G24000,
       G24001,G24002,G24003,G24004,G24005,G24006,G24007,G24008,G24009,G24010,G24011,G24012,G24013,G24014,G24015,G24016,G24017,G24018,G24019,G24020,
       G24021,G24022,G24023,G24024,G24025,G24026,G24027,G24028,G24029,G24030,G24031,G24032,G24033,G24034,G24035,G24036,G24037,G24038,G24039,G24040,
       G24041,G24042,G24043,G24044,G24045,G24046,G24047,G24048,G24049,G24050,G24051,G24052,G24053,G24054,G24055,G24056,G24057,G24058,G24059,G24060,
       G24061,G24062,G24063,G24064,G24065,G24066,G24067,G24068,G24069,G24070,G24071,G24072,G24073,G24074,G24075,G24076,G24077,G24078,G24079,G24080,
       G24081,G24082,G24083,G24084,G24085,G24086,G24087,G24088,G24089,G24090,G24091,G24092,G24093,G24094,G24095,G24096,G24097,G24098,G24099,G24100,
       G24101,G24102,G24103,G24104,G24105,G24106,G24107,G24108,G24109,G24110,G24111,G24112,G24113,G24114,G24115,G24116,G24117,G24118,G24119,G24120,
       G24121,G24122,G24123,G24124,G24125,G24126,G24127,G24128,G24129,G24130,G24131,G24132,G24133,G24134,G24135,G24136,G24137,G24138,G24139,G24140,
       G24141,G24142,G24143,G24144,G24145,G24146,G24147,G24148,G24149,G24150,G24151,G24152,G24153,G24154,G24155,G24156,G24157,G24158,G24159,G24160,
       G24161,G24162,G24163,G24164,G24165,G24166,G24167,G24168,G24169,G24170,G24171,G24172,G24173,G24174,G24175,G24176,G24177,G24178,G24179,G24180,
       G24181,G24182,G24183,G24184,G24185,G24186,G24187,G24188,G24189,G24190,G24191,G24192,G24193,G24194,G24195,G24196,G24197,G24198,G24199,G24200,
       G24201,G24202,G24203,G24204,G24205,G24206,G24207,G24208,G24209,G24210,G24211,G24212,G24213,G24214,G24215,G24216,G24217,G24218,G24219,G24220,
       G24221,G24222,G24223,G24224,G24225,G24226,G24227,G24228,G24229,G24230,G24231,G24232,G24233,G24234,G24235,G24236,G24237,G24238,G24239,G24240,
       G24241,G24242,G24243,G24244,G24245,G24246,G24247,G24248,G24249,G24250,G24251,G24252,G24253,G24254,G24255,G24256,G24257,G24258,G24259,G24260,
       G24261,G24262,G24263,G24264,G24265,G24266,G24267,G24268,G24269,G24270,G24271,G24272,G24273,G24274,G24275,G24276,G24277,G24278,G24279,G24280,
       G24281,G24282,G24283,G24284,G24285,G24286,G24287,G24288,G24289,G24290,G24291,G24292,G24293,G24294,G24295,G24296,G24297,G24298,G24299,G24300,
       G24301,G24302,G24303,G24304,G24305,G24306,G24307,G24308,G24309,G24310,G24311,G24312,G24313,G24314,G24315,G24316,G24317,G24318,G24319,G24320,
       G24321,G24322,G24323,G24324,G24325,G24326,G24327,G24328,G24329,G24330,G24331,G24332,G24333,G24334,G24335,G24336,G24337,G24338,G24339,G24340,
       G24341,G24342,G24343,G24344,G24345,G24346,G24347,G24348,G24349,G24350,G24351,G24352,G24353,G24354,G24355,G24356,G24357,G24358,G24359,G24360,
       G24361,G24362,G24363,G24364,G24365,G24366,G24367,G24368,G24369,G24370,G24371,G24372,G24373,G24374,G24375,G24376,G24377,G24378,G24379,G24380,
       G24381,G24382,G24383,G24384,G24385,G24386,G24387,G24388,G24389,G24390,G24391,G24392,G24393,G24394,G24395,G24396,G24397,G24398,G24399,G24400,
       G24401,G24402,G24403,G24404,G24405,G24406,G24407,G24408,G24409,G24410,G24411,G24412,G24413,G24414,G24415,G24416,G24417,G24418,G24419,G24420,
       G24421,G24422,G24423,G24424,G24425,G24426,G24427,G24428,G24429,G24430,G24431,G24432,G24433,G24434,G24435,G24436,G24437,G24438,G24439,G24440,
       G24441,G24442,G24443,G24444,G24445,G24446,G24447,G24448,G24449,G24450,G24451,G24452,G24453,G24454,G24455,G24456,G24457,G24458,G24459,G24460,
       G24461,G24462,G24463,G24464,G24465,G24466,G24467,G24468,G24469,G24470,G24471,G24472,G24473,G24474,G24475,G24476,G24477,G24478,G24479,G24480,
       G24481,G24482,G24483,G24484,G24485,G24486,G24487,G24488,G24489,G24490,G24491,G24492,G24493,G24494,G24495,G24496,G24497,G24498,G24499,G24500,
       G24501,G24502,G24503,G24504,G24505,G24506,G24507,G24508,G24509,G24510,G24511,G24512,G24513,G24514,G24515,G24516,G24517,G24518,G24519,G24520,
       G24521,G24522,G24523,G24524,G24525,G24526,G24527,G24528,G24529,G24530,G24531,G24532,G24533,G24534,G24535,G24536,G24537,G24538,G24539,G24540,
       G24541,G24542,G24543,G24544,G24545,G24546,G24547,G24548,G24549,G24550,G24551,G24552,G24553,G24554,G24555,G24556,G24557,G24558,G24559,G24560,
       G24561,G24562,G24563,G24564,G24565,G24566,G24567,G24568,G24569,G24570,G24571,G24572,G24573,G24574,G24575,G24576,G24577,G24578,G24579,G24580,
       G24581,G24582,G24583,G24584,G24585,G24586,G24587,G24588,G24589,G24590,G24591,G24592,G24593,G24594,G24595,G24596,G24597,G24598,G24599,G24600,
       G24601,G24602,G24603,G24604,G24605,G24606,G24607,G24608,G24609,G24610,G24611,G24612,G24613,G24614,G24615,G24616,G24617,G24618,G24619,G24620,
       G24621,G24622,G24623,G24624,G24625,G24626,G24627,G24628,G24629,G24630,G24631,G24632,G24633,G24634,G24635,G24636,G24637,G24638,G24639,G24640,
       G24641,G24642,G24643,G24644,G24645,G24646,G24647,G24648,G24649,G24650,G24651,G24652,G24653,G24654,G24655,G24656,G24657,G24658,G24659,G24660,
       G24661,G24662,G24663,G24664,G24665,G24666,G24667,G24668,G24669,G24670,G24671,G24672,G24673,G24674,G24675,G24676,G24677,G24678,G24679,G24680,
       G24681,G24682,G24683,G24684,G24685,G24686,G24687,G24688,G24689,G24690,G24691,G24692,G24693,G24694,G24695,G24696,G24697,G24698,G24699,G24700,
       G24701,G24702,G24703,G24704,G24705,G24706,G24707,G24708,G24709,G24710,G24711,G24712,G24713,G24714,G24715,G24716,G24717,G24718,G24719,G24720,
       G24721,G24722,G24723,G24724,G24725,G24726,G24727,G24728,G24729,G24730,G24731,G24732,G24733,G24734,G24735,G24736,G24737,G24738,G24739,G24740,
       G24741,G24742,G24743,G24744,G24745,G24746,G24747,G24748,G24749,G24750,G24751,G24752,G24753,G24754,G24755,G24756,G24757,G24758,G24759,G24760,
       G24761,G24762,G24763,G24764,G24765,G24766,G24767,G24768,G24769,G24770,G24771,G24772,G24773,G24774,G24775,G24776,G24777,G24778,G24779,G24780,
       G24781,G24782,G24783,G24784,G24785,G24786,G24787,G24788,G24789,G24790,G24791,G24792,G24793,G24794,G24795,G24796,G24797,G24798,G24799,G24800,
       G24801,G24802,G24803,G24804,G24805,G24806,G24807,G24808,G24809,G24810,G24811,G24812,G24813,G24814,G24815,G24816,G24817,G24818,G24819,G24820,
       G24821,G24822,G24823,G24824,G24825,G24826,G24827,G24828,G24829,G24830,G24831,G24832,G24833,G24834,G24835,G24836,G24837,G24838,G24839,G24840,
       G24841,G24842,G24843,G24844,G24845,G24846,G24847,G24848,G24849,G24850,G24851,G24852,G24853,G24854,G24855,G24856,G24857,G24858,G24859,G24860,
       G24861,G24862,G24863,G24864,G24865,G24866,G24867,G24868,G24869,G24870,G24871,G24872,G24873,G24874,G24875,G24876,G24877,G24878,G24879,G24880,
       G24881,G24882,G24883,G24884,G24885,G24886,G24887,G24888,G24889,G24890,G24891,G24892,G24893,G24894,G24895,G24896,G24897,G24898,G24899,G24900,
       G24901,G24902,G24903,G24904,G24905,G24906,G24907,G24908,G24909,G24910,G24911,G24912,G24913,G24914,G24915,G24916,G24917,G24918,G24919,G24920,
       G24921,G24922,G24923,G24924,G24925,G24926,G24927,G24928,G24929,G24930,G24931,G24932,G24933,G24934,G24935,G24936,G24937,G24938,G24939,G24940,
       G24941,G24942,G24943,G24944,G24945,G24946,G24947,G24948,G24949,G24950,G24951,G24952,G24953,G24954,G24955,G24956,G24957,G24958,G24959,G24960,
       G24961,G24962,G24963,G24964,G24965,G24966,G24967,G24968,G24969,G24970,G24971,G24972,G24973,G24974,G24975,G24976,G24977,G24978,G24979,G24980,
       G24981,G24982,G24983,G24984,G24985,G24986,G24987,G24988,G24989,G24990,G24991,G24992,G24993,G24994,G24995,G24996,G24997,G24998,G24999,G25000,
       G25001,G25002,G25003,G25004,G25005,G25006,G25007,G25008,G25009,G25010,G25011,G25012,G25013,G25014,G25015,G25016,G25017,G25018,G25019,G25020,
       G25021,G25022,G25023,G25024,G25025,G25026,G25027,G25028,G25029,G25030,G25031,G25032,G25033,G25034,G25035,G25036,G25037,G25038,G25039,G25040,
       G25041,G25042,G25043,G25044,G25045,G25046,G25047,G25048,G25049,G25050,G25051,G25052,G25053,G25054,G25055,G25056,G25057,G25058,G25059,G25060,
       G25061,G25062,G25063,G25064,G25065,G25066,G25067,G25068,G25069,G25070,G25071,G25072,G25073,G25074,G25075,G25076,G25077,G25078,G25079,G25080,
       G25081,G25082,G25083,G25084,G25085,G25086,G25087,G25088,G25089,G25090,G25091,G25092,G25093,G25094,G25095,G25096,G25097,G25098,G25099,G25100,
       G25101,G25102,G25103,G25104,G25105,G25106,G25107,G25108,G25109,G25110,G25111,G25112,G25113,G25114,G25115,G25116,G25117,G25118,G25119,G25120,
       G25121,G25122,G25123,G25124,G25125,G25126,G25127,G25128,G25129,G25130,G25131,G25132,G25133,G25134,G25135,G25136,G25137,G25138,G25139,G25140,
       G25141,G25142,G25143,G25144,G25145,G25146,G25147,G25148,G25149,G25150,G25151,G25152,G25153,G25154,G25155,G25156,G25157,G25158,G25159,G25160,
       G25161,G25162,G25163,G25164,G25165,G25166,G25167,G25168,G25169,G25170,G25171,G25172,G25173,G25174,G25175,G25176,G25177,G25178,G25179,G25180,
       G25181,G25182,G25183,G25184,G25185,G25186,G25187,G25188,G25189,G25190,G25191,G25192,G25193,G25194,G25195,G25196,G25197,G25198,G25199,G25200,
       G25201,G25202,G25203,G25204,G25205,G25206,G25207,G25208,G25209,G25210,G25211,G25212,G25213,G25214,G25215,G25216,G25217,G25218,G25219,G25220,
       G25221,G25222,G25223,G25224,G25225,G25226,G25227,G25228,G25229,G25230,G25231,G25232,G25233,G25234,G25235,G25236,G25237,G25238,G25239,G25240,
       G25241,G25242,G25243,G25244,G25245,G25246,G25247,G25248,G25249,G25250,G25251,G25252,G25253,G25254,G25255,G25256,G25257,G25258,G25259,G25260,
       G25261,G25262,G25263,G25264,G25265,G25266,G25267,G25268,G25269,G25270,G25271,G25272,G25273,G25274,G25275,G25276,G25277,G25278,G25279,G25280,
       G25281,G25282,G25283,G25284,G25285,G25286,G25287,G25288,G25289,G25290,G25291,G25292,G25293,G25294,G25295,G25296,G25297,G25298,G25299,G25300,
       G25301,G25302,G25303,G25304,G25305,G25306,G25307,G25308,G25309,G25310,G25311,G25312,G25313,G25314,G25315,G25316,G25317,G25318,G25319,G25320,
       G25321,G25322,G25323,G25324,G25325,G25326,G25327,G25328,G25329,G25330,G25331,G25332,G25333,G25334,G25335,G25336,G25337,G25338,G25339,G25340,
       G25341,G25342,G25343,G25344,G25345,G25346,G25347,G25348,G25349,G25350,G25351,G25352,G25353,G25354,G25355,G25356,G25357,G25358,G25359,G25360,
       G25361,G25362,G25363,G25364,G25365,G25366,G25367,G25368,G25369,G25370,G25371,G25372,G25373,G25374,G25375,G25376,G25377,G25378,G25379,G25380,
       G25381,G25382,G25383,G25384,G25385,G25386,G25387,G25388,G25389,G25390,G25391,G25392,G25393,G25394,G25395,G25396,G25397,G25398,G25399,G25400,
       G25401,G25402,G25403,G25404,G25405,G25406,G25407,G25408,G25409,G25410,G25411,G25412,G25413,G25414,G25415,G25416,G25417,G25418,G25419,G25420,
       G25421,G25422,G25423,G25424,G25425,G25426,G25427,G25428,G25429,G25430,G25431,G25432,G25433,G25434,G25435,G25436,G25437,G25438,G25439,G25440,
       G25441,G25442,G25443,G25444,G25445,G25446,G25447,G25448,G25449,G25450,G25451,G25452,G25453,G25454,G25455,G25456,G25457,G25458,G25459,G25460,
       G25461,G25462,G25463,G25464,G25465,G25466,G25467,G25468,G25469,G25470,G25471,G25472,G25473,G25474,G25475,G25476,G25477,G25478,G25479,G25480,
       G25481,G25482,G25483,G25484,G25485,G25486,G25487,G25488,G25489,G25490,G25491,G25492,G25493,G25494,G25495,G25496,G25497,G25498,G25499,G25500,
       G25501,G25502,G25503,G25504,G25505,G25506,G25507,G25508,G25509,G25510,G25511,G25512,G25513,G25514,G25515,G25516,G25517,G25518,G25519,G25520,
       G25521,G25522,G25523,G25524,G25525,G25526,G25527,G25528,G25529,G25530,G25531,G25532,G25533,G25534,G25535,G25536,G25537,G25538,G25539,G25540,
       G25541,G25542,G25543,G25544,G25545,G25546,G25547,G25548,G25549,G25550,G25551,G25552,G25553,G25554,G25555,G25556,G25557,G25558,G25559,G25560,
       G25561,G25562,G25563,G25564,G25565,G25566,G25567,G25568,G25569,G25570,G25571,G25572,G25573,G25574,G25575,G25576,G25577,G25578,G25579,G25580,
       G25581,G25582,G25583,G25584,G25585,G25586,G25587,G25588,G25589,G25590,G25591,G25592,G25593,G25594,G25595,G25596,G25597,G25598,G25599,G25600,
       G25601,G25602,G25603,G25604,G25605,G25606,G25607,G25608,G25609,G25610,G25611,G25612,G25613,G25614,G25615,G25616,G25617,G25618,G25619,G25620,
       G25621,G25622,G25623,G25624,G25625,G25626,G25627,G25628,G25629,G25630,G25631,G25632,G25633,G25634,G25635,G25636,G25637,G25638,G25639,G25640,
       G25641,G25642,G25643,G25644,G25645,G25646,G25647,G25648,G25649,G25650,G25651,G25652,G25653,G25654,G25655,G25656,G25657,G25658,G25659,G25660,
       G25661,G25662,G25663,G25664,G25665,G25666,G25667,G25668,G25669,G25670,G25671,G25672,G25673,G25674,G25675,G25676,G25677,G25678,G25679,G25680,
       G25681,G25682,G25683,G25684,G25685,G25686,G25687,G25688,G25689,G25690,G25691,G25692,G25693,G25694,G25695,G25696,G25697,G25698,G25699,G25700,
       G25701,G25702,G25703,G25704,G25705,G25706,G25707,G25708,G25709,G25710,G25711,G25712,G25713,G25714,G25715,G25716,G25717,G25718,G25719,G25720,
       G25721,G25722,G25723,G25724,G25725,G25726,G25727,G25728,G25729,G25730,G25731,G25732,G25733,G25734,G25735,G25736,G25737,G25738,G25739,G25740,
       G25741,G25742,G25743,G25744,G25745,G25746,G25747,G25748,G25749,G25750,G25751,G25752,G25753,G25754,G25755,G25756,G25757,G25758,G25759,G25760,
       G25761,G25762,G25763,G25764,G25765,G25766,G25767,G25768,G25769,G25770,G25771,G25772,G25773,G25774,G25775,G25776,G25777,G25778,G25779,G25780,
       G25781,G25782,G25783,G25784,G25785,G25786,G25787,G25788,G25789,G25790,G25791,G25792,G25793,G25794,G25795,G25796,G25797,G25798,G25799,G25800,
       G25801,G25802,G25803,G25804,G25805,G25806,G25807,G25808,G25809,G25810,G25811,G25812,G25813,G25814,G25815,G25816,G25817,G25818,G25819,G25820,
       G25821,G25822,G25823,G25824,G25825,G25826,G25827,G25828,G25829,G25830,G25831,G25832,G25833,G25834,G25835,G25836,G25837,G25838,G25839,G25840,
       G25841,G25842,G25843,G25844,G25845,G25846,G25847,G25848,G25849,G25850,G25851,G25852,G25853,G25854,G25855,G25856,G25857,G25858,G25859,G25860,
       G25861,G25862,G25863,G25864,G25865,G25866,G25867,G25868,G25869,G25870,G25871,G25872,G25873,G25874,G25875,G25876,G25877,G25878,G25879,G25880,
       G25881,G25882,G25883,G25884,G25885,G25886,G25887,G25888,G25889,G25890,G25891,G25892,G25893,G25894,G25895,G25896,G25897,G25898,G25899,G25900,
       G25901,G25902,G25903,G25904,G25905,G25906,G25907,G25908,G25909,G25910,G25911,G25912,G25913,G25914,G25915,G25916,G25917,G25918,G25919,G25920,
       G25921,G25922,G25923,G25924,G25925,G25926,G25927,G25928,G25929,G25930,G25931,G25932,G25933,G25934,G25935,G25936,G25937,G25938,G25939,G25940,
       G25941,G25942,G25943,G25944,G25945,G25946,G25947,G25948,G25949,G25950,G25951,G25952,G25953,G25954,G25955,G25956,G25957,G25958,G25959,G25960,
       G25961,G25962,G25963,G25964,G25965,G25966,G25967,G25968,G25969,G25970,G25971,G25972,G25973,G25974,G25975,G25976,G25977,G25978,G25979,G25980,
       G25981,G25982,G25983,G25984,G25985,G25986,G25987,G25988,G25989,G25990,G25991,G25992,G25993,G25994,G25995,G25996,G25997,G25998,G25999,G26000,
       G26001,G26002,G26003,G26004,G26005,G26006,G26007,G26008,G26009,G26010,G26011,G26012,G26013,G26014,G26015,G26016,G26017,G26018,G26019,G26020,
       G26021,G26022,G26023,G26024,G26025,G26026,G26027,G26028,G26029,G26030,G26031,G26032,G26033,G26034,G26035,G26036,G26037,G26038,G26039,G26040,
       G26041,G26042,G26043,G26044,G26045,G26046,G26047,G26048,G26049,G26050,G26051,G26052,G26053,G26054,G26055,G26056,G26057,G26058,G26059,G26060,
       G26061,G26062,G26063,G26064,G26065,G26066,G26067,G26068,G26069,G26070,G26071,G26072,G26073,G26074,G26075,G26076,G26077,G26078,G26079,G26080,
       G26081,G26082,G26083,G26084,G26085,G26086,G26087,G26088,G26089,G26090,G26091,G26092,G26093,G26094,G26095,G26096,G26097,G26098,G26099,G26100,
       G26101,G26102,G26103,G26104,G26105,G26106,G26107,G26108,G26109,G26110,G26111,G26112,G26113,G26114,G26115,G26116,G26117,G26118,G26119,G26120,
       G26121,G26122,G26123,G26124,G26125,G26126,G26127,G26128,G26129,G26130,G26131,G26132,G26133,G26134,G26135,G26136,G26137,G26138,G26139,G26140,
       G26141,G26142,G26143,G26144,G26145,G26146,G26147,G26148,G26149,G26150,G26151,G26152,G26153,G26154,G26155,G26156,G26157,G26158,G26159,G26160,
       G26161,G26162,G26163,G26164,G26165,G26166,G26167,G26168,G26169,G26170,G26171,G26172,G26173,G26174,G26175,G26176,G26177,G26178,G26179,G26180,
       G26181,G26182,G26183,G26184,G26185,G26186,G26187,G26188,G26189,G26190,G26191,G26192,G26193,G26194,G26195,G26196,G26197,G26198,G26199,G26200,
       G26201,G26202,G26203,G26204,G26205,G26206,G26207,G26208,G26209,G26210,G26211,G26212,G26213,G26214,G26215,G26216,G26217,G26218,G26219,G26220,
       G26221,G26222,G26223,G26224,G26225,G26226,G26227,G26228,G26229,G26230,G26231,G26232,G26233,G26234,G26235,G26236,G26237,G26238,G26239,G26240,
       G26241,G26242,G26243,G26244,G26245,G26246,G26247,G26248,G26249,G26250,G26251,G26252,G26253,G26254,G26255,G26256,G26257,G26258,G26259,G26260,
       G26261,G26262,G26263,G26264,G26265,G26266,G26267,G26268,G26269,G26270,G26271,G26272,G26273,G26274,G26275,G26276,G26277,G26278,G26279,G26280,
       G26281,G26282,G26283,G26284,G26285,G26286,G26287,G26288,G26289,G26290,G26291,G26292,G26293,G26294,G26295,G26296,G26297,G26298,G26299,G26300,
       G26301,G26302,G26303,G26304,G26305,G26306,G26307,G26308,G26309,G26310,G26311,G26312,G26313,G26314,G26315,G26316,G26317,G26318,G26319,G26320,
       G26321,G26322,G26323,G26324,G26325,G26326,G26327,G26328,G26329,G26330,G26331,G26332,G26333,G26334,G26335,G26336,G26337,G26338,G26339,G26340,
       G26341,G26342,G26343,G26344,G26345,G26346,G26347,G26348,G26349,G26350,G26351,G26352,G26353,G26354,G26355,G26356,G26357,G26358,G26359,G26360,
       G26361,G26362,G26363,G26364,G26365,G26366,G26367,G26368,G26369,G26370,G26371,G26372,G26373,G26374,G26375,G26376,G26377,G26378,G26379,G26380,
       G26381,G26382,G26383,G26384,G26385,G26386,G26387,G26388,G26389,G26390,G26391,G26392,G26393,G26394,G26395,G26396,G26397,G26398,G26399,G26400,
       G26401,G26402,G26403,G26404,G26405,G26406,G26407,G26408,G26409,G26410,G26411,G26412,G26413,G26414,G26415,G26416,G26417,G26418,G26419,G26420,
       G26421,G26422,G26423,G26424,G26425,G26426,G26427,G26428,G26429,G26430,G26431,G26432,G26433,G26434,G26435,G26436,G26437,G26438,G26439,G26440,
       G26441,G26442,G26443,G26444,G26445,G26446,G26447,G26448,G26449,G26450,G26451,G26452,G26453,G26454,G26455,G26456,G26457,G26458,G26459,G26460,
       G26461,G26462,G26463,G26464,G26465,G26466,G26467,G26468,G26469,G26470,G26471,G26472,G26473,G26474,G26475,G26476,G26477,G26478,G26479,G26480,
       G26481,G26482,G26483,G26484,G26485,G26486,G26487,G26488,G26489,G26490,G26491,G26492,G26493,G26494,G26495,G26496,G26497,G26498,G26499,G26500,
       G26501,G26502,G26503,G26504,G26505,G26506,G26507,G26508,G26509,G26510,G26511,G26512,G26513,G26514,G26515,G26516,G26517,G26518,G26519,G26520,
       G26521,G26522,G26523,G26524,G26525,G26526,G26527,G26528,G26529,G26530,G26531,G26532,G26533,G26534,G26535,G26536,G26537,G26538,G26539,G26540,
       G26541,G26542,G26543,G26544,G26545,G26546,G26547,G26548,G26549,G26550,G26551,G26552,G26553,G26554,G26555,G26556,G26557,G26558,G26559,G26560,
       G26561,G26562,G26563,G26564,G26565,G26566,G26567,G26568,G26569,G26570,G26571,G26572,G26573,G26574,G26575,G26576,G26577,G26578,G26579,G26580,
       G26581,G26582,G26583,G26584,G26585,G26586,G26587,G26588,G26589,G26590,G26591,G26592,G26593,G26594,G26595,G26596,G26597,G26598,G26599,G26600,
       G26601,G26602,G26603,G26604,G26605,G26606,G26607,G26608,G26609,G26610,G26611,G26612,G26613,G26614,G26615,G26616,G26617,G26618,G26619,G26620,
       G26621,G26622,G26623,G26624,G26625,G26626,G26627,G26628,G26629,G26630,G26631,G26632,G26633,G26634,G26635,G26636,G26637,G26638,G26639,G26640,
       G26641,G26642,G26643,G26644,G26645,G26646,G26647,G26648,G26649,G26650,G26651,G26652,G26653,G26654,G26655,G26656,G26657,G26658,G26659,G26660,
       G26661,G26662,G26663,G26664,G26665,G26666,G26667,G26668,G26669,G26670,G26671,G26672,G26673,G26674,G26675,G26676,G26677,G26678,G26679,G26680,
       G26681,G26682,G26683,G26684,G26685,G26686,G26687,G26688,G26689,G26690,G26691,G26692,G26693,G26694,G26695,G26696,G26697,G26698,G26699,G26700,
       G26701,G26702,G26703,G26704,G26705,G26706,G26707,G26708,G26709,G26710,G26711,G26712,G26713,G26714,G26715,G26716,G26717,G26718,G26719,G26720,
       G26721,G26722,G26723,G26724,G26725,G26726,G26727,G26728,G26729,G26730,G26731,G26732,G26733,G26734,G26735,G26736,G26737,G26738,G26739,G26740,
       G26741,G26742,G26743,G26744,G26745,G26746,G26747,G26748,G26749,G26750,G26751,G26752,G26753,G26754,G26755,G26756,G26757,G26758,G26759,G26760,
       G26761,G26762,G26763,G26764,G26765,G26766,G26767,G26768,G26769,G26770,G26771,G26772,G26773,G26774,G26775,G26776,G26777,G26778,G26779,G26780,
       G26781,G26782,G26783,G26784,G26785,G26786,G26787,G26788,G26789,G26790,G26791,G26792,G26793,G26794,G26795,G26796,G26797,G26798,G26799,G26800,
       G26801,G26802,G26803,G26804,G26805,G26806,G26807,G26808,G26809,G26810,G26811,G26812,G26813,G26814,G26815,G26816,G26817,G26818,G26819,G26820,
       G26821,G26822,G26823,G26824,G26825,G26826,G26827,G26828,G26829,G26830,G26831,G26832,G26833,G26834,G26835,G26836,G26837,G26838,G26839,G26840,
       G26841,G26842,G26843,G26844,G26845,G26846,G26847,G26848,G26849,G26850,G26851,G26852,G26853,G26854,G26855,G26856,G26857,G26858,G26859,G26860,
       G26861,G26862,G26863,G26864,G26865,G26866,G26867,G26868,G26869,G26870,G26871,G26872,G26873,G26874,G26875,G26876,G26877,G26878,G26879,G26880,
       G26881,G26882,G26883,G26884,G26885,G26886,G26887,G26888,G26889,G26890,G26891,G26892,G26893,G26894,G26895,G26896,G26897,G26898,G26899,G26900,
       G26901,G26902,G26903,G26904,G26905,G26906,G26907,G26908,G26909,G26910,G26911,G26912,G26913,G26914,G26915,G26916,G26917,G26918,G26919,G26920,
       G26921,G26922,G26923,G26924,G26925,G26926,G26927,G26928,G26929,G26930,G26931,G26932,G26933,G26934,G26935,G26936,G26937,G26938,G26939,G26940,
       G26941,G26942,G26943,G26944,G26945,G26946,G26947,G26948,G26949,G26950,G26951,G26952,G26953,G26954,G26955,G26956,G26957,G26958,G26959,G26960,
       G26961,G26962,G26963,G26964,G26965,G26966,G26967,G26968,G26969,G26970,G26971,G26972,G26973,G26974,G26975,G26976,G26977,G26978,G26979,G26980,
       G26981,G26982,G26983,G26984,G26985,G26986,G26987,G26988,G26989,G26990,G26991,G26992,G26993,G26994,G26995,G26996,G26997,G26998,G26999,G27000,
       G27001,G27002,G27003,G27004,G27005,G27006,G27007,G27008,G27009,G27010,G27011,G27012,G27013,G27014,G27015,G27016,G27017,G27018,G27019,G27020,
       G27021,G27022,G27023,G27024,G27025,G27026,G27027,G27028,G27029,G27030,G27031,G27032,G27033,G27034,G27035,G27036,G27037,G27038,G27039,G27040,
       G27041,G27042,G27043,G27044,G27045,G27046,G27047,G27048,G27049,G27050,G27051,G27052,G27053,G27054,G27055,G27056,G27057,G27058,G27059,G27060,
       G27061,G27062,G27063,G27064,G27065,G27066,G27067,G27068,G27069,G27070,G27071,G27072,G27073,G27074,G27075,G27076,G27077,G27078,G27079,G27080,
       G27081,G27082,G27083,G27084,G27085,G27086,G27087,G27088,G27089,G27090,G27091,G27092,G27093,G27094,G27095,G27096,G27097,G27098,G27099,G27100,
       G27101,G27102,G27103,G27104,G27105,G27106,G27107,G27108,G27109,G27110,G27111,G27112,G27113,G27114,G27115,G27116,G27117,G27118,G27119,G27120,
       G27121,G27122,G27123,G27124,G27125,G27126,G27127,G27128,G27129,G27130,G27131,G27132,G27133,G27134,G27135,G27136,G27137,G27138,G27139,G27140,
       G27141,G27142,G27143,G27144,G27145,G27146,G27147,G27148,G27149,G27150,G27151,G27152,G27153,G27154,G27155,G27156,G27157,G27158,G27159,G27160,
       G27161,G27162,G27163,G27164,G27165,G27166,G27167,G27168,G27169,G27170,G27171,G27172,G27173,G27174,G27175,G27176,G27177,G27178,G27179,G27180,
       G27181,G27182,G27183,G27184,G27185,G27186,G27187,G27188,G27189,G27190,G27191,G27192,G27193,G27194,G27195,G27196,G27197,G27198,G27199,G27200,
       G27201,G27202,G27203,G27204,G27205,G27206,G27207,G27208,G27209,G27210,G27211,G27212,G27213,G27214,G27215,G27216,G27217,G27218,G27219,G27220,
       G27221,G27222,G27223,G27224,G27225,G27226,G27227,G27228,G27229,G27230,G27231,G27232,G27233,G27234,G27235,G27236,G27237,G27238,G27239,G27240,
       G27241,G27242,G27243,G27244,G27245,G27246,G27247,G27248,G27249,G27250,G27251,G27252,G27253,G27254,G27255,G27256,G27257,G27258,G27259,G27260,
       G27261,G27262,G27263,G27264,G27265,G27266,G27267,G27268,G27269,G27270,G27271,G27272,G27273,G27274,G27275,G27276,G27277,G27278,G27279,G27280,
       G27281,G27282,G27283,G27284,G27285,G27286,G27287,G27288,G27289,G27290,G27291,G27292,G27293,G27294,G27295,G27296,G27297,G27298,G27299,G27300,
       G27301,G27302,G27303,G27304,G27305,G27306,G27307,G27308,G27309,G27310,G27311,G27312,G27313,G27314,G27315,G27316,G27317,G27318,G27319,G27320,
       G27321,G27322,G27323,G27324,G27325,G27326,G27327,G27328,G27329,G27330,G27331,G27332,G27333,G27334,G27335,G27336,G27337,G27338,G27339,G27340,
       G27341,G27342,G27343,G27344,G27345,G27346,G27347,G27348,G27349,G27350,G27351,G27352,G27353,G27354,G27355,G27356,G27357,G27358,G27359,G27360,
       G27361,G27362,G27363,G27364,G27365,G27366,G27367,G27368,G27369,G27370,G27371,G27372,G27373,G27374,G27375,G27376,G27377,G27378,G27379,G27380,
       G27381,G27382,G27383,G27384,G27385,G27386,G27387,G27388,G27389,G27390,G27391,G27392,G27393,G27394,G27395,G27396,G27397,G27398,G27399,G27400,
       G27401,G27402,G27403,G27404,G27405,G27406,G27407,G27408,G27409,G27410,G27411,G27412,G27413,G27414,G27415,G27416,G27417,G27418,G27419,G27420,
       G27421,G27422,G27423,G27424,G27425,G27426,G27427,G27428,G27429,G27430,G27431,G27432,G27433,G27434,G27435,G27436,G27437,G27438,G27439,G27440,
       G27441,G27442,G27443,G27444,G27445,G27446,G27447,G27448,G27449,G27450,G27451,G27452,G27453,G27454,G27455,G27456,G27457,G27458,G27459,G27460,
       G27461,G27462,G27463,G27464,G27465,G27466,G27467,G27468,G27469,G27470,G27471,G27472,G27473,G27474,G27475,G27476,G27477,G27478,G27479,G27480,
       G27481,G27482,G27483,G27484,G27485,G27486,G27487,G27488,G27489,G27490,G27491,G27492,G27493,G27494,G27495,G27496,G27497,G27498,G27499,G27500,
       G27501,G27502,G27503,G27504,G27505,G27506,G27507,G27508,G27509,G27510,G27511,G27512,G27513,G27514,G27515,G27516,G27517,G27518,G27519,G27520,
       G27521,G27522,G27523,G27524,G27525,G27526,G27527,G27528,G27529,G27530,G27531,G27532,G27533,G27534,G27535,G27536,G27537,G27538,G27539,G27540,
       G27541,G27542,G27543,G27544,G27545,G27546,G27547,G27548,G27549,G27550,G27551,G27552,G27553,G27554,G27555,G27556,G27557,G27558,G27559,G27560,
       G27561,G27562,G27563,G27564,G27565,G27566,G27567,G27568,G27569,G27570,G27571,G27572,G27573,G27574,G27575,G27576,G27577,G27578,G27579,G27580,
       G27581,G27582,G27583,G27584,G27585,G27586,G27587,G27588,G27589,G27590,G27591,G27592,G27593,G27594,G27595,G27596,G27597,G27598,G27599,G27600,
       G27601,G27602,G27603,G27604,G27605,G27606,G27607,G27608,G27609,G27610,G27611,G27612,G27613,G27614,G27615,G27616,G27617,G27618,G27619,G27620,
       G27621,G27622,G27623,G27624,G27625,G27626,G27627,G27628,G27629,G27630,G27631,G27632,G27633,G27634,G27635,G27636,G27637,G27638,G27639,G27640,
       G27641,G27642,G27643,G27644,G27645,G27646,G27647,G27648,G27649,G27650,G27651,G27652,G27653,G27654,G27655,G27656,G27657,G27658,G27659,G27660,
       G27661,G27662,G27663,G27664,G27665,G27666,G27667,G27668,G27669,G27670,G27671,G27672,G27673,G27674,G27675,G27676,G27677,G27678,G27679,G27680,
       G27681,G27682,G27683,G27684,G27685,G27686,G27687,G27688,G27689,G27690,G27691,G27692,G27693,G27694,G27695,G27696,G27697,G27698,G27699,G27700,
       G27701,G27702,G27703,G27704,G27705,G27706,G27707,G27708,G27709,G27710,G27711,G27712,G27713,G27714,G27715,G27716,G27717,G27718,G27719,G27720,
       G27721,G27722,G27723,G27724,G27725,G27726,G27727,G27728,G27729,G27730,G27731,G27732,G27733,G27734,G27735,G27736,G27737,G27738,G27739,G27740,
       G27741,G27742,G27743,G27744,G27745,G27746,G27747,G27748,G27749,G27750,G27751,G27752,G27753,G27754,G27755,G27756,G27757,G27758,G27759,G27760,
       G27761,G27762,G27763,G27764,G27765,G27766,G27767,G27768,G27769,G27770,G27771,G27772,G27773,G27774,G27775,G27776,G27777,G27778,G27779,G27780,
       G27781,G27782,G27783,G27784,G27785,G27786,G27787,G27788,G27789,G27790,G27791,G27792,G27793,G27794,G27795,G27796,G27797,G27798,G27799,G27800,
       G27801,G27802,G27803,G27804,G27805,G27806,G27807,G27808,G27809,G27810,G27811,G27812,G27813,G27814,G27815,G27816,G27817,G27818,G27819,G27820,
       G27821,G27822,G27823,G27824,G27825,G27826,G27827,G27828,G27829,G27830,G27831,G27832,G27833,G27834,G27835,G27836,G27837,G27838,G27839,G27840,
       G27841,G27842,G27843,G27844,G27845,G27846,G27847,G27848,G27849,G27850,G27851,G27852,G27853,G27854,G27855,G27856,G27857,G27858,G27859,G27860,
       G27861,G27862,G27863,G27864,G27865,G27866,G27867,G27868,G27869,G27870,G27871,G27872,G27873,G27874,G27875,G27876,G27877,G27878,G27879,G27880,
       G27881,G27882,G27883,G27884,G27885,G27886,G27887,G27888,G27889,G27890,G27891,G27892,G27893,G27894,G27895,G27896,G27897,G27898,G27899,G27900,
       G27901,G27902,G27903,G27904,G27905,G27906,G27907,G27908,G27909,G27910,G27911,G27912,G27913,G27914,G27915,G27916,G27917,G27918,G27919,G27920,
       G27921,G27922,G27923,G27924,G27925,G27926,G27927,G27928,G27929,G27930,G27931,G27932,G27933,G27934,G27935,G27936,G27937,G27938,G27939,G27940,
       G27941,G27942,G27943,G27944,G27945,G27946,G27947,G27948,G27949,G27950,G27951,G27952,G27953,G27954,G27955,G27956,G27957,G27958,G27959,G27960,
       G27961,G27962,G27963,G27964,G27965,G27966,G27967,G27968,G27969,G27970,G27971,G27972,G27973,G27974,G27975,G27976,G27977,G27978,G27979,G27980,
       G27981,G27982,G27983,G27984,G27985,G27986,G27987,G27988,G27989,G27990,G27991,G27992,G27993,G27994,G27995,G27996,G27997,G27998,G27999,G28000,
       G28001,G28002,G28003,G28004,G28005,G28006,G28007,G28008,G28009,G28010,G28011,G28012,G28013,G28014,G28015,G28016,G28017,G28018,G28019,G28020,
       G28021,G28022,G28023,G28024,G28025,G28026,G28027,G28028,G28029,G28030,G28031,G28032,G28033,G28034,G28035,G28036,G28037,G28038,G28039,G28040,
       G28041,G28042,G28043,G28044,G28045,G28046,G28047,G28048,G28049,G28050,G28051,G28052,G28053,G28054,G28055,G28056,G28057,G28058,G28059,G28060,
       G28061,G28062,G28063,G28064,G28065,G28066,G28067,G28068,G28069,G28070,G28071,G28072,G28073,G28074,G28075,G28076,G28077,G28078,G28079,G28080,
       G28081,G28082,G28083,G28084,G28085,G28086,G28087,G28088,G28089,G28090,G28091,G28092,G28093,G28094,G28095,G28096,G28097,G28098,G28099,G28100,
       G28101,G28102,G28103,G28104,G28105,G28106,G28107,G28108,G28109,G28110,G28111,G28112,G28113,G28114,G28115,G28116,G28117,G28118,G28119,G28120,
       G28121,G28122,G28123,G28124,G28125,G28126,G28127,G28128,G28129,G28130,G28131,G28132,G28133,G28134,G28135,G28136,G28137,G28138,G28139,G28140,
       G28141,G28142,G28143,G28144,G28145,G28146,G28147,G28148,G28149,G28150,G28151,G28152,G28153,G28154,G28155,G28156,G28157,G28158,G28159,G28160,
       G28161,G28162,G28163,G28164,G28165,G28166,G28167,G28168,G28169,G28170,G28171,G28172,G28173,G28174,G28175,G28176,G28177,G28178,G28179,G28180,
       G28181,G28182,G28183,G28184,G28185,G28186,G28187,G28188,G28189,G28190,G28191,G28192,G28193,G28194,G28195,G28196,G28197,G28198,G28199,G28200,
       G28201,G28202,G28203,G28204,G28205,G28206,G28207,G28208,G28209,G28210,G28211,G28212,G28213,G28214,G28215,G28216,G28217,G28218,G28219,G28220,
       G28221,G28222,G28223,G28224,G28225,G28226,G28227,G28228,G28229,G28230,G28231,G28232,G28233,G28234,G28235,G28236,G28237,G28238,G28239,G28240,
       G28241,G28242,G28243,G28244,G28245,G28246,G28247,G28248,G28249,G28250,G28251,G28252,G28253,G28254,G28255,G28256,G28257,G28258,G28259,G28260,
       G28261,G28262,G28263,G28264,G28265,G28266,G28267,G28268,G28269,G28270,G28271,G28272,G28273,G28274,G28275,G28276,G28277,G28278,G28279,G28280,
       G28281,G28282,G28283,G28284,G28285,G28286,G28287,G28288,G28289,G28290,G28291,G28292,G28293,G28294,G28295,G28296,G28297,G28298,G28299,G28300,
       G28301,G28302,G28303,G28304,G28305,G28306,G28307,G28308,G28309,G28310,G28311,G28312,G28313,G28314,G28315,G28316,G28317,G28318,G28319,G28320,
       G28321,G28322,G28323,G28324,G28325,G28326,G28327,G28328,G28329,G28330,G28331,G28332,G28333,G28334,G28335,G28336,G28337,G28338,G28339,G28340,
       G28341,G28342,G28343,G28344,G28345,G28346,G28347,G28348,G28349,G28350,G28351,G28352,G28353,G28354,G28355,G28356,G28357,G28358,G28359,G28360,
       G28361,G28362,G28363,G28364,G28365,G28366,G28367,G28368,G28369,G28370,G28371,G28372,G28373,G28374,G28375,G28376,G28377,G28378,G28379,G28380,
       G28381,G28382,G28383,G28384,G28385,G28386,G28387,G28388,G28389,G28390,G28391,G28392,G28393,G28394,G28395,G28396,G28397,G28398,G28399,G28400,
       G28401,G28402,G28403,G28404,G28405,G28406,G28407,G28408,G28409,G28410,G28411,G28412,G28413,G28414,G28415,G28416,G28417,G28418,G28419,G28420,
       G28421,G28422,G28423,G28424,G28425,G28426,G28427,G28428,G28429,G28430,G28431,G28432,G28433,G28434,G28435,G28436,G28437,G28438,G28439,G28440,
       G28441,G28442,G28443,G28444,G28445,G28446,G28447,G28448,G28449,G28450,G28451,G28452,G28453,G28454,G28455,G28456,G28457,G28458,G28459,G28460,
       G28461,G28462,G28463,G28464,G28465,G28466,G28467,G28468,G28469,G28470,G28471,G28472,G28473,G28474,G28475,G28476,G28477,G28478,G28479,G28480,
       G28481,G28482,G28483,G28484,G28485,G28486,G28487,G28488,G28489,G28490,G28491,G28492,G28493,G28494,G28495,G28496,G28497,G28498,G28499,G28500,
       G28501,G28502,G28503,G28504,G28505,G28506,G28507,G28508,G28509,G28510,G28511,G28512,G28513,G28514,G28515,G28516,G28517,G28518,G28519,G28520,
       G28521,G28522,G28523,G28524,G28525,G28526,G28527,G28528,G28529,G28530,G28531,G28532,G28533,G28534,G28535,G28536,G28537,G28538,G28539,G28540,
       G28541,G28542,G28543,G28544,G28545,G28546,G28547,G28548,G28549,G28550,G28551,G28552,G28553,G28554,G28555,G28556,G28557,G28558,G28559,G28560,
       G28561,G28562,G28563,G28564,G28565,G28566,G28567,G28568,G28569,G28570,G28571,G28572,G28573,G28574,G28575,G28576,G28577,G28578,G28579,G28580,
       G28581,G28582,G28583,G28584,G28585,G28586,G28587,G28588,G28589,G28590,G28591,G28592,G28593,G28594,G28595,G28596,G28597,G28598,G28599,G28600,
       G28601,G28602,G28603,G28604,G28605,G28606,G28607,G28608,G28609,G28610,G28611,G28612,G28613,G28614,G28615,G28616,G28617,G28618,G28619,G28620,
       G28621,G28622,G28623,G28624,G28625,G28626,G28627,G28628,G28629,G28630,G28631,G28632,G28633,G28634,G28635,G28636,G28637,G28638,G28639,G28640,
       G28641,G28642,G28643,G28644,G28645,G28646,G28647,G28648,G28649,G28650,G28651,G28652,G28653,G28654,G28655,G28656,G28657,G28658,G28659,G28660,
       G28661,G28662,G28663,G28664,G28665,G28666,G28667,G28668,G28669,G28670,G28671,G28672,G28673,G28674,G28675,G28676,G28677,G28678,G28679,G28680,
       G28681,G28682,G28683,G28684,G28685,G28686,G28687,G28688,G28689,G28690,G28691,G28692,G28693,G28694,G28695,G28696,G28697,G28698,G28699,G28700,
       G28701,G28702,G28703,G28704,G28705,G28706,G28707,G28708,G28709,G28710,G28711,G28712,G28713,G28714,G28715,G28716,G28717,G28718,G28719,G28720,
       G28721,G28722,G28723,G28724,G28725,G28726,G28727,G28728,G28729,G28730,G28731,G28732,G28733,G28734,G28735,G28736,G28737,G28738,G28739,G28740,
       G28741,G28742,G28743,G28744,G28745,G28746,G28747,G28748,G28749,G28750,G28751,G28752,G28753,G28754,G28755,G28756,G28757,G28758,G28759,G28760,
       G28761,G28762,G28763,G28764,G28765,G28766,G28767,G28768,G28769,G28770,G28771,G28772,G28773,G28774,G28775,G28776,G28777,G28778,G28779,G28780,
       G28781,G28782,G28783,G28784,G28785,G28786,G28787,G28788,G28789,G28790,G28791,G28792,G28793,G28794,G28795,G28796,G28797,G28798,G28799,G28800,
       G28801,G28802,G28803,G28804,G28805,G28806,G28807,G28808,G28809,G28810,G28811,G28812,G28813,G28814,G28815,G28816,G28817,G28818,G28819,G28820,
       G28821,G28822,G28823,G28824,G28825,G28826,G28827,G28828,G28829,G28830,G28831,G28832,G28833,G28834,G28835,G28836,G28837,G28838,G28839,G28840,
       G28841,G28842,G28843,G28844,G28845,G28846,G28847,G28848,G28849,G28850,G28851,G28852,G28853,G28854,G28855,G28856,G28857,G28858,G28859,G28860,
       G28861,G28862,G28863,G28864,G28865,G28866,G28867,G28868,G28869,G28870,G28871,G28872,G28873,G28874,G28875,G28876,G28877,G28878,G28879,G28880,
       G28881,G28882,G28883,G28884,G28885,G28886,G28887,G28888,G28889,G28890,G28891,G28892,G28893,G28894,G28895,G28896,G28897,G28898,G28899,G28900,
       G28901,G28902,G28903,G28904,G28905,G28906,G28907,G28908,G28909,G28910,G28911,G28912,G28913,G28914,G28915,G28916,G28917,G28918,G28919,G28920,
       G28921,G28922,G28923,G28924,G28925,G28926,G28927,G28928,G28929,G28930,G28931,G28932,G28933,G28934,G28935,G28936,G28937,G28938,G28939,G28940,
       G28941,G28942,G28943,G28944,G28945,G28946,G28947,G28948,G28949,G28950,G28951,G28952,G28953,G28954,G28955,G28956,G28957,G28958,G28959,G28960,
       G28961,G28962,G28963,G28964,G28965,G28966,G28967,G28968,G28969,G28970,G28971,G28972,G28973,G28974,G28975,G28976,G28977,G28978,G28979,G28980,
       G28981,G28982,G28983,G28984,G28985,G28986,G28987,G28988,G28989,G28990,G28991,G28992,G28993,G28994,G28995,G28996,G28997,G28998,G28999,G29000,
       G29001,G29002,G29003,G29004,G29005,G29006,G29007,G29008,G29009,G29010,G29011,G29012,G29013,G29014,G29015,G29016,G29017,G29018,G29019,G29020,
       G29021,G29022,G29023,G29024,G29025,G29026,G29027,G29028,G29029,G29030,G29031,G29032,G29033,G29034,G29035,G29036,G29037,G29038,G29039,G29040,
       G29041,G29042,G29043,G29044,G29045,G29046,G29047,G29048,G29049,G29050,G29051,G29052,G29053,G29054,G29055,G29056,G29057,G29058,G29059,G29060,
       G29061,G29062,G29063,G29064,G29065,G29066,G29067,G29068,G29069,G29070,G29071,G29072,G29073,G29074,G29075,G29076,G29077,G29078,G29079,G29080,
       G29081,G29082,G29083,G29084,G29085,G29086,G29087,G29088,G29089,G29090,G29091,G29092,G29093,G29094,G29095,G29096,G29097,G29098,G29099,G29100,
       G29101,G29102,G29103,G29104,G29105,G29106,G29107,G29108,G29109,G29110,G29111,G29112,G29113,G29114,G29115,G29116,G29117,G29118,G29119,G29120,
       G29121,G29122,G29123,G29124,G29125,G29126,G29127,G29128,G29129,G29130,G29131,G29132,G29133,G29134,G29135,G29136,G29137,G29138,G29139,G29140,
       G29141,G29142,G29143,G29144,G29145,G29146,G29147,G29148,G29149,G29150,G29151,G29152,G29153,G29154,G29155,G29156,G29157,G29158,G29159,G29160,
       G29161,G29162,G29163,G29164,G29165,G29166,G29167,G29168,G29169,G29170,G29171,G29172,G29173,G29174,G29175,G29176,G29177,G29178,G29179,G29180,
       G29181,G29182,G29183,G29184,G29185,G29186,G29187,G29188,G29189,G29190,G29191,G29192,G29193,G29194,G29195,G29196,G29197,G29198,G29199,G29200,
       G29201,G29202,G29203,G29204,G29205,G29206,G29207,G29208,G29209,G29210,G29211,G29212,G29213,G29214,G29215,G29216,G29217,G29218,G29219,G29220,
       G29221,G29222,G29223,G29224,G29225,G29226,G29227,G29228,G29229,G29230,G29231,G29232,G29233,G29234,G29235,G29236,G29237,G29238,G29239,G29240,
       G29241,G29242,G29243,G29244,G29245,G29246,G29247,G29248,G29249,G29250,G29251,G29252,G29253,G29254,G29255,G29256,G29257,G29258,G29259,G29260,
       G29261,G29262,G29263,G29264,G29265,G29266,G29267,G29268,G29269,G29270,G29271,G29272,G29273,G29274,G29275,G29276,G29277,G29278,G29279,G29280,
       G29281,G29282,G29283,G29284,G29285,G29286,G29287,G29288,G29289,G29290,G29291,G29292,G29293,G29294,G29295,G29296,G29297,G29298,G29299,G29300,
       G29301,G29302,G29303,G29304,G29305,G29306,G29307,G29308,G29309,G29310,G29311,G29312,G29313,G29314,G29315,G29316,G29317,G29318,G29319,G29320,
       G29321,G29322,G29323,G29324,G29325,G29326,G29327,G29328,G29329,G29330,G29331,G29332,G29333,G29334,G29335,G29336,G29337,G29338,G29339,G29340,
       G29341,G29342,G29343,G29344,G29345,G29346,G29347,G29348,G29349,G29350,G29351,G29352,G29353,G29354,G29355,G29356,G29357,G29358,G29359,G29360,
       G29361,G29362,G29363,G29364,G29365,G29366,G29367,G29368,G29369,G29370,G29371,G29372,G29373,G29374,G29375,G29376,G29377,G29378,G29379,G29380,
       G29381,G29382,G29383,G29384,G29385,G29386,G29387,G29388,G29389,G29390,G29391,G29392,G29393,G29394,G29395,G29396,G29397,G29398,G29399,G29400,
       G29401,G29402,G29403,G29404,G29405,G29406,G29407,G29408,G29409,G29410,G29411,G29412,G29413,G29414,G29415,G29416,G29417,G29418,G29419,G29420,
       G29421,G29422,G29423,G29424,G29425,G29426,G29427,G29428,G29429,G29430,G29431,G29432,G29433,G29434,G29435,G29436,G29437,G29438,G29439,G29440,
       G29441,G29442,G29443,G29444,G29445,G29446,G29447,G29448,G29449,G29450,G29451,G29452,G29453,G29454,G29455,G29456,G29457,G29458,G29459,G29460,
       G29461,G29462,G29463,G29464,G29465,G29466,G29467,G29468,G29469,G29470,G29471,G29472,G29473,G29474,G29475,G29476,G29477,G29478,G29479,G29480,
       G29481,G29482,G29483,G29484,G29485,G29486,G29487,G29488,G29489,G29490,G29491,G29492,G29493,G29494,G29495,G29496,G29497,G29498,G29499,G29500,
       G29501,G29502,G29503,G29504,G29505,G29506,G29507,G29508,G29509,G29510,G29511,G29512,G29513,G29514,G29515,G29516,G29517,G29518,G29519,G29520,
       G29521,G29522,G29523,G29524,G29525,G29526,G29527,G29528,G29529,G29530,G29531,G29532,G29533,G29534,G29535,G29536,G29537,G29538,G29539,G29540,
       G29541,G29542,G29543,G29544,G29545,G29546,G29547,G29548,G29549,G29550,G29551,G29552,G29553,G29554,G29555,G29556,G29557,G29558,G29559,G29560,
       G29561,G29562,G29563,G29564,G29565,G29566,G29567,G29568,G29569,G29570,G29571,G29572,G29573,G29574,G29575,G29576,G29577,G29578,G29579,G29580,
       G29581,G29582,G29583,G29584,G29585,G29586,G29587,G29588,G29589,G29590,G29591,G29592,G29593,G29594,G29595,G29596,G29597,G29598,G29599,G29600,
       G29601,G29602,G29603,G29604,G29605,G29606,G29607,G29608,G29609,G29610,G29611,G29612,G29613,G29614,G29615,G29616,G29617,G29618,G29619,G29620,
       G29621,G29622,G29623,G29624,G29625,G29626,G29627,G29628,G29629,G29630,G29631,G29632,G29633,G29634,G29635,G29636,G29637,G29638,G29639,G29640,
       G29641,G29642,G29643,G29644,G29645,G29646,G29647,G29648,G29649,G29650,G29651,G29652,G29653,G29654,G29655,G29656,G29657,G29658,G29659,G29660,
       G29661,G29662,G29663,G29664,G29665,G29666,G29667,G29668,G29669,G29670,G29671,G29672,G29673,G29674,G29675,G29676,G29677,G29678,G29679,G29680,
       G29681,G29682,G29683,G29684,G29685,G29686,G29687,G29688,G29689,G29690,G29691,G29692,G29693,G29694,G29695,G29696,G29697,G29698,G29699,G29700,
       G29701,G29702,G29703,G29704,G29705,G29706,G29707,G29708,G29709,G29710,G29711,G29712,G29713,G29714,G29715,G29716,G29717,G29718,G29719,G29720,
       G29721,G29722,G29723,G29724,G29725,G29726,G29727,G29728,G29729,G29730,G29731,G29732,G29733,G29734,G29735,G29736,G29737,G29738,G29739,G29740,
       G29741,G29742,G29743,G29744,G29745,G29746,G29747,G29748,G29749,G29750,G29751,G29752,G29753,G29754,G29755,G29756,G29757,G29758,G29759,G29760,
       G29761,G29762,G29763,G29764,G29765,G29766,G29767,G29768,G29769,G29770,G29771,G29772,G29773,G29774,G29775,G29776,G29777,G29778,G29779,G29780,
       G29781,G29782,G29783,G29784,G29785,G29786,G29787,G29788,G29789,G29790,G29791,G29792,G29793,G29794,G29795,G29796,G29797,G29798,G29799,G29800,
       G29801,G29802,G29803,G29804,G29805,G29806,G29807,G29808,G29809,G29810,G29811,G29812,G29813,G29814,G29815,G29816,G29817,G29818,G29819,G29820,
       G29821,G29822,G29823,G29824,G29825,G29826,G29827,G29828,G29829,G29830,G29831,G29832,G29833,G29834,G29835,G29836,G29837,G29838,G29839,G29840,
       G29841,G29842,G29843,G29844,G29845,G29846,G29847,G29848,G29849,G29850,G29851,G29852,G29853,G29854,G29855,G29856,G29857,G29858,G29859,G29860,
       G29861,G29862,G29863,G29864,G29865,G29866,G29867,G29868,G29869,G29870,G29871,G29872,G29873,G29874,G29875,G29876,G29877,G29878,G29879,G29880,
       G29881,G29882,G29883,G29884,G29885,G29886,G29887,G29888,G29889,G29890,G29891,G29892,G29893,G29894,G29895,G29896,G29897,G29898,G29899,G29900,
       G29901,G29902,G29903,G29904,G29905,G29906,G29907,G29908,G29909,G29910,G29911,G29912,G29913,G29914,G29915,G29916,G29917,G29918,G29919,G29920,
       G29921,G29922,G29923,G29924,G29925,G29926,G29927,G29928,G29929,G29930,G29931,G29932,G29933,G29934,G29935,G29936,G29937,G29938,G29939,G29940,
       G29941,G29942,G29943,G29944,G29945,G29946,G29947,G29948,G29949,G29950,G29951,G29952,G29953,G29954,G29955,G29956,G29957,G29958,G29959,G29960,
       G29961,G29962,G29963,G29964,G29965,G29966,G29967,G29968,G29969,G29970,G29971,G29972,G29973,G29974,G29975,G29976,G29977,G29978,G29979,G29980,
       G29981,G29982,G29983,G29984,G29985,G29986,G29987,G29988,G29989,G29990,G29991,G29992,G29993,G29994,G29995,G29996,G29997,G29998,G29999,G30000,
       G30001,G30002,G30003,G30004,G30005,G30006,G30007,G30008,G30009,G30010,G30011,G30012,G30013,G30014,G30015,G30016,G30017,G30018,G30019,G30020,
       G30021,G30022,G30023,G30024,G30025,G30026,G30027,G30028,G30029,G30030,G30031,G30032,G30033,G30034,G30035,G30036,G30037,G30038,G30039,G30040,
       G30041,G30042,G30043,G30044,G30045,G30046,G30047,G30048,G30049,G30050,G30051,G30052,G30053,G30054,G30055,G30056,G30057,G30058,G30059,G30060,
       G30061,G30062,G30063,G30064,G30065,G30066,G30067,G30068,G30069,G30070,G30071,G30072,G30073,G30074,G30075,G30076,G30077,G30078,G30079,G30080,
       G30081,G30082,G30083,G30084,G30085,G30086,G30087,G30088,G30089,G30090,G30091,G30092,G30093,G30094,G30095,G30096,G30097,G30098,G30099,G30100,
       G30101,G30102,G30103,G30104,G30105,G30106,G30107,G30108,G30109,G30110,G30111,G30112,G30113,G30114,G30115,G30116,G30117,G30118,G30119,G30120,
       G30121,G30122,G30123,G30124,G30125,G30126,G30127,G30128,G30129,G30130,G30131,G30132,G30133,G30134,G30135,G30136,G30137,G30138,G30139,G30140,
       G30141,G30142,G30143,G30144,G30145,G30146,G30147,G30148,G30149,G30150,G30151,G30152,G30153,G30154,G30155,G30156,G30157,G30158,G30159,G30160,
       G30161,G30162,G30163,G30164,G30165,G30166,G30167,G30168,G30169,G30170,G30171,G30172,G30173,G30174,G30175,G30176,G30177,G30178,G30179,G30180,
       G30181,G30182,G30183,G30184,G30185,G30186,G30187,G30188,G30189,G30190,G30191,G30192,G30193,G30194,G30195,G30196,G30197,G30198,G30199,G30200,
       G30201,G30202,G30203,G30204,G30205,G30206,G30207,G30208,G30209,G30210,G30211,G30212,G30213,G30214,G30215,G30216,G30217,G30218,G30219,G30220,
       G30221,G30222,G30223,G30224,G30225,G30226,G30227,G30228,G30229,G30230,G30231,G30232,G30233,G30234,G30235,G30236,G30237,G30238,G30239,G30240,
       G30241,G30242,G30243,G30244,G30245,G30246,G30247,G30248,G30249,G30250,G30251,G30252,G30253,G30254,G30255,G30256,G30257,G30258,G30259,G30260,
       G30261,G30262,G30263,G30264,G30265,G30266,G30267,G30268,G30269,G30270,G30271,G30272,G30273,G30274,G30275,G30276,G30277,G30278,G30279,G30280,
       G30281,G30282,G30283,G30284,G30285,G30286,G30287,G30288,G30289,G30290,G30291,G30292,G30293,G30294,G30295,G30296,G30297,G30298,G30299,G30300,
       G30301,G30302,G30303,G30304,G30305,G30306,G30307,G30308,G30309,G30310,G30311,G30312,G30313,G30314,G30315,G30316,G30317,G30318,G30319,G30320,
       G30321,G30322,G30323,G30324,G30325,G30326,G30327,G30328,G30329,G30330,G30331,G30332,G30333,G30334,G30335,G30336,G30337,G30338,G30339,G30340,
       G30341,G30342,G30343,G30344,G30345,G30346,G30347,G30348,G30349,G30350,G30351,G30352,G30353,G30354,G30355,G30356,G30357,G30358,G30359,G30360,
       G30361,G30362,G30363,G30364,G30365,G30366,G30367,G30368,G30369,G30370,G30371,G30372,G30373,G30374,G30375,G30376,G30377,G30378,G30379,G30380,
       G30381,G30382,G30383,G30384,G30385,G30386,G30387,G30388,G30389,G30390,G30391,G30392,G30393,G30394,G30395,G30396,G30397,G30398,G30399,G30400,
       G30401,G30402,G30403,G30404,G30405,G30406,G30407,G30408,G30409,G30410,G30411,G30412,G30413,G30414,G30415,G30416,G30417,G30418,G30419,G30420,
       G30421,G30422,G30423,G30424,G30425,G30426,G30427,G30428,G30429,G30430,G30431,G30432,G30433,G30434,G30435,G30436,G30437,G30438,G30439,G30440,
       G30441,G30442,G30443,G30444,G30445,G30446,G30447,G30448,G30449,G30450,G30451,G30452,G30453,G30454,G30455,G30456,G30457,G30458,G30459,G30460,
       G30461,G30462,G30463,G30464,G30465,G30466,G30467,G30468,G30469,G30470,G30471,G30472,G30473,G30474,G30475,G30476,G30477,G30478,G30479,G30480,
       G30481,G30482,G30483,G30484,G30485,G30486,G30487,G30488,G30489,G30490,G30491,G30492,G30493,G30494,G30495,G30496,G30497,G30498,G30499,G30500,
       G30501,G30502,G30503,G30504,G30505,G30506,G30507,G30508,G30509,G30510,G30511,G30512,G30513,G30514,G30515,G30516,G30517,G30518,G30519,G30520,
       G30521,G30522,G30523,G30524,G30525,G30526,G30527,G30528,G30529,G30530,G30531,G30532,G30533,G30534,G30535,G30536,G30537,G30538,G30539,G30540,
       G30541,G30542,G30543,G30544,G30545,G30546,G30547,G30548,G30549,G30550,G30551,G30552,G30553,G30554,G30555,G30556,G30557,G30558,G30559,G30560,
       G30561,G30562,G30563,G30564,G30565,G30566,G30567,G30568,G30569,G30570,G30571,G30572,G30573,G30574,G30575,G30576,G30577,G30578,G30579,G30580,
       G30581,G30582,G30583,G30584,G30585,G30586,G30587,G30588,G30589,G30590,G30591,G30592,G30593,G30594,G30595,G30596,G30597,G30598,G30599,G30600,
       G30601,G30602,G30603,G30604,G30605,G30606,G30607,G30608,G30609,G30610,G30611,G30612,G30613,G30614,G30615,G30616,G30617,G30618,G30619,G30620,
       G30621,G30622,G30623,G30624,G30625,G30626,G30627,G30628,G30629,G30630,G30631,G30632,G30633,G30634,G30635,G30636,G30637,G30638,G30639,G30640,
       G30641,G30642,G30643,G30644,G30645,G30646,G30647,G30648,G30649,G30650,G30651,G30652,G30653,G30654,G30655,G30656,G30657,G30658,G30659,G30660,
       G30661,G30662,G30663,G30664,G30665,G30666,G30667,G30668,G30669,G30670,G30671,G30672,G30673,G30674,G30675,G30676,G30677,G30678,G30679,G30680,
       G30681,G30682,G30683,G30684,G30685,G30686,G30687,G30688,G30689,G30690,G30691,G30692,G30693,G30694,G30695,G30696,G30697,G30698,G30699,G30700,
       G30701,G30702,G30703,G30704,G30705,G30706,G30707,G30708,G30709,G30710,G30711,G30712,G30713,G30714,G30715,G30716,G30717,G30718,G30719,G30720,
       G30721,G30722,G30723,G30724,G30725,G30726,G30727,G30728,G30729,G30730,G30731,G30732,G30733,G30734,G30735,G30736,G30737,G30738,G30739,G30740,
       G30741,G30742,G30743,G30744,G30745,G30746,G30747,G30748,G30749,G30750,G30751,G30752,G30753,G30754,G30755,G30756,G30757,G30758,G30759,G30760,
       G30761,G30762,G30763,G30764,G30765,G30766,G30767,G30768,G30769,G30770,G30771,G30772,G30773,G30774,G30775,G30776,G30777,G30778,G30779,G30780,
       G30781,G30782,G30783,G30784,G30785,G30786,G30787,G30788,G30789,G30790,G30791,G30792,G30793,G30794,G30795,G30796,G30797,G30798,G30799,G30800,
       G30801,G30802,G30803,G30804,G30805,G30806,G30807,G30808,G30809,G30810,G30811,G30812,G30813,G30814,G30815,G30816,G30817,G30818,G30819,G30820,
       G30821,G30822,G30823,G30824,G30825,G30826,G30827,G30828,G30829,G30830,G30831,G30832,G30833,G30834,G30835,G30836,G30837,G30838,G30839,G30840,
       G30841,G30842,G30843,G30844,G30845,G30846,G30847,G30848,G30849,G30850,G30851,G30852,G30853,G30854,G30855,G30856,G30857,G30858,G30859,G30860,
       G30861,G30862,G30863,G30864,G30865,G30866,G30867,G30868,G30869,G30870,G30871,G30872,G30873,G30874,G30875,G30876,G30877,G30878,G30879,G30880,
       G30881,G30882,G30883,G30884,G30885,G30886,G30887,G30888,G30889,G30890,G30891,G30892,G30893,G30894,G30895,G30896,G30897,G30898,G30899,G30900,
       G30901,G30902,G30903,G30904,G30905,G30906,G30907,G30908,G30909,G30910,G30911,G30912,G30913,G30914,G30915,G30916,G30917,G30918,G30919,G30920,
       G30921,G30922,G30923,G30924,G30925,G30926,G30927,G30928,G30929,G30930,G30931,G30932,G30933,G30934,G30935,G30936,G30937,G30938,G30939,G30940,
       G30941,G30942,G30943,G30944,G30945,G30946,G30947,G30948,G30949,G30950,G30951,G30952,G30953,G30954,G30955,G30956,G30957,G30958,G30959,G30960,
       G30961,G30962,G30963,G30964,G30965,G30966,G30967,G30968,G30969,G30970,G30971,G30972,G30973,G30974,G30975,G30976,G30977,G30978,G30979,G30980,
       G30981,G30982,G30983,G30984,G30985,G30986,G30987,G30988,G30989,G30990,G30991,G30992,G30993,G30994,G30995,G30996,G30997,G30998,G30999,G31000,
       G31001,G31002,G31003,G31004,G31005,G31006,G31007,G31008,G31009,G31010,G31011,G31012,G31013,G31014,G31015,G31016,G31017,G31018,G31019,G31020,
       G31021,G31022,G31023,G31024,G31025,G31026,G31027,G31028,G31029,G31030,G31031,G31032,G31033,G31034,G31035,G31036,G31037,G31038,G31039,G31040,
       G31041,G31042,G31043,G31044,G31045,G31046,G31047,G31048,G31049,G31050,G31051,G31052,G31053,G31054,G31055,G31056,G31057,G31058,G31059,G31060,
       G31061,G31062,G31063,G31064,G31065,G31066,G31067,G31068,G31069,G31070,G31071,G31072,G31073,G31074,G31075,G31076,G31077,G31078,G31079,G31080,
       G31081,G31082,G31083,G31084,G31085,G31086,G31087,G31088,G31089,G31090,G31091,G31092,G31093,G31094,G31095,G31096,G31097,G31098,G31099,G31100,
       G31101,G31102,G31103,G31104,G31105,G31106,G31107,G31108,G31109,G31110,G31111,G31112,G31113,G31114,G31115,G31116,G31117,G31118,G31119,G31120,
       G31121,G31122,G31123,G31124,G31125,G31126,G31127,G31128,G31129,G31130,G31131,G31132,G31133,G31134,G31135,G31136,G31137,G31138,G31139,G31140,
       G31141,G31142,G31143,G31144,G31145,G31146,G31147,G31148,G31149,G31150,G31151,G31152,G31153,G31154,G31155,G31156,G31157,G31158,G31159,G31160,
       G31161,G31162,G31163,G31164,G31165,G31166,G31167,G31168,G31169,G31170,G31171,G31172,G31173,G31174,G31175,G31176,G31177,G31178,G31179,G31180,
       G31181,G31182,G31183,G31184,G31185,G31186,G31187,G31188,G31189,G31190,G31191,G31192,G31193,G31194,G31195,G31196,G31197,G31198,G31199,G31200,
       G31201,G31202,G31203,G31204,G31205,G31206,G31207,G31208,G31209,G31210,G31211,G31212,G31213,G31214,G31215,G31216,G31217,G31218,G31219,G31220,
       G31221,G31222,G31223,G31224,G31225,G31226,G31227,G31228,G31229,G31230,G31231,G31232,G31233,G31234,G31235,G31236,G31237,G31238,G31239,G31240,
       G31241,G31242,G31243,G31244,G31245,G31246,G31247,G31248,G31249,G31250,G31251,G31252,G31253,G31254,G31255,G31256,G31257,G31258,G31259,G31260,
       G31261,G31262,G31263,G31264,G31265,G31266,G31267,G31268,G31269,G31270,G31271,G31272,G31273,G31274,G31275,G31276,G31277,G31278,G31279,G31280,
       G31281,G31282,G31283,G31284,G31285,G31286,G31287,G31288,G31289,G31290,G31291,G31292,G31293,G31294,G31295,G31296,G31297,G31298,G31299,G31300,
       G31301,G31302,G31303,G31304,G31305,G31306,G31307,G31308,G31309,G31310,G31311,G31312,G31313,G31314,G31315,G31316,G31317,G31318,G31319,G31320,
       G31321,G31322,G31323,G31324,G31325,G31326,G31327,G31328,G31329,G31330,G31331,G31332,G31333,G31334,G31335,G31336,G31337,G31338,G31339,G31340,
       G31341,G31342,G31343,G31344,G31345,G31346,G31347,G31348,G31349,G31350,G31351,G31352,G31353,G31354,G31355,G31356,G31357,G31358,G31359,G31360,
       G31361,G31362,G31363,G31364,G31365,G31366,G31367,G31368,G31369,G31370,G31371,G31372,G31373,G31374,G31375,G31376,G31377,G31378,G31379,G31380,
       G31381,G31382,G31383,G31384,G31385,G31386,G31387,G31388,G31389,G31390,G31391,G31392,G31393,G31394,G31395,G31396,G31397,G31398,G31399,G31400,
       G31401,G31402,G31403,G31404,G31405,G31406,G31407,G31408,G31409,G31410,G31411,G31412,G31413,G31414,G31415,G31416,G31417,G31418,G31419,G31420,
       G31421,G31422,G31423,G31424,G31425,G31426,G31427,G31428,G31429,G31430,G31431,G31432,G31433,G31434,G31435,G31436,G31437,G31438,G31439,G31440,
       G31441,G31442,G31443,G31444,G31445,G31446,G31447,G31448,G31449,G31450,G31451,G31452,G31453,G31454,G31455,G31456,G31457,G31458,G31459,G31460,
       G31461,G31462,G31463,G31464,G31465,G31466,G31467,G31468,G31469,G31470,G31471,G31472,G31473,G31474,G31475,G31476,G31477,G31478,G31479,G31480,
       G31481,G31482,G31483,G31484,G31485,G31486,G31487,G31488,G31489,G31490,G31491,G31492,G31493,G31494,G31495,G31496,G31497,G31498,G31499,G31500,
       G31501,G31502,G31503,G31504,G31505,G31506,G31507,G31508,G31509,G31510,G31511,G31512,G31513,G31514,G31515,G31516,G31517,G31518,G31519,G31520,
       G31521,G31522,G31523,G31524,G31525,G31526,G31527,G31528,G31529,G31530,G31531,G31532,G31533,G31534,G31535,G31536,G31537,G31538,G31539,G31540,
       G31541,G31542,G31543,G31544,G31545,G31546,G31547,G31548,G31549,G31550,G31551,G31552,G31553,G31554,G31555,G31556,G31557,G31558,G31559,G31560,
       G31561,G31562,G31563,G31564,G31565,G31566,G31567,G31568,G31569,G31570,G31571,G31572,G31573,G31574,G31575,G31576,G31577,G31578,G31579,G31580,
       G31581,G31582,G31583,G31584,G31585,G31586,G31587,G31588,G31589,G31590,G31591,G31592,G31593,G31594,G31595,G31596,G31597,G31598,G31599,G31600,
       G31601,G31602,G31603,G31604,G31605,G31606,G31607,G31608,G31609,G31610,G31611,G31612,G31613,G31614,G31615,G31616,G31617,G31618,G31619,G31620,
       G31621,G31622,G31623,G31624,G31625,G31626,G31627,G31628,G31629,G31630,G31631,G31632,G31633,G31634,G31635,G31636,G31637,G31638,G31639,G31640,
       G31641,G31642,G31643,G31644,G31645,G31646,G31647,G31648,G31649,G31650,G31651,G31652,G31653,G31654,G31655,G31656,G31657,G31658,G31659,G31660,
       G31661,G31662,G31663,G31664,G31665,G31666,G31667,G31668,G31669,G31670,G31671,G31672,G31673,G31674,G31675,G31676,G31677,G31678,G31679,G31680,
       G31681,G31682,G31683,G31684,G31685,G31686,G31687,G31688,G31689,G31690,G31691,G31692,G31693,G31694,G31695,G31696,G31697,G31698,G31699,G31700,
       G31701,G31702,G31703,G31704,G31705,G31706,G31707,G31708,G31709,G31710,G31711,G31712,G31713,G31714,G31715,G31716,G31717,G31718,G31719,G31720,
       G31721,G31722,G31723,G31724,G31725,G31726,G31727,G31728,G31729,G31730,G31731,G31732,G31733,G31734,G31735,G31736,G31737,G31738,G31739,G31740,
       G31741,G31742,G31743,G31744,G31745,G31746,G31747,G31748,G31749,G31750,G31751,G31752,G31753,G31754,G31755,G31756,G31757,G31758,G31759,G31760,
       G31761,G31762,G31763,G31764,G31765,G31766,G31767,G31768,G31769,G31770,G31771,G31772,G31773,G31774,G31775,G31776,G31777,G31778,G31779,G31780,
       G31781,G31782,G31783,G31784,G31785,G31786,G31787,G31788,G31789,G31790,G31791,G31792,G31793,G31794,G31795,G31796,G31797,G31798,G31799,G31800,
       G31801,G31802,G31803,G31804,G31805,G31806,G31807,G31808,G31809,G31810,G31811,G31812,G31813,G31814,G31815,G31816,G31817,G31818,G31819,G31820,
       G31821,G31822,G31823,G31824,G31825,G31826,G31827,G31828,G31829,G31830,G31831,G31832,G31833,G31834,G31835,G31836,G31837,G31838,G31839,G31840,
       G31841,G31842,G31843,G31844,G31845,G31846,G31847,G31848,G31849,G31850,G31851,G31852,G31853,G31854,G31855,G31856,G31857,G31858,G31859,G31860,
       G31861,G31862,G31863,G31864,G31865,G31866,G31867,G31868,G31869,G31870,G31871,G31872,G31873,G31874,G31875,G31876,G31877,G31878,G31879,G31880,
       G31881,G31882,G31883,G31884,G31885,G31886,G31887,G31888,G31889,G31890,G31891,G31892,G31893,G31894,G31895,G31896,G31897,G31898,G31899,G31900,
       G31901,G31902,G31903,G31904,G31905,G31906,G31907,G31908,G31909,G31910,G31911,G31912,G31913,G31914,G31915,G31916,G31917,G31918,G31919,G31920,
       G31921,G31922,G31923,G31924,G31925,G31926,G31927,G31928,G31929,G31930,G31931,G31932,G31933,G31934,G31935,G31936,G31937,G31938,G31939,G31940,
       G31941,G31942,G31943,G31944,G31945,G31946,G31947,G31948,G31949,G31950,G31951,G31952,G31953,G31954,G31955,G31956,G31957,G31958,G31959,G31960,
       G31961,G31962,G31963,G31964,G31965,G31966,G31967,G31968,G31969,G31970,G31971,G31972,G31973,G31974,G31975,G31976,G31977,G31978,G31979,G31980,
       G31981,G31982,G31983,G31984,G31985,G31986,G31987,G31988,G31989,G31990,G31991,G31992,G31993,G31994,G31995,G31996,G31997,G31998,G31999,G32000,
       G32001,G32002,G32003,G32004,G32005,G32006,G32007,G32008,G32009,G32010,G32011,G32012,G32013,G32014,G32015,G32016,G32017,G32018,G32019,G32020,
       G32021,G32022,G32023,G32024,G32025,G32026,G32027,G32028,G32029,G32030,G32031,G32032,G32033,G32034,G32035,G32036,G32037,G32038,G32039,G32040,
       G32041,G32042,G32043,G32044,G32045,G32046,G32047,G32048,G32049,G32050,G32051,G32052,G32053,G32054,G32055,G32056,G32057,G32058,G32059,G32060,
       G32061,G32062,G32063,G32064,G32065,G32066,G32067,G32068,G32069,G32070,G32071,G32072,G32073,G32074,G32075,G32076,G32077,G32078,G32079,G32080,
       G32081,G32082,G32083,G32084,G32085,G32086,G32087,G32088,G32089,G32090,G32091,G32092,G32093,G32094,G32095,G32096,G32097,G32098,G32099,G32100,
       G32101,G32102,G32103,G32104,G32105,G32106,G32107,G32108,G32109,G32110,G32111,G32112,G32113,G32114,G32115,G32116,G32117,G32118,G32119,G32120,
       G32121,G32122,G32123,G32124,G32125,G32126,G32127,G32128,G32129,G32130,G32131,G32132,G32133,G32134,G32135,G32136,G32137,G32138,G32139,G32140,
       G32141,G32142,G32143,G32144,G32145,G32146,G32147,G32148,G32149,G32150,G32151,G32152,G32153,G32154,G32155,G32156,G32157,G32158,G32159,G32160,
       G32161,G32162,G32163,G32164,G32165,G32166,G32167,G32168,G32169,G32170,G32171,G32172,G32173,G32174,G32175,G32176,G32177,G32178,G32179,G32180,
       G32181,G32182,G32183,G32184,G32185,G32186,G32187,G32188,G32189,G32190,G32191,G32192,G32193,G32194,G32195,G32196,G32197,G32198,G32199,G32200,
       G32201,G32202,G32203,G32204,G32205,G32206,G32207,G32208,G32209,G32210,G32211,G32212,G32213,G32214,G32215,G32216,G32217,G32218,G32219,G32220,
       G32221,G32222,G32223,G32224,G32225,G32226,G32227,G32228,G32229,G32230,G32231,G32232,G32233,G32234,G32235,G32236,G32237,G32238,G32239,G32240,
       G32241,G32242,G32243,G32244,G32245,G32246,G32247,G32248,G32249,G32250,G32251,G32252,G32253,G32254,G32255,G32256,G32257,G32258,G32259,G32260,
       G32261,G32262,G32263,G32264,G32265,G32266,G32267,G32268,G32269,G32270,G32271,G32272,G32273,G32274,G32275,G32276,G32277,G32278,G32279,G32280,
       G32281,G32282,G32283,G32284,G32285,G32286,G32287,G32288,G32289,G32290,G32291,G32292,G32293,G32294,G32295,G32296,G32297,G32298,G32299,G32300,
       G32301,G32302,G32303,G32304,G32305,G32306,G32307,G32308,G32309,G32310,G32311,G32312,G32313,G32314,G32315,G32316,G32317,G32318,G32319,G32320,
       G32321,G32322,G32323,G32324,G32325,G32326,G32327,G32328,G32329,G32330,G32331,G32332,G32333,G32334,G32335,G32336,G32337,G32338,G32339,G32340,
       G32341,G32342,G32343,G32344,G32345,G32346,G32347,G32348,G32349,G32350,G32351,G32352,G32353,G32354,G32355,G32356,G32357,G32358,G32359,G32360,
       G32361,G32362,G32363,G32364,G32365,G32366,G32367,G32368,G32369,G32370,G32371,G32372,G32373,G32374,G32375,G32376,G32377,G32378,G32379,G32380,
       G32381,G32382,G32383,G32384,G32385,G32386,G32387,G32388,G32389,G32390,G32391,G32392,G32393,G32394,G32395,G32396,G32397,G32398,G32399,G32400,
       G32401,G32402,G32403,G32404,G32405,G32406,G32407,G32408,G32409,G32410,G32411,G32412,G32413,G32414,G32415,G32416,G32417,G32418,G32419,G32420,
       G32421,G32422,G32423,G32424,G32425,G32426,G32427,G32428,G32429,G32430,G32431,G32432,G32433,G32434,G32435,G32436,G32437,G32438,G32439,G32440,
       G32441,G32442,G32443,G32444,G32445,G32446,G32447,G32448,G32449,G32450,G32451,G32452,G32453,G32454,G32455,G32456,G32457,G32458,G32459,G32460,
       G32461,G32462,G32463,G32464,G32465,G32466,G32467,G32468,G32469,G32470,G32471,G32472,G32473,G32474,G32475,G32476,G32477,G32478,G32479,G32480,
       G32481,G32482,G32483,G32484,G32485,G32486,G32487,G32488,G32489,G32490,G32491,G32492,G32493,G32494,G32495,G32496,G32497,G32498,G32499,G32500,
       G32501,G32502,G32503,G32504,G32505,G32506,G32507,G32508,G32509,G32510,G32511,G32512,G32513,G32514,G32515,G32516,G32517,G32518,G32519,G32520,
       G32521,G32522,G32523,G32524,G32525,G32526,G32527,G32528,G32529,G32530,G32531,G32532,G32533,G32534,G32535,G32536,G32537,G32538,G32539,G32540,
       G32541,G32542,G32543,G32544,G32545,G32546,G32547,G32548,G32549,G32550,G32551,G32552,G32553,G32554,G32555,G32556,G32557,G32558,G32559,G32560,
       G32561,G32562,G32563,G32564,G32565,G32566,G32567,G32568,G32569,G32570,G32571,G32572,G32573,G32574,G32575,G32576,G32577,G32578,G32579,G32580,
       G32581,G32582,G32583,G32584,G32585,G32586,G32587,G32588,G32589,G32590,G32591,G32592,G32593,G32594,G32595,G32596,G32597,G32598,G32599,G32600,
       G32601,G32602,G32603,G32604,G32605,G32606,G32607,G32608,G32609,G32610,G32611,G32612,G32613,G32614,G32615,G32616,G32617,G32618,G32619,G32620,
       G32621,G32622,G32623,G32624,G32625,G32626,G32627,G32628,G32629,G32630,G32631,G32632,G32633,G32634,G32635,G32636,G32637,G32638,G32639,G32640,
       G32641,G32642,G32643,G32644,G32645,G32646,G32647,G32648,G32649,G32650,G32651,G32652,G32653,G32654,G32655,G32656,G32657,G32658,G32659,G32660,
       G32661,G32662,G32663,G32664,G32665,G32666,G32667,G32668,G32669,G32670,G32671,G32672,G32673,G32674,G32675,G32676,G32677,G32678,G32679,G32680,
       G32681,G32682,G32683,G32684,G32685,G32686,G32687,G32688,G32689,G32690,G32691,G32692,G32693,G32694,G32695,G32696,G32697,G32698,G32699,G32700,
       G32701,G32702,G32703,G32704,G32705,G32706,G32707,G32708,G32709,G32710,G32711,G32712,G32713,G32714,G32715,G32716,G32717,G32718,G32719,G32720,
       G32721,G32722,G32723,G32724,G32725,G32726,G32727,G32728,G32729,G32730,G32731,G32732,G32733,G32734,G32735,G32736,G32737,G32738,G32739,G32740,
       G32741,G32742,G32743,G32744,G32745,G32746,G32747,G32748,G32749,G32750,G32751,G32752,G32753,G32754,G32755,G32756,G32757,G32758,G32759,G32760,
       G32761,G32762,G32763,G32764,G32765,G32766,G32767,G32768,G32769,G32770,G32771,G32772,G32773,G32774,G32775,G32776,G32777,G32778,G32779,G32780,
       G32781,G32782,G32783,G32784,G32785,G32786,G32787,G32788,G32789,G32790,G32791,G32792,G32793,G32794,G32795,G32796,G32797,G32798,G32799,G32800,
       G32801,G32802,G32803,G32804,G32805,G32806,G32807,G32808,G32809,G32810,G32811,G32812,G32813,G32814,G32815,G32816,G32817,G32818,G32819,G32820,
       G32821,G32822,G32823,G32824,G32825,G32826,G32827,G32828,G32829,G32830,G32831,G32832,G32833,G32834,G32835,G32836,G32837,G32838,G32839,G32840,
       G32841,G32842,G32843,G32844,G32845,G32846,G32847,G32848,G32849,G32850,G32851,G32852,G32853,G32854,G32855,G32856,G32857,G32858,G32859,G32860,
       G32861,G32862,G32863,G32864,G32865,G32866,G32867,G32868,G32869,G32870,G32871,G32872,G32873,G32874,G32875,G32876,G32877,G32878,G32879,G32880,
       G32881,G32882,G32883,G32884,G32885,G32886,G32887,G32888,G32889,G32890,G32891,G32892,G32893,G32894,G32895,G32896,G32897,G32898,G32899,G32900,
       G32901,G32902,G32903,G32904,G32905,G32906,G32907,G32908,G32909,G32910,G32911,G32912,G32913,G32914,G32915,G32916,G32917,G32918,G32919,G32920,
       G32921,G32922,G32923,G32924,G32925,G32926,G32927,G32928,G32929,G32930,G32931,G32932,G32933,G32934,G32935,G32936,G32937,G32938,G32939,G32940,
       G32941,G32942,G32943,G32944,G32945,G32946,G32947,G32948,G32949,G32950,G32951,G32952,G32953,G32954,G32955,G32956,G32957,G32958,G32959,G32960,
       G32961,G32962,G32963,G32964,G32965,G32966,G32967,G32968,G32969,G32970,G32971,G32972,G32973,G32974,G32975,G32976,G32977,G32978,G32979,G32980,
       G32981,G32982,G32983,G32984,G32985,G32986,G32987,G32988,G32989,G32990,G32991,G32992,G32993,G32994,G32995,G32996,G32997,G32998,G32999,G33000,
       G33001,G33002,G33003,G33004,G33005,G33006,G33007,G33008,G33009,G33010,G33011,G33012,G33013,G33014,G33015,G33016,G33017,G33018,G33019,G33020,
       G33021,G33022,G33023,G33024,G33025,G33026,G33027,G33028,G33029,G33030,G33031,G33032,G33033,G33034,G33035,G33036,G33037,G33038,G33039,G33040,
       G33041,G33042,G33043,G33044,G33045,G33046,G33047,G33048,G33049,G33050,G33051,G33052,G33053,G33054,G33055,G33056,G33057,G33058,G33059,G33060,
       G33061,G33062,G33063,G33064,G33065,G33066,G33067,G33068,G33069,G33070,G33071,G33072,G33073,G33074,G33075,G33076,G33077,G33078,G33079,G33080,
       G33081,G33082,G33083,G33084,G33085,G33086,G33087,G33088,G33089,G33090,G33091,G33092,G33093,G33094,G33095,G33096,G33097,G33098,G33099,G33100,
       G33101,G33102,G33103,G33104,G33105,G33106,G33107,G33108,G33109,G33110,G33111,G33112,G33113,G33114,G33115,G33116,G33117,G33118,G33119,G33120,
       G33121,G33122,G33123,G33124,G33125,G33126,G33127,G33128,G33129,G33130,G33131,G33132,G33133,G33134,G33135,G33136,G33137,G33138,G33139,G33140,
       G33141,G33142,G33143,G33144,G33145,G33146,G33147,G33148,G33149,G33150,G33151,G33152,G33153,G33154,G33155,G33156,G33157,G33158,G33159,G33160,
       G33161,G33162,G33163,G33164,G33165,G33166,G33167,G33168,G33169,G33170,G33171,G33172,G33173,G33174,G33175,G33176,G33177,G33178,G33179,G33180,
       G33181,G33182,G33183,G33184,G33185,G33186,G33187,G33188,G33189,G33190,G33191,G33192,G33193,G33194,G33195,G33196,G33197,G33198,G33199,G33200,
       G33201,G33202,G33203,G33204,G33205,G33206,G33207,G33208,G33209,G33210,G33211,G33212,G33213,G33214,G33215,G33216,G33217,G33218,G33219,G33220,
       G33221,G33222,G33223,G33224,G33225,G33226,G33227,G33228,G33229,G33230,G33231,G33232,G33233,G33234,G33235,G33236,G33237,G33238,G33239,G33240,
       G33241,G33242,G33243,G33244,G33245,G33246,G33247,G33248,G33249,G33250,G33251,G33252,G33253,G33254,G33255,G33256,G33257,G33258,G33259,G33260,
       G33261,G33262,G33263,G33264,G33265,G33266,G33267,G33268,G33269,G33270,G33271,G33272,G33273,G33274,G33275,G33276,G33277,G33278,G33279,G33280,
       G33281,G33282,G33283,G33284,G33285,G33286,G33287,G33288,G33289,G33290,G33291,G33292,G33293,G33294,G33295,G33296,G33297,G33298,G33299,G33300,
       G33301,G33302,G33303,G33304,G33305,G33306,G33307,G33308,G33309,G33310,G33311,G33312,G33313,G33314,G33315,G33316,G33317,G33318,G33319,G33320,
       G33321,G33322,G33323,G33324,G33325,G33326,G33327,G33328,G33329,G33330,G33331,G33332,G33333,G33334,G33335,G33336,G33337,G33338,G33339,G33340,
       G33341,G33342,G33343,G33344,G33345,G33346,G33347,G33348,G33349,G33350,G33351,G33352,G33353,G33354,G33355,G33356,G33357,G33358,G33359,G33360,
       G33361,G33362,G33363,G33364,G33365,G33366,G33367,G33368,G33369,G33370,G33371,G33372,G33373,G33374,G33375,G33376,G33377,G33378,G33379,G33380,
       G33381,G33382,G33383,G33384,G33385,G33386,G33387,G33388,G33389,G33390,G33391,G33392,G33393,G33394,G33395,G33396,G33397,G33398,G33399,G33400,
       G33401,G33402,G33403,G33404,G33405,G33406,G33407,G33408,G33409,G33410,G33411,G33412,G33413,G33414,G33415,G33416,G33417,G33418,G33419,G33420,
       G33421,G33422,G33423,G33424,G33425,G33426,G33427,G33428,G33429,G33430,G33431,G33432,G33433,G33434,G33435,G33436,G33437,G33438,G33439,G33440,
       G33441,G33442,G33443,G33444,G33445,G33446,G33447,G33448,G33449,G33450,G33451,G33452,G33453,G33454,G33455,G33456,G33457,G33458,G33459,G33460,
       G33461,G33462,G33463,G33464,G33465,G33466,G33467,G33468,G33469,G33470,G33471,G33472,G33473,G33474,G33475,G33476,G33477,G33478,G33479,G33480,
       G33481,G33482,G33483,G33484,G33485,G33486,G33487,G33488,G33489,G33490,G33491,G33492,G33493,G33494,G33495,G33496,G33497,G33498,G33499,G33500,
       G33501,G33502,G33503,G33504,G33505,G33506,G33507,G33508,G33509,G33510,G33511,G33512,G33513,G33514,G33515,G33516,G33517,G33518,G33519,G33520,
       G33521,G33522,G33523,G33524,G33525,G33526,G33527,G33528,G33529,G33530,G33531,G33532,G33533,G33534,G33535,G33536,G33537,G33538,G33539,G33540,
       G33541,G33542,G33543,G33544,G33545,G33546,G33547,G33548,G33549,G33550,G33551,G33552,G33553,G33554,G33555,G33556,G33557,G33558,G33559,G33560,
       G33561,G33562,G33563,G33564,G33565,G33566,G33567,G33568,G33569,G33570,G33571,G33572,G33573,G33574,G33575,G33576,G33577,G33578,G33579,G33580,
       G33581,G33582,G33583,G33584,G33585,G33586,G33587,G33588,G33589,G33590,G33591,G33592,G33593,G33594,G33595,G33596,G33597,G33598,G33599,G33600,
       G33601,G33602,G33603,G33604,G33605,G33606,G33607,G33608,G33609,G33610,G33611,G33612,G33613,G33614,G33615,G33616,G33617,G33618,G33619,G33620,
       G33621,G33622,G33623,G33624,G33625,G33626,G33627,G33628,G33629,G33630,G33631,G33632,G33633,G33634,G33635,G33636,G33637,G33638,G33639,G33640,
       G33641,G33642,G33643,G33644,G33645,G33646,G33647,G33648,G33649,G33650,G33651,G33652,G33653,G33654,G33655,G33656,G33657,G33658,G33659,G33660,
       G33661,G33662,G33663,G33664,G33665,G33666,G33667,G33668,G33669,G33670,G33671,G33672,G33673,G33674,G33675,G33676,G33677,G33678,G33679,G33680,
       G33681,G33682,G33683,G33684,G33685,G33686,G33687,G33688,G33689,G33690,G33691,G33692,G33693,G33694,G33695,G33696,G33697,G33698,G33699,G33700,
       G33701,G33702,G33703,G33704,G33705,G33706,G33707,G33708,G33709,G33710,G33711,G33712,G33713,G33714,G33715,G33716,G33717,G33718,G33719,G33720,
       G33721,G33722,G33723,G33724,G33725,G33726,G33727,G33728,G33729,G33730,G33731,G33732,G33733,G33734,G33735,G33736,G33737,G33738,G33739,G33740,
       G33741,G33742,G33743,G33744,G33745,G33746,G33747,G33748,G33749,G33750,G33751,G33752,G33753,G33754,G33755,G33756,G33757,G33758,G33759,G33760,
       G33761,G33762,G33763,G33764,G33765,G33766,G33767,G33768,G33769,G33770,G33771,G33772,G33773,G33774,G33775,G33776,G33777,G33778,G33779,G33780,
       G33781,G33782,G33783,G33784,G33785,G33786,G33787,G33788,G33789,G33790,G33791,G33792,G33793,G33794,G33795,G33796,G33797,G33798,G33799,G33800,
       G33801,G33802,G33803,G33804,G33805,G33806,G33807,G33808,G33809,G33810,G33811,G33812,G33813,G33814,G33815,G33816,G33817,G33818,G33819,G33820,
       G33821,G33822,G33823,G33824,G33825,G33826,G33827,G33828,G33829,G33830,G33831,G33832,G33833,G33834,G33835,G33836,G33837,G33838,G33839,G33840,
       G33841,G33842,G33843,G33844,G33845,G33846,G33847,G33848,G33849,G33850,G33851,G33852,G33853,G33854,G33855,G33856,G33857,G33858,G33859,G33860,
       G33861,G33862,G33863,G33864,G33865,G33866,G33867,G33868,G33869,G33870,G33871,G33872,G33873,G33874,G33875,G33876,G33877,G33878,G33879,G33880,
       G33881,G33882,G33883,G33884,G33885,G33886,G33887,G33888,G33889,G33890,G33891,G33892,G33893,G33894,G33895,G33896,G33897,G33898,G33899,G33900,
       G33901,G33902,G33903,G33904,G33905,G33906,G33907,G33908,G33909,G33910,G33911,G33912,G33913,G33914,G33915,G33916,G33917,G33918,G33919,G33920,
       G33921,G33922,G33923,G33924,G33925,G33926,G33927,G33928,G33929,G33930,G33931,G33932,G33933,G33934,G33935,G33936,G33937,G33938,G33939,G33940,
       G33941,G33942,G33943,G33944,G33945,G33946,G33947,G33948,G33949,G33950,G33951,G33952,G33953,G33954,G33955,G33956,G33957,G33958,G33959,G33960,
       G33961,G33962,G33963,G33964,G33965,G33966,G33967,G33968,G33969,G33970,G33971,G33972,G33973,G33974,G33975,G33976,G33977,G33978,G33979,G33980,
       G33981,G33982,G33983,G33984,G33985,G33986,G33987,G33988,G33989,G33990,G33991,G33992,G33993,G33994,G33995,G33996,G33997,G33998,G33999,G34000,
       G34001,G34002,G34003,G34004,G34005,G34006,G34007,G34008,G34009,G34010,G34011,G34012,G34013,G34014,G34015,G34016,G34017,G34018,G34019,G34020,
       G34021,G34022,G34023,G34024,G34025,G34026,G34027,G34028,G34029,G34030,G34031,G34032,G34033,G34034,G34035,G34036,G34037,G34038,G34039,G34040,
       G34041,G34042,G34043,G34044,G34045,G34046,G34047,G34048,G34049,G34050,G34051,G34052,G34053,G34054,G34055,G34056,G34057,G34058,G34059,G34060,
       G34061,G34062,G34063,G34064,G34065,G34066,G34067,G34068,G34069,G34070,G34071,G34072,G34073,G34074,G34075,G34076,G34077,G34078,G34079,G34080,
       G34081,G34082,G34083,G34084,G34085,G34086,G34087,G34088,G34089,G34090,G34091,G34092,G34093,G34094,G34095,G34096,G34097,G34098,G34099,G34100,
       G34101,G34102,G34103,G34104,G34105,G34106,G34107,G34108,G34109,G34110,G34111,G34112,G34113,G34114,G34115,G34116,G34117,G34118,G34119,G34120,
       G34121,G34122,G34123,G34124,G34125,G34126,G34127,G34128,G34129,G34130,G34131,G34132,G34133,G34134,G34135,G34136,G34137,G34138,G34139,G34140,
       G34141,G34142,G34143,G34144,G34145,G34146,G34147,G34148,G34149,G34150,G34151,G34152,G34153,G34154,G34155,G34156,G34157,G34158,G34159,G34160,
       G34161,G34162,G34163,G34164,G34165,G34166,G34167,G34168,G34169,G34170,G34171,G34172,G34173,G34174,G34175,G34176,G34177,G34178,G34179,G34180,
       G34181,G34182,G34183,G34184,G34185,G34186,G34187,G34188,G34189,G34190,G34191,G34192,G34193,G34194,G34195,G34196,G34197,G34198,G34199,G34200,
       G34201,G34202,G34203,G34204,G34205,G34206,G34207,G34208,G34209,G34210,G34211,G34212,G34213,G34214,G34215,G34216,G34217,G34218,G34219,G34220,
       G34221,G34222,G34223,G34224,G34225,G34226,G34227,G34228,G34229,G34230,G34231,G34232,G34233,G34234,G34235,G34236,G34237,G34238,G34239,G34240,
       G34241,G34242,G34243,G34244,G34245,G34246,G34247,G34248,G34249,G34250,G34251,G34252,G34253,G34254,G34255,G34256,G34257,G34258,G34259,G34260,
       G34261,G34262,G34263,G34264,G34265,G34266,G34267,G34268,G34269,G34270,G34271,G34272,G34273,G34274,G34275,G34276,G34277,G34278,G34279,G34280,
       G34281,G34282,G34283,G34284,G34285,G34286,G34287,G34288,G34289,G34290,G34291,G34292,G34293,G34294,G34295,G34296,G34297,G34298,G34299,G34300,
       G34301,G34302,G34303,G34304,G34305,G34306,G34307,G34308,G34309,G34310,G34311,G34312,G34313,G34314,G34315,G34316,G34317,G34318,G34319,G34320,
       G34321,G34322,G34323,G34324,G34325,G34326,G34327,G34328,G34329,G34330,G34331,G34332,G34333,G34334,G34335,G34336,G34337,G34338,G34339,G34340,
       G34341,G34342,G34343,G34344,G34345,G34346,G34347,G34348,G34349,G34350,G34351,G34352,G34353,G34354,G34355,G34356,G34357,G34358,G34359,G34360,
       G34361,G34362,G34363,G34364,G34365,G34366,G34367,G34368,G34369,G34370,G34371,G34372,G34373,G34374,G34375,G34376,G34377,G34378,G34379,G34380,
       G34381,G34382,G34383,G34384,G34385,G34386,G34387,G34388,G34389,G34390,G34391,G34392,G34393,G34394,G34395,G34396,G34397,G34398,G34399,G34400,
       G34401,G34402,G34403,G34404,G34405,G34406,G34407,G34408,G34409,G34410,G34411,G34412,G34413,G34414,G34415,G34416,G34417,G34418,G34419,G34420,
       G34421,G34422,G34423,G34424,G34425,G34426,G34427,G34428,G34429,G34430,G34431,G34432,G34433,G34434,G34435,G34436,G34437,G34438,G34439,G34440,
       G34441,G34442,G34443,G34444,G34445,G34446,G34447,G34448,G34449,G34450,G34451,G34452,G34453,G34454,G34455,G34456,G34457,G34458,G34459,G34460,
       G34461,G34462,G34463,G34464,G34465,G34466,G34467,G34468,G34469,G34470,G34471,G34472,G34473,G34474,G34475,G34476,G34477,G34478,G34479,G34480,
       G34481,G34482,G34483,G34484,G34485,G34486,G34487,G34488,G34489,G34490,G34491,G34492,G34493,G34494,G34495,G34496,G34497,G34498,G34499,G34500,
       G34501,G34502,G34503,G34504,G34505,G34506,G34507,G34508,G34509,G34510,G34511,G34512,G34513,G34514,G34515,G34516,G34517,G34518,G34519,G34520,
       G34521,G34522,G34523,G34524,G34525,G34526,G34527,G34528,G34529,G34530,G34531,G34532,G34533,G34534,G34535,G34536,G34537,G34538,G34539,G34540,
       G34541,G34542,G34543,G34544,G34545,G34546,G34547,G34548,G34549,G34550,G34551,G34552,G34553,G34554,G34555,G34556,G34557,G34558,G34559,G34560,
       G34561,G34562,G34563,G34564,G34565,G34566,G34567,G34568,G34569,G34570,G34571,G34572,G34573,G34574,G34575,G34576,G34577,G34578,G34579,G34580,
       G34581,G34582,G34583,G34584,G34585,G34586,G34587,G34588,G34589,G34590,G34591,G34592,G34593,G34594,G34595,G34596,G34597,G34598,G34599,G34600,
       G34601,G34602,G34603,G34604,G34605,G34606,G34607,G34608,G34609,G34610,G34611,G34612,G34613,G34614,G34615,G34616,G34617,G34618,G34619,G34620,
       G34621,G34622,G34623,G34624,G34625,G34626,G34627,G34628,G34629,G34630,G34631,G34632,G34633,G34634,G34635,G34636,G34637,G34638,G34639,G34640,
       G34641,G34642,G34643,G34644,G34645,G34646,G34647,G34648,G34649,G34650,G34651,G34652,G34653,G34654,G34655,G34656,G34657,G34658,G34659,G34660,
       G34661,G34662,G34663,G34664,G34665,G34666,G34667,G34668,G34669,G34670,G34671,G34672,G34673,G34674,G34675,G34676,G34677,G34678,G34679,G34680,
       G34681,G34682,G34683,G34684,G34685,G34686,G34687,G34688,G34689,G34690,G34691,G34692,G34693,G34694,G34695,G34696,G34697,G34698,G34699,G34700,
       G34701,G34702,G34703,G34704,G34705,G34706,G34707,G34708,G34709,G34710,G34711,G34712,G34713,G34714,G34715,G34716,G34717,G34718,G34719,G34720,
       G34721,G34722,G34723,G34724,G34725,G34726,G34727,G34728,G34729,G34730,G34731,G34732,G34733,G34734,G34735,G34736,G34737,G34738,G34739,G34740,
       G34741,G34742,G34743,G34744,G34745,G34746,G34747,G34748,G34749,G34750,G34751,G34752,G34753,G34754,G34755,G34756,G34757,G34758,G34759,G34760,
       G34761,G34762,G34763,G34764,G34765,G34766,G34767,G34768,G34769,G34770,G34771,G34772,G34773,G34774,G34775,G34776,G34777,G34778,G34779,G34780,
       G34781,G34782,G34783,G34784,G34785,G34786,G34787,G34788,G34789,G34790,G34791,G34792,G34793,G34794,G34795,G34796,G34797,G34798,G34799,G34800,
       G34801,G34802,G34803,G34804,G34805,G34806,G34807,G34808,G34809,G34810,G34811,G34812,G34813,G34814,G34815,G34816,G34817,G34818,G34819,G34820,
       G34821,G34822,G34823,G34824,G34825,G34826,G34827,G34828,G34829,G34830,G34831,G34832,G34833,G34834,G34835,G34836,G34837,G34838,G34839,G34840,
       G34841,G34842,G34843,G34844,G34845,G34846,G34847,G34848,G34849,G34850,G34851,G34852,G34853,G34854,G34855,G34856,G34857,G34858,G34859,G34860,
       G34861,G34862,G34863,G34864,G34865,G34866,G34867,G34868,G34869,G34870,G34871,G34872,G34873,G34874,G34875,G34876,G34877,G34878,G34879,G34880,
       G34881,G34882,G34883,G34884,G34885,G34886,G34887,G34888,G34889,G34890,G34891,G34892,G34893,G34894,G34895,G34896,G34897,G34898,G34899,G34900,
       G34901,G34902,G34903,G34904,G34905,G34906,G34907,G34908,G34909,G34910,G34911,G34912,G34913,G34914,G34915,G34916,G34917,G34918,G34919,G34920,
       G34921,G34922,G34923,G34924,G34925,G34926,G34927,G34928,G34929,G34930,G34931,G34932,G34933,G34934,G34935,G34936,G34937,G34938,G34939,G34940,
       G34941,G34942,G34943,G34944,G34945,G34946,G34947,G34948,G34949,G34950,G34951,G34952,G34953,G34954,G34955,G34956,G34957,G34958,G34959,G34960,
       G34961,G34962,G34963,G34964,G34965,G34966,G34967,G34968,G34969,G34970,G34971,G34972,G34973,G34974,G34975,G34976,G34977,G34978,G34979,G34980,
       G34981,G34982,G34983,G34984,G34985,G34986,G34987,G34988,G34989,G34990,G34991,G34992,G34993,G34994,G34995,G34996,G34997,G34998,G34999,G35000,
       G35001,G35002,G35003,G35004,G35005,G35006,G35007,G35008,G35009,G35010,G35011,G35012,G35013,G35014,G35015,G35016,G35017,G35018,G35019,G35020,
       G35021,G35022,G35023,G35024,G35025,G35026,G35027,G35028,G35029,G35030,G35031,G35032,G35033,G35034,G35035,G35036,G35037,G35038,G35039,G35040,
       G35041,G35042,G35043,G35044,G35045,G35046,G35047,G35048,G35049,G35050,G35051,G35052,G35053,G35054,G35055,G35056,G35057,G35058,G35059,G35060,
       G35061,G35062,G35063,G35064,G35065,G35066,G35067,G35068,G35069,G35070,G35071,G35072,G35073,G35074,G35075,G35076,G35077,G35078,G35079,G35080,
       G35081,G35082,G35083,G35084,G35085,G35086,G35087,G35088,G35089,G35090,G35091,G35092,G35093,G35094,G35095,G35096,G35097,G35098,G35099,G35100,
       G35101,G35102,G35103,G35104,G35105,G35106,G35107,G35108,G35109,G35110,G35111,G35112,G35113,G35114,G35115,G35116,G35117,G35118,G35119,G35120,
       G35121,G35122,G35123,G35124,G35125,G35126,G35127,G35128,G35129,G35130,G35131,G35132,G35133,G35134,G35135,G35136,G35137,G35138,G35139,G35140,
       G35141,G35142,G35143,G35144,G35145,G35146,G35147,G35148,G35149,G35150,G35151,G35152,G35153,G35154,G35155,G35156,G35157,G35158,G35159,G35160,
       G35161,G35162,G35163,G35164,G35165,G35166,G35167,G35168,G35169,G35170,G35171,G35172,G35173,G35174,G35175,G35176,G35177,G35178,G35179,G35180,
       G35181,G35182,G35183,G35184,G35185,G35186,G35187,G35188,G35189,G35190,G35191,G35192,G35193,G35194,G35195,G35196,G35197,G35198,G35199,G35200,
       G35201,G35202,G35203,G35204,G35205,G35206,G35207,G35208,G35209,G35210,G35211,G35212,G35213,G35214,G35215,G35216,G35217,G35218,G35219,G35220,
       G35221,G35222,G35223,G35224,G35225,G35226,G35227,G35228,G35229,G35230,G35231,G35232,G35233,G35234,G35235,G35236,G35237,G35238,G35239,G35240,
       G35241,G35242,G35243,G35244,G35245,G35246,G35247,G35248,G35249,G35250,G35251,G35252,G35253,G35254,G35255,G35256,G35257,G35258,G35259,G35260,
       G35261,G35262,G35263,G35264,G35265,G35266,G35267,G35268,G35269,G35270,G35271,G35272,G35273,G35274,G35275,G35276,G35277,G35278,G35279,G35280,
       G35281,G35282,G35283,G35284,G35285,G35286,G35287,G35288,G35289,G35290,G35291,G35292,G35293,G35294,G35295,G35296,G35297,G35298,G35299,G35300,
       G35301,G35302,G35303,G35304,G35305,G35306,G35307,G35308,G35309,G35310,G35311,G35312,G35313,G35314,G35315,G35316,G35317,G35318,G35319,G35320,
       G35321,G35322,G35323,G35324,G35325,G35326,G35327,G35328,G35329,G35330,G35331,G35332,G35333,G35334,G35335,G35336,G35337,G35338,G35339,G35340,
       G35341,G35342,G35343,G35344,G35345,G35346,G35347,G35348,G35349,G35350,G35351,G35352,G35353,G35354,G35355,G35356,G35357,G35358,G35359,G35360,
       G35361,G35362,G35363,G35364,G35365,G35366,G35367,G35368,G35369,G35370,G35371,G35372,G35373,G35374,G35375,G35376,G35377,G35378,G35379,G35380,
       G35381,G35382,G35383,G35384,G35385,G35386,G35387,G35388,G35389,G35390,G35391,G35392,G35393,G35394,G35395,G35396,G35397,G35398,G35399,G35400,
       G35401,G35402,G35403,G35404,G35405,G35406,G35407,G35408,G35409,G35410,G35411,G35412,G35413,G35414,G35415,G35416,G35417,G35418,G35419,G35420,
       G35421,G35422,G35423,G35424,G35425,G35426,G35427,G35428,G35429,G35430,G35431,G35432,G35433,G35434,G35435,G35436,G35437,G35438,G35439,G35440,
       G35441,G35442,G35443,G35444,G35445,G35446,G35447,G35448,G35449,G35450,G35451,G35452,G35453,G35454,G35455,G35456,G35457,G35458,G35459,G35460,
       G35461,G35462,G35463,G35464,G35465,G35466,G35467,G35468,G35469,G35470,G35471,G35472,G35473,G35474,G35475,G35476,G35477,G35478,G35479,G35480,
       G35481,G35482,G35483,G35484,G35485,G35486,G35487,G35488,G35489,G35490,G35491,G35492,G35493,G35494,G35495,G35496,G35497,G35498,G35499,G35500,
       G35501,G35502,G35503,G35504,G35505,G35506,G35507,G35508,G35509,G35510,G35511,G35512,G35513,G35514,G35515,G35516,G35517,G35518,G35519,G35520,
       G35521,G35522,G35523,G35524,G35525,G35526,G35527,G35528,G35529,G35530,G35531,G35532,G35533,G35534,G35535,G35536,G35537,G35538,G35539,G35540,
       G35541,G35542,G35543,G35544,G35545,G35546,G35547,G35548,G35549,G35550,G35551,G35552,G35553,G35554,G35555,G35556,G35557,G35558,G35559,G35560,
       G35561,G35562,G35563,G35564,G35565,G35566,G35567,G35568,G35569,G35570,G35571,G35572,G35573,G35574,G35575,G35576,G35577,G35578,G35579,G35580,
       G35581,G35582,G35583,G35584,G35585,G35586,G35587,G35588,G35589,G35590,G35591,G35592,G35593,G35594,G35595,G35596,G35597,G35598,G35599,G35600,
       G35601,G35602,G35603,G35604,G35605,G35606,G35607,G35608,G35609,G35610,G35611,G35612,G35613,G35614,G35615,G35616,G35617,G35618,G35619,G35620,
       G35621,G35622,G35623,G35624,G35625,G35626,G35627,G35628,G35629,G35630,G35631,G35632,G35633,G35634,G35635,G35636,G35637,G35638,G35639,G35640,
       G35641,G35642,G35643,G35644,G35645,G35646,G35647,G35648,G35649,G35650,G35651,G35652,G35653,G35654,G35655,G35656,G35657,G35658,G35659,G35660,
       G35661,G35662,G35663,G35664,G35665,G35666,G35667,G35668,G35669,G35670,G35671,G35672,G35673,G35674,G35675,G35676,G35677,G35678,G35679,G35680,
       G35681,G35682,G35683,G35684,G35685,G35686,G35687,G35688,G35689,G35690,G35691,G35692,G35693,G35694,G35695,G35696,G35697,G35698,G35699,G35700,
       G35701,G35702,G35703,G35704,G35705,G35706,G35707,G35708,G35709,G35710,G35711,G35712,G35713,G35714,G35715,G35716,G35717,G35718,G35719,G35720,
       G35721,G35722,G35723,G35724,G35725,G35726,G35727,G35728,G35729,G35730,G35731,G35732,G35733,G35734,G35735,G35736,G35737,G35738,G35739,G35740,
       G35741,G35742,G35743,G35744,G35745,G35746,G35747,G35748,G35749,G35750,G35751,G35752,G35753,G35754,G35755,G35756,G35757,G35758,G35759,G35760,
       G35761,G35762,G35763,G35764,G35765,G35766,G35767,G35768,G35769,G35770,G35771,G35772,G35773,G35774,G35775,G35776,G35777,G35778,G35779,G35780,
       G35781,G35782,G35783,G35784,G35785,G35786,G35787,G35788,G35789,G35790,G35791,G35792,G35793,G35794,G35795,G35796,G35797,G35798,G35799,G35800,
       G35801,G35802,G35803,G35804,G35805,G35806,G35807,G35808,G35809,G35810,G35811,G35812,G35813,G35814,G35815,G35816,G35817,G35818,G35819,G35820,
       G35821,G35822,G35823,G35824,G35825,G35826,G35827,G35828,G35829,G35830,G35831,G35832,G35833,G35834,G35835,G35836,G35837,G35838,G35839,G35840,
       G35841,G35842,G35843,G35844,G35845,G35846,G35847,G35848,G35849,G35850,G35851,G35852,G35853,G35854,G35855,G35856,G35857,G35858,G35859,G35860,
       G35861,G35862,G35863,G35864,G35865,G35866,G35867,G35868,G35869,G35870,G35871,G35872,G35873,G35874,G35875,G35876,G35877,G35878,G35879,G35880,
       G35881,G35882,G35883,G35884,G35885,G35886,G35887,G35888,G35889,G35890,G35891,G35892,G35893,G35894,G35895,G35896,G35897,G35898,G35899,G35900,
       G35901,G35902,G35903,G35904,G35905,G35906,G35907,G35908,G35909,G35910,G35911,G35912,G35913,G35914,G35915,G35916,G35917,G35918,G35919,G35920,
       G35921,G35922,G35923,G35924,G35925,G35926,G35927,G35928,G35929,G35930,G35931,G35932,G35933,G35934,G35935,G35936,G35937,G35938,G35939,G35940,
       G35941,G35942,G35943,G35944,G35945,G35946,G35947,G35948,G35949,G35950,G35951,G35952,G35953,G35954,G35955,G35956,G35957,G35958,G35959,G35960,
       G35961,G35962,G35963,G35964,G35965,G35966,G35967,G35968,G35969,G35970,G35971,G35972,G35973,G35974,G35975,G35976,G35977,G35978,G35979,G35980,
       G35981,G35982,G35983,G35984,G35985,G35986,G35987,G35988,G35989,G35990,G35991,G35992,G35993,G35994,G35995,G35996,G35997,G35998,G35999,G36000,
       G36001,G36002,G36003,G36004,G36005,G36006,G36007,G36008,G36009,G36010,G36011,G36012,G36013,G36014,G36015,G36016,G36017,G36018,G36019,G36020,
       G36021,G36022,G36023,G36024,G36025,G36026,G36027,G36028,G36029,G36030,G36031,G36032,G36033,G36034,G36035,G36036,G36037,G36038,G36039,G36040,
       G36041,G36042,G36043,G36044,G36045,G36046,G36047,G36048,G36049,G36050,G36051,G36052,G36053,G36054,G36055,G36056,G36057,G36058,G36059,G36060,
       G36061,G36062,G36063,G36064,G36065,G36066,G36067,G36068,G36069,G36070,G36071,G36072,G36073,G36074,G36075,G36076,G36077,G36078,G36079,G36080,
       G36081,G36082,G36083,G36084,G36085,G36086,G36087,G36088,G36089,G36090,G36091,G36092,G36093,G36094,G36095,G36096,G36097,G36098,G36099,G36100,
       G36101,G36102,G36103,G36104,G36105,G36106,G36107,G36108,G36109,G36110,G36111,G36112,G36113,G36114,G36115,G36116,G36117,G36118,G36119,G36120,
       G36121,G36122,G36123,G36124,G36125,G36126,G36127,G36128,G36129,G36130,G36131,G36132,G36133,G36134,G36135,G36136,G36137,G36138,G36139,G36140,
       G36141,G36142,G36143,G36144,G36145,G36146,G36147,G36148,G36149,G36150,G36151,G36152,G36153,G36154,G36155,G36156,G36157,G36158,G36159,G36160,
       G36161,G36162,G36163,G36164,G36165,G36166,G36167,G36168,G36169,G36170,G36171,G36172,G36173,G36174,G36175,G36176,G36177,G36178,G36179,G36180,
       G36181,G36182,G36183,G36184,G36185,G36186,G36187,G36188,G36189,G36190,G36191,G36192,G36193,G36194,G36195,G36196,G36197,G36198,G36199,G36200,
       G36201,G36202,G36203,G36204,G36205,G36206,G36207,G36208,G36209,G36210,G36211,G36212,G36213,G36214,G36215,G36216,G36217,G36218,G36219,G36220,
       G36221,G36222,G36223,G36224,G36225,G36226,G36227,G36228,G36229,G36230,G36231,G36232,G36233,G36234,G36235,G36236,G36237,G36238,G36239,G36240,
       G36241,G36242,G36243,G36244,G36245,G36246,G36247,G36248,G36249,G36250,G36251,G36252,G36253,G36254,G36255,G36256,G36257,G36258,G36259,G36260,
       G36261,G36262,G36263,G36264,G36265,G36266,G36267,G36268,G36269,G36270,G36271,G36272,G36273,G36274,G36275,G36276,G36277,G36278,G36279,G36280,
       G36281,G36282,G36283,G36284,G36285,G36286,G36287,G36288,G36289,G36290,G36291,G36292,G36293,G36294,G36295,G36296,G36297,G36298,G36299,G36300,
       G36301,G36302,G36303,G36304,G36305,G36306,G36307,G36308,G36309,G36310,G36311,G36312,G36313,G36314,G36315,G36316,G36317,G36318,G36319,G36320,
       G36321,G36322,G36323,G36324,G36325,G36326,G36327,G36328,G36329,G36330,G36331,G36332,G36333,G36334,G36335,G36336,G36337,G36338,G36339,G36340,
       G36341,G36342,G36343,G36344,G36345,G36346,G36347,G36348,G36349,G36350,G36351,G36352,G36353,G36354,G36355,G36356,G36357,G36358,G36359,G36360,
       G36361,G36362,G36363,G36364,G36365,G36366,G36367,G36368,G36369,G36370,G36371,G36372,G36373,G36374,G36375,G36376,G36377,G36378,G36379,G36380,
       G36381,G36382,G36383,G36384,G36385,G36386,G36387,G36388,G36389,G36390,G36391,G36392,G36393,G36394,G36395,G36396,G36397,G36398,G36399,G36400,
       G36401,G36402,G36403,G36404,G36405,G36406,G36407,G36408,G36409,G36410,G36411,G36412,G36413,G36414,G36415,G36416,G36417,G36418,G36419,G36420,
       G36421,G36422,G36423,G36424,G36425,G36426,G36427,G36428,G36429,G36430,G36431,G36432,G36433,G36434,G36435,G36436,G36437,G36438,G36439,G36440,
       G36441,G36442,G36443,G36444,G36445,G36446,G36447,G36448,G36449,G36450,G36451,G36452,G36453,G36454,G36455,G36456,G36457,G36458,G36459,G36460,
       G36461,G36462,G36463,G36464,G36465,G36466,G36467,G36468,G36469,G36470,G36471,G36472,G36473,G36474,G36475,G36476,G36477,G36478,G36479,G36480,
       G36481,G36482,G36483,G36484,G36485,G36486,G36487,G36488,G36489,G36490,G36491,G36492,G36493,G36494,G36495,G36496,G36497,G36498,G36499,G36500,
       G36501,G36502,G36503,G36504,G36505,G36506,G36507,G36508,G36509,G36510,G36511,G36512,G36513,G36514,G36515,G36516,G36517,G36518,G36519,G36520,
       G36521,G36522,G36523,G36524,G36525,G36526,G36527,G36528,G36529,G36530,G36531,G36532,G36533,G36534,G36535,G36536,G36537,G36538,G36539,G36540,
       G36541,G36542,G36543,G36544,G36545,G36546,G36547,G36548,G36549,G36550,G36551,G36552,G36553,G36554,G36555,G36556,G36557,G36558,G36559,G36560,
       G36561,G36562,G36563,G36564,G36565,G36566,G36567,G36568,G36569,G36570,G36571,G36572,G36573,G36574,G36575,G36576,G36577,G36578,G36579,G36580,
       G36581,G36582,G36583,G36584,G36585,G36586,G36587,G36588,G36589,G36590,G36591,G36592,G36593,G36594,G36595,G36596,G36597,G36598,G36599,G36600,
       G36601,G36602,G36603,G36604,G36605,G36606,G36607,G36608,G36609,G36610,G36611,G36612,G36613,G36614,G36615,G36616,G36617,G36618,G36619,G36620,
       G36621,G36622,G36623,G36624,G36625,G36626,G36627,G36628,G36629,G36630,G36631,G36632,G36633,G36634,G36635,G36636,G36637,G36638,G36639,G36640,
       G36641,G36642,G36643,G36644,G36645,G36646,G36647,G36648,G36649,G36650,G36651,G36652,G36653,G36654,G36655,G36656,G36657,G36658,G36659,G36660,
       G36661,G36662,G36663,G36664,G36665,G36666,G36667,G36668,G36669,G36670,G36671,G36672,G36673,G36674,G36675,G36676,G36677,G36678,G36679,G36680,
       G36681,G36682,G36683,G36684,G36685,G36686,G36687,G36688,G36689,G36690,G36691,G36692,G36693,G36694,G36695,G36696,G36697,G36698,G36699,G36700,
       G36701,G36702,G36703,G36704,G36705,G36706,G36707,G36708,G36709,G36710,G36711,G36712,G36713,G36714,G36715,G36716,G36717,G36718,G36719,G36720,
       G36721,G36722,G36723,G36724,G36725,G36726,G36727,G36728,G36729,G36730,G36731,G36732,G36733,G36734,G36735,G36736,G36737,G36738,G36739,G36740,
       G36741,G36742,G36743,G36744,G36745,G36746,G36747,G36748,G36749,G36750,G36751,G36752,G36753,G36754,G36755,G36756,G36757,G36758,G36759,G36760,
       G36761,G36762,G36763,G36764,G36765,G36766,G36767,G36768,G36769,G36770,G36771,G36772,G36773,G36774,G36775,G36776,G36777,G36778,G36779,G36780,
       G36781,G36782,G36783,G36784,G36785,G36786,G36787,G36788,G36789,G36790,G36791,G36792,G36793,G36794,G36795,G36796,G36797,G36798,G36799,G36800,
       G36801,G36802,G36803,G36804,G36805,G36806,G36807,G36808,G36809,G36810,G36811,G36812,G36813,G36814,G36815,G36816,G36817,G36818,G36819,G36820,
       G36821,G36822,G36823,G36824,G36825,G36826,G36827,G36828,G36829,G36830,G36831,G36832,G36833,G36834,G36835,G36836,G36837,G36838,G36839,G36840,
       G36841,G36842,G36843,G36844,G36845,G36846,G36847,G36848,G36849,G36850,G36851,G36852,G36853,G36854,G36855,G36856,G36857,G36858,G36859,G36860,
       G36861,G36862,G36863,G36864,G36865,G36866,G36867,G36868,G36869,G36870,G36871,G36872,G36873,G36874,G36875,G36876,G36877,G36878,G36879,G36880,
       G36881,G36882,G36883,G36884,G36885,G36886,G36887,G36888,G36889,G36890,G36891,G36892,G36893,G36894,G36895,G36896,G36897,G36898,G36899,G36900,
       G36901,G36902,G36903,G36904,G36905,G36906,G36907,G36908,G36909,G36910,G36911,G36912,G36913,G36914,G36915,G36916,G36917,G36918,G36919,G36920,
       G36921,G36922,G36923,G36924,G36925,G36926,G36927,G36928,G36929,G36930,G36931,G36932,G36933,G36934,G36935,G36936,G36937,G36938,G36939,G36940,
       G36941,G36942,G36943,G36944,G36945,G36946,G36947,G36948,G36949,G36950,G36951,G36952,G36953,G36954,G36955,G36956,G36957,G36958,G36959,G36960,
       G36961,G36962,G36963,G36964,G36965,G36966,G36967,G36968,G36969,G36970,G36971,G36972,G36973,G36974,G36975,G36976,G36977,G36978,G36979,G36980,
       G36981,G36982,G36983,G36984,G36985,G36986,G36987,G36988,G36989,G36990,G36991,G36992,G36993,G36994,G36995,G36996,G36997,G36998,G36999,G37000,
       G37001,G37002,G37003,G37004,G37005,G37006,G37007,G37008,G37009,G37010,G37011,G37012,G37013,G37014,G37015,G37016,G37017,G37018,G37019,G37020,
       G37021,G37022,G37023,G37024,G37025,G37026,G37027,G37028,G37029,G37030,G37031,G37032,G37033,G37034,G37035,G37036,G37037,G37038,G37039,G37040,
       G37041,G37042,G37043,G37044,G37045,G37046,G37047,G37048,G37049,G37050,G37051,G37052,G37053,G37054,G37055,G37056,G37057,G37058,G37059,G37060,
       G37061,G37062,G37063,G37064,G37065,G37066,G37067,G37068,G37069,G37070,G37071,G37072,G37073,G37074,G37075,G37076,G37077,G37078,G37079,G37080,
       G37081,G37082,G37083,G37084,G37085,G37086,G37087,G37088,G37089,G37090,G37091,G37092,G37093,G37094,G37095,G37096,G37097,G37098,G37099,G37100,
       G37101,G37102,G37103,G37104,G37105,G37106,G37107,G37108,G37109,G37110,G37111,G37112,G37113,G37114,G37115,G37116,G37117,G37118,G37119,G37120,
       G37121,G37122,G37123,G37124,G37125,G37126,G37127,G37128,G37129,G37130,G37131,G37132,G37133,G37134,G37135,G37136,G37137,G37138,G37139,G37140,
       G37141,G37142,G37143,G37144,G37145,G37146,G37147,G37148,G37149,G37150,G37151,G37152,G37153,G37154,G37155,G37156,G37157,G37158,G37159,G37160,
       G37161,G37162,G37163,G37164,G37165,G37166,G37167,G37168,G37169,G37170,G37171,G37172,G37173,G37174,G37175,G37176,G37177,G37178,G37179,G37180,
       G37181,G37182,G37183,G37184,G37185,G37186,G37187,G37188,G37189,G37190,G37191,G37192,G37193,G37194,G37195,G37196,G37197,G37198,G37199,G37200,
       G37201,G37202,G37203,G37204,G37205,G37206,G37207,G37208,G37209,G37210,G37211,G37212,G37213,G37214,G37215,G37216,G37217,G37218,G37219,G37220,
       G37221,G37222,G37223,G37224,G37225,G37226,G37227,G37228,G37229,G37230,G37231,G37232,G37233,G37234,G37235,G37236,G37237,G37238,G37239,G37240,
       G37241,G37242,G37243,G37244,G37245,G37246,G37247,G37248,G37249,G37250,G37251,G37252,G37253,G37254,G37255,G37256,G37257,G37258,G37259,G37260,
       G37261,G37262,G37263,G37264,G37265,G37266,G37267,G37268,G37269,G37270,G37271,G37272,G37273,G37274,G37275,G37276,G37277,G37278,G37279,G37280,
       G37281,G37282,G37283,G37284,G37285,G37286,G37287,G37288,G37289,G37290,G37291,G37292,G37293,G37294,G37295,G37296,G37297,G37298,G37299,G37300,
       G37301,G37302,G37303,G37304,G37305,G37306,G37307,G37308,G37309,G37310,G37311,G37312,G37313,G37314,G37315,G37316,G37317,G37318,G37319,G37320,
       G37321,G37322,G37323,G37324,G37325,G37326,G37327,G37328,G37329,G37330,G37331,G37332,G37333,G37334,G37335,G37336,G37337,G37338,G37339,G37340,
       G37341,G37342,G37343,G37344,G37345,G37346,G37347,G37348,G37349,G37350,G37351,G37352,G37353,G37354,G37355,G37356,G37357,G37358,G37359,G37360,
       G37361,G37362,G37363,G37364,G37365,G37366,G37367,G37368,G37369,G37370,G37371,G37372,G37373,G37374,G37375,G37376,G37377,G37378,G37379,G37380,
       G37381,G37382,G37383,G37384,G37385,G37386,G37387,G37388,G37389,G37390,G37391,G37392,G37393,G37394,G37395,G37396,G37397,G37398,G37399,G37400,
       G37401,G37402,G37403,G37404,G37405,G37406,G37407,G37408,G37409,G37410,G37411,G37412,G37413,G37414,G37415,G37416,G37417,G37418,G37419,G37420,
       G37421,G37422,G37423,G37424,G37425,G37426,G37427,G37428,G37429,G37430,G37431,G37432,G37433,G37434,G37435,G37436,G37437,G37438,G37439,G37440,
       G37441,G37442,G37443,G37444,G37445,G37446,G37447,G37448,G37449,G37450,G37451,G37452,G37453,G37454,G37455,G37456,G37457,G37458,G37459,G37460,
       G37461,G37462,G37463,G37464,G37465,G37466,G37467,G37468,G37469,G37470,G37471,G37472,G37473,G37474,G37475,G37476,G37477,G37478,G37479,G37480,
       G37481,G37482,G37483,G37484,G37485,G37486,G37487,G37488,G37489,G37490,G37491,G37492,G37493,G37494,G37495,G37496,G37497,G37498,G37499,G37500,
       G37501,G37502,G37503,G37504,G37505,G37506,G37507,G37508,G37509,G37510,G37511,G37512,G37513,G37514,G37515,G37516,G37517,G37518,G37519,G37520,
       G37521,G37522,G37523,G37524,G37525,G37526,G37527,G37528,G37529,G37530,G37531,G37532,G37533,G37534,G37535,G37536,G37537,G37538,G37539,G37540,
       G37541,G37542,G37543,G37544,G37545,G37546,G37547,G37548,G37549,G37550,G37551,G37552,G37553,G37554,G37555,G37556,G37557,G37558,G37559,G37560,
       G37561,G37562,G37563,G37564,G37565,G37566,G37567,G37568,G37569,G37570,G37571,G37572,G37573,G37574,G37575,G37576,G37577,G37578,G37579,G37580,
       G37581,G37582,G37583,G37584,G37585,G37586,G37587,G37588,G37589,G37590,G37591,G37592,G37593,G37594,G37595,G37596,G37597,G37598,G37599,G37600,
       G37601,G37602,G37603,G37604,G37605,G37606,G37607,G37608,G37609,G37610,G37611,G37612,G37613,G37614,G37615,G37616,G37617,G37618,G37619,G37620,
       G37621,G37622,G37623,G37624,G37625,G37626,G37627,G37628,G37629,G37630,G37631,G37632,G37633,G37634,G37635,G37636,G37637,G37638,G37639,G37640,
       G37641,G37642,G37643,G37644,G37645,G37646,G37647,G37648,G37649,G37650,G37651,G37652,G37653,G37654,G37655,G37656,G37657,G37658,G37659,G37660,
       G37661,G37662,G37663,G37664,G37665,G37666,G37667,G37668,G37669,G37670,G37671,G37672,G37673,G37674,G37675,G37676,G37677,G37678,G37679,G37680,
       G37681,G37682,G37683,G37684,G37685,G37686,G37687,G37688,G37689,G37690,G37691,G37692,G37693,G37694,G37695,G37696,G37697,G37698,G37699,G37700,
       G37701,G37702,G37703,G37704,G37705,G37706,G37707,G37708,G37709,G37710,G37711,G37712,G37713,G37714,G37715,G37716,G37717,G37718,G37719,G37720,
       G37721,G37722,G37723,G37724,G37725,G37726,G37727,G37728,G37729,G37730,G37731,G37732,G37733,G37734,G37735,G37736,G37737,G37738,G37739,G37740,
       G37741,G37742,G37743,G37744,G37745,G37746,G37747,G37748,G37749,G37750,G37751,G37752,G37753,G37754,G37755,G37756,G37757,G37758,G37759,G37760,
       G37761,G37762,G37763,G37764,G37765,G37766,G37767,G37768,G37769,G37770,G37771,G37772,G37773,G37774,G37775,G37776,G37777,G37778,G37779,G37780,
       G37781,G37782,G37783,G37784,G37785,G37786,G37787,G37788,G37789,G37790,G37791,G37792,G37793,G37794,G37795,G37796,G37797,G37798,G37799,G37800,
       G37801,G37802,G37803,G37804,G37805,G37806,G37807,G37808,G37809,G37810,G37811,G37812,G37813,G37814,G37815,G37816,G37817,G37818,G37819,G37820,
       G37821,G37822,G37823,G37824,G37825,G37826,G37827,G37828,G37829,G37830,G37831,G37832,G37833,G37834,G37835,G37836,G37837,G37838,G37839,G37840,
       G37841,G37842,G37843,G37844,G37845,G37846,G37847,G37848,G37849,G37850,G37851,G37852,G37853,G37854,G37855,G37856,G37857,G37858,G37859,G37860,
       G37861,G37862,G37863,G37864,G37865,G37866,G37867,G37868,G37869,G37870,G37871,G37872,G37873,G37874,G37875,G37876,G37877,G37878,G37879,G37880,
       G37881,G37882,G37883,G37884,G37885,G37886,G37887,G37888,G37889,G37890,G37891,G37892,G37893,G37894,G37895,G37896,G37897,G37898,G37899,G37900,
       G37901,G37902,G37903,G37904,G37905,G37906,G37907,G37908,G37909,G37910,G37911,G37912,G37913,G37914,G37915,G37916,G37917,G37918,G37919,G37920,
       G37921,G37922,G37923,G37924,G37925,G37926,G37927,G37928,G37929,G37930,G37931,G37932,G37933,G37934,G37935,G37936,G37937,G37938,G37939,G37940,
       G37941,G37942,G37943,G37944,G37945,G37946,G37947,G37948,G37949,G37950,G37951,G37952,G37953,G37954,G37955,G37956,G37957,G37958,G37959,G37960,
       G37961,G37962,G37963,G37964,G37965,G37966,G37967,G37968,G37969,G37970,G37971,G37972,G37973,G37974,G37975,G37976,G37977,G37978,G37979,G37980,
       G37981,G37982,G37983,G37984,G37985,G37986,G37987,G37988,G37989,G37990,G37991,G37992,G37993,G37994,G37995,G37996,G37997,G37998,G37999,G38000,
       G38001,G38002,G38003,G38004,G38005,G38006,G38007,G38008,G38009,G38010,G38011,G38012,G38013,G38014,G38015,G38016,G38017,G38018,G38019,G38020,
       G38021,G38022,G38023,G38024,G38025,G38026,G38027,G38028,G38029,G38030,G38031,G38032,G38033,G38034,G38035,G38036,G38037,G38038,G38039,G38040,
       G38041,G38042,G38043,G38044,G38045,G38046,G38047,G38048,G38049,G38050,G38051,G38052,G38053,G38054,G38055,G38056,G38057,G38058,G38059,G38060,
       G38061,G38062,G38063,G38064,G38065,G38066,G38067,G38068,G38069,G38070,G38071,G38072,G38073,G38074,G38075,G38076,G38077,G38078,G38079,G38080,
       G38081,G38082,G38083,G38084,G38085,G38086,G38087,G38088,G38089,G38090,G38091,G38092,G38093,G38094,G38095,G38096,G38097,G38098,G38099,G38100,
       G38101,G38102,G38103,G38104,G38105,G38106,G38107,G38108,G38109,G38110,G38111,G38112,G38113,G38114,G38115,G38116,G38117,G38118,G38119,G38120,
       G38121,G38122,G38123,G38124,G38125,G38126,G38127,G38128,G38129,G38130,G38131,G38132,G38133,G38134,G38135,G38136,G38137,G38138,G38139,G38140,
       G38141,G38142,G38143,G38144,G38145,G38146,G38147,G38148,G38149,G38150,G38151,G38152,G38153,G38154,G38155,G38156,G38157,G38158,G38159,G38160,
       G38161,G38162,G38163,G38164,G38165,G38166,G38167,G38168,G38169,G38170,G38171,G38172,G38173,G38174,G38175,G38176,G38177,G38178,G38179,G38180,
       G38181,G38182,G38183,G38184,G38185,G38186,G38187,G38188,G38189,G38190,G38191,G38192,G38193,G38194,G38195,G38196,G38197,G38198,G38199,G38200,
       G38201,G38202,G38203,G38204,G38205,G38206,G38207,G38208,G38209,G38210,G38211,G38212,G38213,G38214,G38215,G38216,G38217,G38218,G38219,G38220,
       G38221,G38222,G38223,G38224,G38225,G38226,G38227,G38228,G38229,G38230,G38231,G38232,G38233,G38234,G38235,G38236,G38237,G38238,G38239,G38240,
       G38241,G38242,G38243,G38244,G38245,G38246,G38247,G38248,G38249,G38250,G38251,G38252,G38253,G38254,G38255,G38256,G38257,G38258,G38259,G38260,
       G38261,G38262,G38263,G38264,G38265,G38266,G38267,G38268,G38269,G38270,G38271,G38272,G38273,G38274,G38275,G38276,G38277,G38278,G38279,G38280,
       G38281,G38282,G38283,G38284,G38285,G38286,G38287,G38288,G38289,G38290,G38291,G38292,G38293,G38294,G38295,G38296,G38297,G38298,G38299,G38300,
       G38301,G38302,G38303,G38304,G38305,G38306,G38307,G38308,G38309,G38310,G38311,G38312,G38313,G38314,G38315,G38316,G38317,G38318,G38319,G38320,
       G38321,G38322,G38323,G38324,G38325,G38326,G38327,G38328,G38329,G38330,G38331,G38332,G38333,G38334,G38335,G38336,G38337,G38338,G38339,G38340,
       G38341,G38342,G38343,G38344,G38345,G38346,G38347,G38348,G38349,G38350,G38351,G38352,G38353,G38354,G38355,G38356,G38357,G38358,G38359,G38360,
       G38361,G38362,G38363,G38364,G38365,G38366,G38367,G38368,G38369,G38370,G38371,G38372,G38373,G38374,G38375,G38376,G38377,G38378,G38379,G38380,
       G38381,G38382,G38383,G38384,G38385,G38386,G38387,G38388,G38389,G38390,G38391,G38392,G38393,G38394,G38395,G38396,G38397,G38398,G38399,G38400,
       G38401,G38402,G38403,G38404,G38405,G38406,G38407,G38408,G38409,G38410,G38411,G38412,G38413,G38414,G38415,G38416,G38417,G38418,G38419,G38420,
       G38421,G38422,G38423,G38424,G38425,G38426,G38427,G38428,G38429,G38430,G38431,G38432,G38433,G38434,G38435,G38436,G38437,G38438,G38439,G38440,
       G38441,G38442,G38443,G38444,G38445,G38446,G38447,G38448,G38449,G38450,G38451,G38452,G38453,G38454,G38455,G38456,G38457,G38458,G38459,G38460,
       G38461,G38462,G38463,G38464,G38465,G38466,G38467,G38468,G38469,G38470,G38471,G38472,G38473,G38474,G38475,G38476,G38477,G38478,G38479,G38480,
       G38481,G38482,G38483,G38484,G38485,G38486,G38487,G38488,G38489,G38490,G38491,G38492,G38493,G38494,G38495,G38496,G38497,G38498,G38499,G38500,
       G38501,G38502,G38503,G38504,G38505,G38506,G38507,G38508,G38509,G38510,G38511,G38512,G38513,G38514,G38515,G38516,G38517,G38518,G38519,G38520,
       G38521,G38522,G38523,G38524,G38525,G38526,G38527,G38528,G38529,G38530,G38531,G38532,G38533,G38534,G38535,G38536,G38537,G38538,G38539,G38540,
       G38541,G38542,G38543,G38544,G38545,G38546,G38547,G38548,G38549,G38550,G38551,G38552,G38553,G38554,G38555,G38556,G38557,G38558,G38559,G38560,
       G38561,G38562,G38563,G38564,G38565,G38566,G38567,G38568,G38569,G38570,G38571,G38572,G38573,G38574,G38575,G38576,G38577,G38578,G38579,G38580,
       G38581,G38582,G38583,G38584,G38585,G38586,G38587,G38588,G38589,G38590,G38591,G38592,G38593,G38594,G38595,G38596,G38597,G38598,G38599,G38600,
       G38601,G38602,G38603,G38604,G38605,G38606,G38607,G38608,G38609,G38610,G38611,G38612,G38613,G38614,G38615,G38616,G38617,G38618,G38619,G38620,
       G38621,G38622,G38623,G38624,G38625,G38626,G38627,G38628,G38629,G38630,G38631,G38632,G38633,G38634,G38635,G38636,G38637,G38638,G38639,G38640,
       G38641,G38642,G38643,G38644,G38645,G38646,G38647,G38648,G38649,G38650,G38651,G38652,G38653,G38654,G38655,G38656,G38657,G38658,G38659,G38660,
       G38661,G38662,G38663,G38664,G38665,G38666,G38667,G38668,G38669,G38670,G38671,G38672,G38673,G38674,G38675,G38676,G38677,G38678,G38679,G38680,
       G38681,G38682,G38683,G38684,G38685,G38686,G38687,G38688,G38689,G38690,G38691,G38692,G38693,G38694,G38695,G38696,G38697,G38698,G38699,G38700,
       G38701,G38702,G38703,G38704,G38705,G38706,G38707,G38708,G38709,G38710,G38711,G38712,G38713,G38714,G38715,G38716,G38717,G38718,G38719,G38720,
       G38721,G38722,G38723,G38724,G38725,G38726,G38727,G38728,G38729,G38730,G38731,G38732,G38733,G38734,G38735,G38736,G38737,G38738,G38739,G38740,
       G38741,G38742,G38743,G38744,G38745,G38746,G38747,G38748,G38749,G38750,G38751,G38752,G38753,G38754,G38755,G38756,G38757,G38758,G38759,G38760,
       G38761,G38762,G38763,G38764,G38765,G38766,G38767,G38768,G38769,G38770,G38771,G38772,G38773,G38774,G38775,G38776,G38777,G38778,G38779,G38780,
       G38781,G38782,G38783,G38784,G38785,G38786,G38787,G38788,G38789,G38790,G38791,G38792,G38793,G38794,G38795,G38796,G38797,G38798,G38799,G38800,
       G38801,G38802,G38803,G38804,G38805,G38806,G38807,G38808,G38809,G38810,G38811,G38812,G38813,G38814,G38815,G38816,G38817,G38818,G38819,G38820,
       G38821,G38822,G38823,G38824,G38825,G38826,G38827,G38828,G38829,G38830,G38831,G38832,G38833,G38834,G38835,G38836,G38837,G38838,G38839,G38840,
       G38841,G38842,G38843,G38844,G38845,G38846,G38847,G38848,G38849,G38850,G38851,G38852,G38853,G38854,G38855,G38856,G38857,G38858,G38859,G38860,
       G38861,G38862,G38863,G38864,G38865,G38866,G38867,G38868,G38869,G38870,G38871,G38872,G38873,G38874,G38875,G38876,G38877,G38878,G38879,G38880,
       G38881,G38882,G38883,G38884,G38885,G38886,G38887,G38888,G38889,G38890,G38891,G38892,G38893,G38894,G38895,G38896,G38897,G38898,G38899,G38900,
       G38901,G38902,G38903,G38904,G38905,G38906,G38907,G38908,G38909,G38910,G38911,G38912,G38913,G38914,G38915,G38916,G38917,G38918,G38919,G38920,
       G38921,G38922,G38923,G38924,G38925,G38926,G38927,G38928,G38929,G38930,G38931,G38932,G38933,G38934,G38935,G38936,G38937,G38938,G38939,G38940,
       G38941,G38942,G38943,G38944,G38945,G38946,G38947,G38948,G38949,G38950,G38951,G38952,G38953,G38954,G38955,G38956,G38957,G38958,G38959,G38960,
       G38961,G38962,G38963,G38964,G38965,G38966,G38967,G38968,G38969,G38970,G38971,G38972,G38973,G38974,G38975,G38976,G38977,G38978,G38979,G38980,
       G38981,G38982,G38983,G38984,G38985,G38986,G38987,G38988,G38989,G38990,G38991,G38992,G38993,G38994,G38995,G38996,G38997,G38998,G38999,G39000,
       G39001,G39002,G39003,G39004,G39005,G39006,G39007,G39008,G39009,G39010,G39011,G39012,G39013,G39014,G39015,G39016,G39017,G39018,G39019,G39020,
       G39021,G39022,G39023,G39024,G39025,G39026,G39027,G39028,G39029,G39030,G39031,G39032,G39033,G39034,G39035,G39036,G39037,G39038,G39039,G39040,
       G39041,G39042,G39043,G39044,G39045,G39046,G39047,G39048,G39049,G39050,G39051,G39052,G39053,G39054,G39055,G39056,G39057,G39058,G39059,G39060,
       G39061,G39062,G39063,G39064,G39065,G39066,G39067,G39068,G39069,G39070,G39071,G39072,G39073,G39074,G39075,G39076,G39077,G39078,G39079,G39080,
       G39081,G39082,G39083,G39084,G39085,G39086,G39087,G39088,G39089,G39090,G39091,G39092,G39093,G39094,G39095,G39096,G39097,G39098,G39099,G39100,
       G39101,G39102,G39103,G39104,G39105,G39106,G39107,G39108,G39109,G39110,G39111,G39112,G39113,G39114,G39115,G39116,G39117,G39118,G39119,G39120,
       G39121,G39122,G39123,G39124,G39125,G39126,G39127,G39128,G39129,G39130,G39131,G39132,G39133,G39134,G39135,G39136,G39137,G39138,G39139,G39140,
       G39141,G39142,G39143,G39144,G39145,G39146,G39147,G39148,G39149,G39150,G39151,G39152,G39153,G39154,G39155,G39156,G39157,G39158,G39159,G39160,
       G39161,G39162,G39163,G39164,G39165,G39166,G39167,G39168,G39169,G39170,G39171,G39172,G39173,G39174,G39175,G39176,G39177,G39178,G39179,G39180,
       G39181,G39182,G39183,G39184,G39185,G39186,G39187,G39188,G39189,G39190,G39191,G39192,G39193,G39194,G39195,G39196,G39197,G39198,G39199,G39200,
       G39201,G39202,G39203,G39204,G39205,G39206,G39207,G39208,G39209,G39210,G39211,G39212,G39213,G39214,G39215,G39216,G39217,G39218,G39219,G39220,
       G39221,G39222,G39223,G39224,G39225,G39226,G39227,G39228,G39229,G39230,G39231,G39232,G39233,G39234,G39235,G39236,G39237,G39238,G39239,G39240,
       G39241,G39242,G39243,G39244,G39245,G39246,G39247,G39248,G39249,G39250,G39251,G39252,G39253,G39254,G39255,G39256,G39257,G39258,G39259,G39260,
       G39261,G39262,G39263,G39264,G39265,G39266,G39267,G39268,G39269,G39270,G39271,G39272,G39273,G39274,G39275,G39276,G39277,G39278,G39279,G39280,
       G39281,G39282,G39283,G39284,G39285,G39286,G39287,G39288,G39289,G39290,G39291,G39292,G39293,G39294,G39295,G39296,G39297,G39298,G39299,G39300,
       G39301,G39302,G39303,G39304,G39305,G39306,G39307,G39308,G39309,G39310,G39311,G39312,G39313,G39314,G39315,G39316,G39317,G39318,G39319,G39320,
       G39321,G39322,G39323,G39324,G39325,G39326,G39327,G39328,G39329,G39330,G39331,G39332,G39333,G39334,G39335,G39336,G39337,G39338,G39339,G39340,
       G39341,G39342,G39343,G39344,G39345,G39346,G39347,G39348,G39349,G39350,G39351,G39352,G39353,G39354,G39355,G39356,G39357,G39358,G39359,G39360,
       G39361,G39362,G39363,G39364,G39365,G39366,G39367,G39368,G39369,G39370,G39371,G39372,G39373,G39374,G39375,G39376,G39377,G39378,G39379,G39380,
       G39381,G39382,G39383,G39384,G39385,G39386,G39387,G39388,G39389,G39390,G39391,G39392,G39393,G39394,G39395,G39396,G39397,G39398,G39399,G39400,
       G39401,G39402,G39403,G39404,G39405,G39406,G39407,G39408,G39409,G39410,G39411,G39412,G39413,G39414,G39415,G39416,G39417,G39418,G39419,G39420,
       G39421,G39422,G39423,G39424,G39425,G39426,G39427,G39428,G39429,G39430,G39431,G39432,G39433,G39434,G39435,G39436,G39437,G39438,G39439,G39440,
       G39441,G39442,G39443,G39444,G39445,G39446,G39447,G39448,G39449,G39450,G39451,G39452,G39453,G39454,G39455,G39456,G39457,G39458,G39459,G39460,
       G39461,G39462,G39463,G39464,G39465,G39466,G39467,G39468,G39469,G39470,G39471,G39472,G39473,G39474,G39475,G39476,G39477,G39478,G39479,G39480,
       G39481,G39482,G39483,G39484,G39485,G39486,G39487,G39488,G39489,G39490,G39491,G39492,G39493,G39494,G39495,G39496,G39497,G39498,G39499,G39500,
       G39501,G39502,G39503,G39504,G39505,G39506,G39507,G39508,G39509,G39510,G39511,G39512,G39513,G39514,G39515,G39516,G39517,G39518,G39519,G39520,
       G39521,G39522,G39523,G39524,G39525,G39526,G39527,G39528,G39529,G39530,G39531,G39532,G39533,G39534,G39535,G39536,G39537,G39538,G39539,G39540,
       G39541,G39542,G39543,G39544,G39545,G39546,G39547,G39548,G39549,G39550,G39551,G39552,G39553,G39554,G39555,G39556,G39557,G39558,G39559,G39560,
       G39561,G39562,G39563,G39564,G39565,G39566,G39567,G39568,G39569,G39570,G39571,G39572,G39573,G39574,G39575,G39576,G39577,G39578,G39579,G39580,
       G39581,G39582,G39583,G39584,G39585,G39586,G39587,G39588,G39589,G39590,G39591,G39592,G39593,G39594,G39595,G39596,G39597,G39598,G39599,G39600,
       G39601,G39602,G39603,G39604,G39605,G39606,G39607,G39608,G39609,G39610,G39611,G39612,G39613,G39614,G39615,G39616,G39617,G39618,G39619,G39620,
       G39621,G39622,G39623,G39624,G39625,G39626,G39627,G39628,G39629,G39630,G39631,G39632,G39633,G39634,G39635,G39636,G39637,G39638,G39639,G39640,
       G39641,G39642,G39643,G39644,G39645,G39646,G39647,G39648,G39649,G39650,G39651,G39652,G39653,G39654,G39655,G39656,G39657,G39658,G39659,G39660,
       G39661,G39662,G39663,G39664,G39665,G39666,G39667,G39668,G39669,G39670,G39671,G39672,G39673,G39674,G39675,G39676,G39677,G39678,G39679,G39680,
       G39681,G39682,G39683,G39684,G39685,G39686,G39687,G39688,G39689,G39690,G39691,G39692,G39693,G39694,G39695,G39696,G39697,G39698,G39699,G39700,
       G39701,G39702,G39703,G39704,G39705,G39706,G39707,G39708,G39709,G39710,G39711,G39712,G39713,G39714,G39715,G39716,G39717,G39718,G39719,G39720,
       G39721,G39722,G39723,G39724,G39725,G39726,G39727,G39728,G39729,G39730,G39731,G39732,G39733,G39734,G39735,G39736,G39737,G39738,G39739,G39740,
       G39741,G39742,G39743,G39744,G39745,G39746,G39747,G39748,G39749,G39750,G39751,G39752,G39753,G39754,G39755,G39756,G39757,G39758,G39759,G39760,
       G39761,G39762,G39763,G39764,G39765,G39766,G39767,G39768,G39769,G39770,G39771,G39772,G39773,G39774,G39775,G39776,G39777,G39778,G39779,G39780,
       G39781,G39782,G39783,G39784,G39785,G39786,G39787,G39788,G39789,G39790,G39791,G39792,G39793,G39794,G39795,G39796,G39797,G39798,G39799,G39800,
       G39801,G39802,G39803,G39804,G39805,G39806,G39807,G39808,G39809,G39810,G39811,G39812,G39813,G39814,G39815,G39816,G39817,G39818,G39819,G39820,
       G39821,G39822,G39823,G39824,G39825,G39826,G39827,G39828,G39829,G39830,G39831,G39832,G39833,G39834,G39835,G39836,G39837,G39838,G39839,G39840,
       G39841,G39842,G39843,G39844,G39845,G39846,G39847,G39848,G39849,G39850,G39851,G39852,G39853,G39854,G39855,G39856,G39857,G39858,G39859,G39860,
       G39861,G39862,G39863,G39864,G39865,G39866,G39867,G39868,G39869,G39870,G39871,G39872,G39873,G39874,G39875,G39876,G39877,G39878,G39879,G39880,
       G39881,G39882,G39883,G39884,G39885,G39886,G39887,G39888,G39889,G39890,G39891,G39892,G39893,G39894,G39895,G39896,G39897,G39898,G39899,G39900,
       G39901,G39902,G39903,G39904,G39905,G39906,G39907,G39908,G39909,G39910,G39911,G39912,G39913,G39914,G39915,G39916,G39917,G39918,G39919,G39920,
       G39921,G39922,G39923,G39924,G39925,G39926,G39927,G39928,G39929,G39930,G39931,G39932,G39933,G39934,G39935,G39936,G39937,G39938,G39939,G39940,
       G39941,G39942,G39943,G39944,G39945,G39946,G39947,G39948,G39949,G39950,G39951,G39952,G39953,G39954,G39955,G39956,G39957,G39958,G39959,G39960,
       G39961,G39962,G39963,G39964,G39965,G39966,G39967,G39968,G39969,G39970,G39971,G39972,G39973,G39974,G39975,G39976,G39977,G39978,G39979,G39980,
       G39981,G39982,G39983,G39984,G39985,G39986,G39987,G39988,G39989,G39990,G39991,G39992,G39993,G39994,G39995,G39996,G39997,G39998,G39999,G40000,
       G40001,G40002,G40003,G40004,G40005,G40006,G40007,G40008,G40009,G40010,G40011,G40012,G40013,G40014,G40015,G40016,G40017,G40018,G40019,G40020,
       G40021,G40022,G40023,G40024,G40025,G40026,G40027,G40028,G40029,G40030,G40031,G40032,G40033,G40034,G40035,G40036,G40037,G40038,G40039,G40040,
       G40041,G40042,G40043,G40044,G40045,G40046,G40047,G40048,G40049,G40050,G40051,G40052,G40053,G40054,G40055,G40056,G40057,G40058,G40059,G40060,
       G40061,G40062,G40063,G40064,G40065,G40066,G40067,G40068,G40069,G40070,G40071,G40072,G40073,G40074,G40075,G40076,G40077,G40078,G40079,G40080,
       G40081,G40082,G40083,G40084,G40085,G40086,G40087,G40088,G40089,G40090,G40091,G40092,G40093,G40094,G40095,G40096,G40097,G40098,G40099,G40100,
       G40101,G40102,G40103,G40104,G40105,G40106,G40107,G40108,G40109,G40110,G40111,G40112,G40113,G40114,G40115,G40116,G40117,G40118,G40119,G40120,
       G40121,G40122,G40123,G40124,G40125,G40126,G40127,G40128,G40129,G40130,G40131,G40132,G40133,G40134,G40135,G40136,G40137,G40138,G40139,G40140,
       G40141,G40142,G40143,G40144,G40145,G40146,G40147,G40148,G40149,G40150,G40151,G40152,G40153,G40154,G40155,G40156,G40157,G40158,G40159,G40160,
       G40161,G40162,G40163,G40164,G40165,G40166,G40167,G40168,G40169,G40170,G40171,G40172,G40173,G40174,G40175,G40176,G40177,G40178,G40179,G40180,
       G40181,G40182,G40183,G40184,G40185,G40186,G40187,G40188,G40189,G40190,G40191,G40192,G40193,G40194,G40195,G40196,G40197,G40198,G40199,G40200,
       G40201,G40202,G40203,G40204,G40205,G40206,G40207,G40208,G40209,G40210,G40211,G40212,G40213,G40214,G40215,G40216,G40217,G40218,G40219,G40220,
       G40221,G40222,G40223,G40224,G40225,G40226,G40227,G40228,G40229,G40230,G40231,G40232,G40233,G40234,G40235,G40236,G40237,G40238,G40239,G40240,
       G40241,G40242,G40243,G40244,G40245,G40246,G40247,G40248,G40249,G40250,G40251,G40252,G40253,G40254,G40255,G40256,G40257,G40258,G40259,G40260,
       G40261,G40262,G40263,G40264,G40265,G40266,G40267,G40268,G40269,G40270,G40271,G40272,G40273,G40274,G40275,G40276,G40277,G40278,G40279,G40280,
       G40281,G40282,G40283,G40284,G40285,G40286,G40287,G40288,G40289,G40290,G40291,G40292,G40293,G40294,G40295,G40296,G40297,G40298,G40299,G40300,
       G40301,G40302,G40303,G40304,G40305,G40306,G40307,G40308,G40309,G40310,G40311,G40312,G40313,G40314,G40315,G40316,G40317,G40318,G40319,G40320,
       G40321,G40322,G40323,G40324,G40325,G40326,G40327,G40328,G40329,G40330,G40331,G40332,G40333,G40334,G40335,G40336,G40337,G40338,G40339,G40340,
       G40341,G40342,G40343,G40344,G40345,G40346,G40347,G40348,G40349,G40350,G40351,G40352,G40353,G40354,G40355,G40356,G40357,G40358,G40359,G40360,
       G40361,G40362,G40363,G40364,G40365,G40366,G40367,G40368,G40369,G40370,G40371,G40372,G40373,G40374,G40375,G40376,G40377,G40378,G40379,G40380,
       G40381,G40382,G40383,G40384,G40385,G40386,G40387,G40388,G40389,G40390,G40391,G40392,G40393,G40394,G40395,G40396,G40397,G40398,G40399,G40400,
       G40401,G40402,G40403,G40404,G40405,G40406,G40407,G40408,G40409,G40410,G40411,G40412,G40413,G40414,G40415,G40416,G40417,G40418,G40419,G40420,
       G40421,G40422,G40423,G40424,G40425,G40426,G40427,G40428,G40429,G40430,G40431,G40432,G40433,G40434,G40435,G40436,G40437,G40438,G40439,G40440,
       G40441,G40442,G40443,G40444,G40445,G40446,G40447,G40448,G40449,G40450,G40451,G40452,G40453,G40454,G40455,G40456,G40457,G40458,G40459,G40460,
       G40461,G40462,G40463,G40464,G40465,G40466,G40467,G40468,G40469,G40470,G40471,G40472,G40473,G40474,G40475,G40476,G40477,G40478,G40479,G40480,
       G40481,G40482,G40483,G40484,G40485,G40486,G40487,G40488,G40489,G40490,G40491,G40492,G40493,G40494,G40495,G40496,G40497,G40498,G40499,G40500,
       G40501,G40502,G40503,G40504,G40505,G40506,G40507,G40508,G40509,G40510,G40511,G40512,G40513,G40514,G40515,G40516,G40517,G40518,G40519,G40520,
       G40521,G40522,G40523,G40524,G40525,G40526,G40527,G40528,G40529,G40530,G40531,G40532,G40533,G40534,G40535,G40536,G40537,G40538,G40539,G40540,
       G40541,G40542,G40543,G40544,G40545,G40546,G40547,G40548,G40549,G40550,G40551,G40552,G40553,G40554,G40555,G40556,G40557,G40558,G40559,G40560,
       G40561,G40562,G40563,G40564,G40565,G40566,G40567,G40568,G40569,G40570,G40571,G40572,G40573,G40574,G40575,G40576,G40577,G40578,G40579,G40580,
       G40581,G40582,G40583,G40584,G40585,G40586,G40587,G40588,G40589,G40590,G40591,G40592,G40593,G40594,G40595,G40596,G40597,G40598,G40599,G40600,
       G40601,G40602,G40603,G40604,G40605,G40606,G40607,G40608,G40609,G40610,G40611,G40612,G40613,G40614,G40615,G40616,G40617,G40618,G40619,G40620,
       G40621,G40622,G40623,G40624,G40625,G40626,G40627,G40628,G40629,G40630,G40631,G40632,G40633,G40634,G40635,G40636,G40637,G40638,G40639,G40640,
       G40641,G40642,G40643,G40644,G40645,G40646,G40647,G40648,G40649,G40650,G40651,G40652,G40653,G40654,G40655,G40656,G40657,G40658,G40659,G40660,
       G40661,G40662,G40663,G40664,G40665,G40666,G40667,G40668,G40669,G40670,G40671,G40672,G40673,G40674,G40675,G40676,G40677,G40678,G40679,G40680,
       G40681,G40682,G40683,G40684,G40685,G40686,G40687,G40688,G40689,G40690,G40691,G40692,G40693,G40694,G40695,G40696,G40697,G40698,G40699,G40700,
       G40701,G40702,G40703,G40704,G40705,G40706,G40707,G40708,G40709,G40710,G40711,G40712,G40713,G40714,G40715,G40716,G40717,G40718,G40719,G40720,
       G40721,G40722,G40723,G40724,G40725,G40726,G40727,G40728,G40729,G40730,G40731,G40732,G40733,G40734,G40735,G40736,G40737,G40738,G40739,G40740,
       G40741,G40742,G40743,G40744,G40745,G40746,G40747,G40748,G40749,G40750,G40751,G40752,G40753,G40754,G40755,G40756,G40757,G40758,G40759,G40760,
       G40761,G40762,G40763,G40764,G40765,G40766,G40767,G40768,G40769,G40770,G40771,G40772,G40773,G40774,G40775,G40776,G40777,G40778,G40779,G40780,
       G40781,G40782,G40783,G40784,G40785,G40786,G40787,G40788,G40789,G40790,G40791,G40792,G40793,G40794,G40795,G40796,G40797,G40798,G40799,G40800,
       G40801,G40802,G40803,G40804,G40805,G40806,G40807,G40808,G40809,G40810,G40811,G40812,G40813,G40814,G40815,G40816,G40817,G40818,G40819,G40820,
       G40821,G40822,G40823,G40824,G40825,G40826,G40827,G40828,G40829,G40830,G40831,G40832,G40833,G40834,G40835,G40836,G40837,G40838,G40839,G40840,
       G40841,G40842,G40843,G40844,G40845,G40846,G40847,G40848,G40849,G40850,G40851,G40852,G40853,G40854,G40855,G40856,G40857,G40858,G40859,G40860,
       G40861,G40862,G40863,G40864,G40865,G40866,G40867,G40868,G40869,G40870,G40871,G40872,G40873,G40874,G40875,G40876,G40877,G40878,G40879,G40880,
       G40881,G40882,G40883,G40884,G40885,G40886,G40887,G40888,G40889,G40890,G40891,G40892,G40893,G40894,G40895,G40896,G40897,G40898,G40899,G40900,
       G40901,G40902,G40903,G40904,G40905,G40906,G40907,G40908,G40909,G40910,G40911,G40912,G40913,G40914,G40915,G40916,G40917,G40918,G40919,G40920,
       G40921,G40922,G40923,G40924,G40925,G40926,G40927,G40928,G40929,G40930,G40931,G40932,G40933,G40934,G40935,G40936,G40937,G40938,G40939,G40940,
       G40941,G40942,G40943,G40944,G40945,G40946,G40947,G40948,G40949,G40950,G40951,G40952,G40953,G40954,G40955,G40956,G40957,G40958,G40959,G40960,
       G40961,G40962,G40963,G40964,G40965,G40966,G40967,G40968,G40969,G40970,G40971,G40972,G40973,G40974,G40975,G40976,G40977,G40978,G40979,G40980,
       G40981,G40982,G40983,G40984,G40985,G40986,G40987,G40988,G40989,G40990,G40991,G40992,G40993,G40994,G40995,G40996,G40997,G40998,G40999,G41000,
       G41001,G41002,G41003,G41004,G41005,G41006,G41007,G41008,G41009,G41010,G41011,G41012,G41013,G41014,G41015,G41016,G41017,G41018,G41019,G41020,
       G41021,G41022,G41023,G41024,G41025,G41026,G41027,G41028,G41029,G41030,G41031,G41032,G41033,G41034,G41035,G41036,G41037,G41038,G41039,G41040,
       G41041,G41042,G41043,G41044,G41045,G41046,G41047,G41048,G41049,G41050,G41051,G41052,G41053,G41054,G41055,G41056,G41057,G41058,G41059,G41060,
       G41061,G41062,G41063,G41064,G41065,G41066,G41067,G41068,G41069,G41070,G41071,G41072,G41073,G41074,G41075,G41076,G41077,G41078,G41079,G41080,
       G41081,G41082,G41083,G41084,G41085,G41086,G41087,G41088,G41089,G41090,G41091,G41092,G41093,G41094,G41095,G41096,G41097,G41098,G41099,G41100,
       G41101,G41102,G41103,G41104,G41105,G41106,G41107,G41108,G41109,G41110,G41111,G41112,G41113,G41114,G41115,G41116,G41117,G41118,G41119,G41120,
       G41121,G41122,G41123,G41124,G41125,G41126,G41127,G41128,G41129,G41130,G41131,G41132,G41133,G41134,G41135,G41136,G41137,G41138,G41139,G41140,
       G41141,G41142,G41143,G41144,G41145,G41146,G41147,G41148,G41149,G41150,G41151,G41152,G41153,G41154,G41155,G41156,G41157,G41158,G41159,G41160,
       G41161,G41162,G41163,G41164,G41165,G41166,G41167,G41168,G41169,G41170,G41171,G41172,G41173,G41174,G41175,G41176,G41177,G41178,G41179,G41180,
       G41181,G41182,G41183,G41184,G41185,G41186,G41187,G41188,G41189,G41190,G41191,G41192,G41193,G41194,G41195,G41196,G41197,G41198,G41199,G41200,
       G41201,G41202,G41203,G41204,G41205,G41206,G41207,G41208,G41209,G41210,G41211,G41212,G41213,G41214,G41215,G41216,G41217,G41218,G41219,G41220,
       G41221,G41222,G41223,G41224,G41225,G41226,G41227,G41228,G41229,G41230,G41231,G41232,G41233,G41234,G41235,G41236,G41237,G41238,G41239,G41240,
       G41241,G41242,G41243,G41244,G41245,G41246,G41247,G41248,G41249,G41250,G41251,G41252,G41253,G41254,G41255,G41256,G41257,G41258,G41259,G41260,
       G41261,G41262,G41263,G41264,G41265,G41266,G41267,G41268,G41269,G41270,G41271,G41272,G41273,G41274,G41275,G41276,G41277,G41278,G41279,G41280,
       G41281,G41282,G41283,G41284,G41285,G41286,G41287,G41288,G41289,G41290,G41291,G41292,G41293,G41294,G41295,G41296,G41297,G41298,G41299,G41300,
       G41301,G41302,G41303,G41304,G41305,G41306,G41307,G41308,G41309,G41310,G41311,G41312,G41313,G41314,G41315,G41316,G41317,G41318,G41319,G41320,
       G41321,G41322,G41323,G41324,G41325,G41326,G41327,G41328,G41329,G41330,G41331,G41332,G41333,G41334,G41335,G41336,G41337,G41338,G41339,G41340,
       G41341,G41342,G41343,G41344,G41345,G41346,G41347,G41348,G41349,G41350,G41351,G41352,G41353,G41354,G41355,G41356,G41357,G41358,G41359,G41360,
       G41361,G41362,G41363,G41364,G41365,G41366,G41367,G41368,G41369,G41370,G41371,G41372,G41373,G41374,G41375,G41376,G41377,G41378,G41379,G41380,
       G41381,G41382,G41383,G41384,G41385,G41386,G41387,G41388,G41389,G41390,G41391,G41392,G41393,G41394,G41395,G41396,G41397,G41398,G41399,G41400,
       G41401,G41402,G41403,G41404,G41405,G41406,G41407,G41408,G41409,G41410,G41411,G41412,G41413,G41414,G41415,G41416,G41417,G41418,G41419,G41420,
       G41421,G41422,G41423,G41424,G41425,G41426,G41427,G41428,G41429,G41430,G41431,G41432,G41433,G41434,G41435,G41436,G41437,G41438,G41439,G41440,
       G41441,G41442,G41443,G41444,G41445,G41446,G41447,G41448,G41449,G41450,G41451,G41452,G41453,G41454,G41455,G41456,G41457,G41458,G41459,G41460,
       G41461,G41462,G41463,G41464,G41465,G41466,G41467,G41468,G41469,G41470,G41471,G41472,G41473,G41474,G41475,G41476,G41477,G41478,G41479,G41480,
       G41481,G41482,G41483,G41484,G41485,G41486,G41487,G41488,G41489,G41490,G41491,G41492,G41493,G41494,G41495,G41496,G41497,G41498,G41499,G41500,
       G41501,G41502,G41503,G41504,G41505,G41506,G41507,G41508,G41509,G41510,G41511,G41512,G41513,G41514,G41515,G41516,G41517,G41518,G41519,G41520,
       G41521,G41522,G41523,G41524,G41525,G41526,G41527,G41528,G41529,G41530,G41531,G41532,G41533,G41534,G41535,G41536,G41537,G41538,G41539,G41540,
       G41541,G41542,G41543,G41544,G41545,G41546,G41547,G41548,G41549,G41550,G41551,G41552,G41553,G41554,G41555,G41556,G41557,G41558,G41559,G41560,
       G41561,G41562,G41563,G41564,G41565,G41566,G41567,G41568,G41569,G41570,G41571,G41572,G41573,G41574,G41575,G41576,G41577,G41578,G41579,G41580,
       G41581,G41582,G41583,G41584,G41585,G41586,G41587,G41588,G41589,G41590,G41591,G41592,G41593,G41594,G41595,G41596,G41597,G41598,G41599,G41600,
       G41601,G41602,G41603,G41604,G41605,G41606,G41607,G41608,G41609,G41610,G41611,G41612,G41613,G41614,G41615,G41616,G41617,G41618,G41619,G41620,
       G41621,G41622,G41623,G41624,G41625,G41626,G41627,G41628,G41629,G41630,G41631,G41632,G41633,G41634,G41635,G41636,G41637,G41638,G41639,G41640,
       G41641,G41642,G41643,G41644,G41645,G41646,G41647,G41648,G41649,G41650,G41651,G41652,G41653,G41654,G41655,G41656,G41657,G41658,G41659,G41660,
       G41661,G41662,G41663,G41664,G41665,G41666,G41667,G41668,G41669,G41670,G41671,G41672,G41673,G41674,G41675,G41676,G41677,G41678,G41679,G41680,
       G41681,G41682,G41683,G41684,G41685,G41686,G41687,G41688,G41689,G41690,G41691,G41692,G41693,G41694,G41695,G41696,G41697,G41698,G41699,G41700,
       G41701,G41702,G41703,G41704,G41705,G41706,G41707,G41708,G41709,G41710,G41711,G41712,G41713,G41714,G41715,G41716,G41717,G41718,G41719,G41720,
       G41721,G41722,G41723,G41724,G41725,G41726,G41727,G41728,G41729,G41730,G41731,G41732,G41733,G41734,G41735,G41736,G41737,G41738,G41739,G41740,
       G41741,G41742,G41743,G41744,G41745,G41746,G41747,G41748,G41749,G41750,G41751,G41752,G41753,G41754,G41755,G41756,G41757,G41758,G41759,G41760,
       G41761,G41762,G41763,G41764,G41765,G41766,G41767,G41768,G41769,G41770,G41771,G41772,G41773,G41774,G41775,G41776,G41777,G41778,G41779,G41780,
       G41781,G41782,G41783,G41784,G41785,G41786,G41787,G41788,G41789,G41790,G41791,G41792,G41793,G41794,G41795,G41796,G41797,G41798,G41799,G41800,
       G41801,G41802,G41803,G41804,G41805,G41806,G41807,G41808,G41809,G41810,G41811,G41812,G41813,G41814,G41815,G41816,G41817,G41818,G41819,G41820,
       G41821,G41822,G41823,G41824,G41825,G41826,G41827,G41828,G41829,G41830,G41831,G41832,G41833,G41834,G41835,G41836,G41837,G41838,G41839,G41840,
       G41841,G41842,G41843,G41844,G41845,G41846,G41847,G41848,G41849,G41850,G41851,G41852,G41853,G41854,G41855,G41856,G41857,G41858,G41859,G41860,
       G41861,G41862,G41863,G41864,G41865,G41866,G41867,G41868,G41869,G41870,G41871,G41872,G41873,G41874,G41875,G41876,G41877,G41878,G41879,G41880,
       G41881,G41882,G41883,G41884,G41885,G41886,G41887,G41888,G41889,G41890,G41891,G41892,G41893,G41894,G41895,G41896,G41897,G41898,G41899,G41900,
       G41901,G41902,G41903,G41904,G41905,G41906,G41907,G41908,G41909,G41910,G41911,G41912,G41913,G41914,G41915,G41916,G41917,G41918,G41919,G41920,
       G41921,G41922,G41923,G41924,G41925,G41926,G41927,G41928,G41929,G41930,G41931,G41932,G41933,G41934,G41935,G41936,G41937,G41938,G41939,G41940,
       G41941,G41942,G41943,G41944,G41945,G41946,G41947,G41948,G41949,G41950,G41951,G41952,G41953,G41954,G41955,G41956,G41957,G41958,G41959,G41960,
       G41961,G41962,G41963,G41964,G41965,G41966,G41967,G41968,G41969,G41970,G41971,G41972,G41973,G41974,G41975,G41976,G41977,G41978,G41979,G41980,
       G41981,G41982,G41983,G41984,G41985,G41986,G41987,G41988,G41989,G41990,G41991,G41992,G41993,G41994,G41995,G41996,G41997,G41998,G41999,G42000,
       G42001,G42002,G42003,G42004,G42005,G42006,G42007,G42008,G42009,G42010,G42011,G42012,G42013,G42014,G42015,G42016,G42017,G42018,G42019,G42020,
       G42021,G42022,G42023,G42024,G42025,G42026,G42027,G42028,G42029,G42030,G42031,G42032,G42033,G42034,G42035,G42036,G42037,G42038,G42039,G42040,
       G42041,G42042,G42043,G42044,G42045,G42046,G42047,G42048,G42049,G42050,G42051,G42052,G42053,G42054,G42055,G42056,G42057,G42058,G42059,G42060,
       G42061,G42062,G42063,G42064,G42065,G42066,G42067,G42068,G42069,G42070,G42071,G42072,G42073,G42074,G42075,G42076,G42077,G42078,G42079,G42080,
       G42081,G42082,G42083,G42084,G42085,G42086,G42087,G42088,G42089,G42090,G42091,G42092,G42093,G42094,G42095,G42096,G42097,G42098,G42099,G42100,
       G42101,G42102,G42103,G42104,G42105,G42106,G42107,G42108,G42109,G42110,G42111,G42112,G42113,G42114,G42115,G42116,G42117,G42118,G42119,G42120,
       G42121,G42122,G42123,G42124,G42125,G42126,G42127,G42128,G42129,G42130,G42131,G42132,G42133,G42134,G42135,G42136,G42137,G42138,G42139,G42140,
       G42141,G42142,G42143,G42144,G42145,G42146,G42147,G42148,G42149,G42150,G42151,G42152,G42153,G42154,G42155,G42156,G42157,G42158,G42159,G42160,
       G42161,G42162,G42163,G42164,G42165,G42166,G42167,G42168,G42169,G42170,G42171,G42172,G42173,G42174,G42175,G42176,G42177,G42178,G42179,G42180,
       G42181,G42182,G42183,G42184,G42185,G42186,G42187,G42188,G42189,G42190,G42191,G42192,G42193,G42194,G42195,G42196,G42197,G42198,G42199,G42200,
       G42201,G42202,G42203,G42204,G42205,G42206,G42207,G42208,G42209,G42210,G42211,G42212,G42213,G42214,G42215,G42216,G42217,G42218,G42219,G42220,
       G42221,G42222,G42223,G42224,G42225,G42226,G42227,G42228,G42229,G42230,G42231,G42232,G42233,G42234,G42235,G42236,G42237,G42238,G42239,G42240,
       G42241,G42242,G42243,G42244,G42245,G42246,G42247,G42248,G42249,G42250,G42251,G42252,G42253,G42254,G42255,G42256,G42257,G42258,G42259,G42260,
       G42261,G42262,G42263,G42264,G42265,G42266,G42267,G42268,G42269,G42270,G42271,G42272,G42273,G42274,G42275,G42276,G42277,G42278,G42279,G42280,
       G42281,G42282,G42283,G42284,G42285,G42286,G42287,G42288,G42289,G42290,G42291,G42292,G42293,G42294,G42295,G42296,G42297,G42298,G42299,G42300,
       G42301,G42302,G42303,G42304,G42305,G42306,G42307,G42308,G42309,G42310,G42311,G42312,G42313,G42314,G42315,G42316,G42317,G42318,G42319,G42320,
       G42321,G42322,G42323,G42324,G42325,G42326,G42327,G42328,G42329,G42330,G42331,G42332,G42333,G42334,G42335,G42336,G42337,G42338,G42339,G42340,
       G42341,G42342,G42343,G42344,G42345,G42346,G42347,G42348,G42349,G42350,G42351,G42352,G42353,G42354,G42355,G42356,G42357,G42358,G42359,G42360,
       G42361,G42362,G42363,G42364,G42365,G42366,G42367,G42368,G42369,G42370,G42371,G42372,G42373,G42374,G42375,G42376,G42377,G42378,G42379,G42380,
       G42381,G42382,G42383,G42384,G42385,G42386,G42387,G42388,G42389,G42390,G42391,G42392,G42393,G42394,G42395,G42396,G42397,G42398,G42399,G42400,
       G42401,G42402,G42403,G42404,G42405,G42406,G42407,G42408,G42409,G42410,G42411,G42412,G42413,G42414,G42415,G42416,G42417,G42418,G42419,G42420,
       G42421,G42422,G42423,G42424,G42425,G42426,G42427,G42428,G42429,G42430,G42431,G42432,G42433,G42434,G42435,G42436,G42437,G42438,G42439,G42440,
       G42441,G42442,G42443,G42444,G42445,G42446,G42447,G42448,G42449,G42450,G42451,G42452,G42453,G42454,G42455,G42456,G42457,G42458,G42459,G42460,
       G42461,G42462,G42463,G42464,G42465,G42466,G42467,G42468,G42469,G42470,G42471,G42472,G42473,G42474,G42475,G42476,G42477,G42478,G42479,G42480,
       G42481,G42482,G42483,G42484,G42485,G42486,G42487,G42488,G42489,G42490,G42491,G42492,G42493,G42494,G42495,G42496,G42497,G42498,G42499,G42500,
       G42501,G42502,G42503,G42504,G42505,G42506,G42507,G42508,G42509,G42510,G42511,G42512,G42513,G42514,G42515,G42516,G42517,G42518,G42519,G42520,
       G42521,G42522,G42523,G42524,G42525,G42526,G42527,G42528,G42529,G42530,G42531,G42532,G42533,G42534,G42535,G42536,G42537,G42538,G42539,G42540,
       G42541,G42542,G42543,G42544,G42545,G42546,G42547,G42548,G42549,G42550,G42551,G42552,G42553,G42554,G42555,G42556,G42557,G42558,G42559,G42560,
       G42561,G42562,G42563,G42564,G42565,G42566,G42567,G42568,G42569,G42570,G42571,G42572,G42573,G42574,G42575,G42576,G42577,G42578,G42579,G42580,
       G42581,G42582,G42583,G42584,G42585,G42586,G42587,G42588,G42589,G42590,G42591,G42592,G42593,G42594,G42595,G42596,G42597,G42598,G42599,G42600,
       G42601,G42602,G42603,G42604,G42605,G42606,G42607,G42608,G42609,G42610,G42611,G42612,G42613,G42614,G42615,G42616,G42617,G42618,G42619,G42620,
       G42621,G42622,G42623,G42624,G42625,G42626,G42627,G42628,G42629,G42630,G42631,G42632,G42633,G42634,G42635,G42636,G42637,G42638,G42639,G42640,
       G42641,G42642,G42643,G42644,G42645,G42646,G42647,G42648,G42649,G42650,G42651,G42652,G42653,G42654,G42655,G42656,G42657,G42658,G42659,G42660,
       G42661,G42662,G42663,G42664,G42665,G42666,G42667,G42668,G42669,G42670,G42671,G42672,G42673,G42674,G42675,G42676,G42677,G42678,G42679,G42680,
       G42681,G42682,G42683,G42684,G42685,G42686,G42687,G42688,G42689,G42690,G42691,G42692,G42693,G42694,G42695,G42696,G42697,G42698,G42699,G42700,
       G42701,G42702,G42703,G42704,G42705,G42706,G42707,G42708,G42709,G42710,G42711,G42712,G42713,G42714,G42715,G42716,G42717,G42718,G42719,G42720,
       G42721,G42722,G42723,G42724,G42725,G42726,G42727,G42728,G42729,G42730,G42731,G42732,G42733,G42734,G42735,G42736,G42737,G42738,G42739,G42740,
       G42741,G42742,G42743,G42744,G42745,G42746,G42747,G42748,G42749,G42750,G42751,G42752,G42753,G42754,G42755,G42756,G42757,G42758,G42759,G42760,
       G42761,G42762,G42763,G42764,G42765,G42766,G42767,G42768,G42769,G42770,G42771,G42772,G42773,G42774,G42775,G42776,G42777,G42778,G42779,G42780,
       G42781,G42782,G42783,G42784,G42785,G42786,G42787,G42788,G42789,G42790,G42791,G42792,G42793,G42794,G42795,G42796,G42797,G42798,G42799,G42800,
       G42801,G42802,G42803,G42804,G42805,G42806,G42807,G42808,G42809,G42810,G42811,G42812,G42813,G42814,G42815,G42816,G42817,G42818,G42819,G42820,
       G42821,G42822,G42823,G42824,G42825,G42826,G42827,G42828,G42829,G42830,G42831,G42832,G42833,G42834,G42835,G42836,G42837,G42838,G42839,G42840,
       G42841,G42842,G42843,G42844,G42845,G42846,G42847,G42848,G42849,G42850,G42851,G42852,G42853,G42854,G42855,G42856,G42857,G42858,G42859,G42860,
       G42861,G42862,G42863,G42864,G42865,G42866,G42867,G42868,G42869,G42870,G42871,G42872,G42873,G42874,G42875,G42876,G42877,G42878,G42879,G42880,
       G42881,G42882,G42883,G42884,G42885,G42886,G42887,G42888,G42889,G42890,G42891,G42892,G42893,G42894,G42895,G42896,G42897,G42898,G42899,G42900,
       G42901,G42902,G42903,G42904,G42905,G42906,G42907,G42908,G42909,G42910,G42911,G42912,G42913,G42914,G42915,G42916,G42917,G42918,G42919,G42920,
       G42921,G42922,G42923,G42924,G42925,G42926,G42927,G42928,G42929,G42930,G42931,G42932,G42933,G42934,G42935,G42936,G42937,G42938,G42939,G42940,
       G42941,G42942,G42943,G42944,G42945,G42946,G42947,G42948,G42949,G42950,G42951,G42952,G42953,G42954,G42955,G42956,G42957,G42958,G42959,G42960,
       G42961,G42962,G42963,G42964,G42965,G42966,G42967,G42968,G42969,G42970,G42971,G42972,G42973,G42974,G42975,G42976,G42977,G42978,G42979,G42980,
       G42981,G42982,G42983,G42984,G42985,G42986,G42987,G42988,G42989,G42990,G42991,G42992,G42993,G42994,G42995,G42996,G42997,G42998,G42999,G43000,
       G43001,G43002,G43003,G43004,G43005,G43006,G43007,G43008,G43009,G43010,G43011,G43012,G43013,G43014,G43015,G43016,G43017,G43018,G43019,G43020,
       G43021,G43022,G43023,G43024,G43025,G43026,G43027,G43028,G43029,G43030,G43031,G43032,G43033,G43034,G43035,G43036,G43037,G43038,G43039,G43040,
       G43041,G43042,G43043,G43044,G43045,G43046,G43047,G43048,G43049,G43050,G43051,G43052,G43053,G43054,G43055,G43056,G43057,G43058,G43059,G43060,
       G43061,G43062,G43063,G43064,G43065,G43066,G43067,G43068,G43069,G43070,G43071,G43072,G43073,G43074,G43075,G43076,G43077,G43078,G43079,G43080,
       G43081,G43082,G43083,G43084,G43085,G43086,G43087,G43088,G43089,G43090,G43091,G43092,G43093,G43094,G43095,G43096,G43097,G43098,G43099,G43100,
       G43101,G43102,G43103,G43104,G43105,G43106,G43107,G43108,G43109,G43110,G43111,G43112,G43113,G43114,G43115,G43116,G43117,G43118,G43119,G43120,
       G43121,G43122,G43123,G43124,G43125,G43126,G43127,G43128,G43129,G43130,G43131,G43132,G43133,G43134,G43135,G43136,G43137,G43138,G43139,G43140,
       G43141,G43142,G43143,G43144,G43145,G43146,G43147,G43148,G43149,G43150,G43151,G43152,G43153,G43154,G43155,G43156,G43157,G43158,G43159,G43160,
       G43161,G43162,G43163,G43164,G43165,G43166,G43167,G43168,G43169,G43170,G43171,G43172,G43173,G43174,G43175,G43176,G43177,G43178,G43179,G43180,
       G43181,G43182,G43183,G43184,G43185,G43186,G43187,G43188,G43189,G43190,G43191,G43192,G43193,G43194,G43195,G43196,G43197,G43198,G43199,G43200,
       G43201,G43202,G43203,G43204,G43205,G43206,G43207,G43208,G43209,G43210,G43211,G43212,G43213,G43214,G43215,G43216,G43217,G43218,G43219,G43220,
       G43221,G43222,G43223,G43224,G43225,G43226,G43227,G43228,G43229,G43230,G43231,G43232,G43233,G43234,G43235,G43236,G43237,G43238,G43239,G43240,
       G43241,G43242,G43243,G43244,G43245,G43246,G43247,G43248,G43249,G43250,G43251,G43252,G43253,G43254,G43255,G43256,G43257,G43258,G43259,G43260,
       G43261,G43262,G43263,G43264,G43265,G43266,G43267,G43268,G43269,G43270,G43271,G43272,G43273,G43274,G43275,G43276,G43277,G43278,G43279,G43280,
       G43281,G43282,G43283,G43284,G43285,G43286,G43287,G43288,G43289,G43290,G43291,G43292,G43293,G43294,G43295,G43296,G43297,G43298,G43299,G43300,
       G43301,G43302,G43303,G43304,G43305,G43306,G43307,G43308,G43309,G43310,G43311,G43312,G43313,G43314,G43315,G43316,G43317,G43318,G43319,G43320,
       G43321,G43322,G43323,G43324,G43325,G43326,G43327,G43328,G43329,G43330,G43331,G43332,G43333,G43334,G43335,G43336,G43337,G43338,G43339,G43340,
       G43341,G43342,G43343,G43344,G43345,G43346,G43347,G43348,G43349,G43350,G43351,G43352,G43353,G43354,G43355,G43356,G43357,G43358,G43359,G43360,
       G43361,G43362,G43363,G43364,G43365,G43366,G43367,G43368,G43369,G43370,G43371,G43372,G43373,G43374,G43375,G43376,G43377,G43378,G43379,G43380,
       G43381,G43382,G43383,G43384,G43385,G43386,G43387,G43388,G43389,G43390,G43391,G43392,G43393,G43394,G43395,G43396,G43397,G43398,G43399,G43400,
       G43401,G43402,G43403,G43404,G43405,G43406,G43407,G43408,G43409,G43410,G43411,G43412,G43413,G43414,G43415,G43416,G43417,G43418,G43419,G43420,
       G43421,G43422,G43423,G43424,G43425,G43426,G43427,G43428,G43429,G43430,G43431,G43432,G43433,G43434,G43435,G43436,G43437,G43438,G43439,G43440,
       G43441,G43442,G43443,G43444,G43445,G43446,G43447,G43448,G43449,G43450,G43451,G43452,G43453,G43454,G43455,G43456,G43457,G43458,G43459,G43460,
       G43461,G43462,G43463,G43464,G43465,G43466,G43467,G43468,G43469,G43470,G43471,G43472,G43473,G43474,G43475,G43476,G43477,G43478,G43479,G43480,
       G43481,G43482,G43483,G43484,G43485,G43486,G43487,G43488,G43489,G43490,G43491,G43492,G43493,G43494,G43495,G43496,G43497,G43498,G43499,G43500,
       G43501,G43502,G43503,G43504,G43505,G43506,G43507,G43508,G43509,G43510,G43511,G43512,G43513,G43514,G43515,G43516,G43517,G43518,G43519,G43520,
       G43521,G43522,G43523,G43524,G43525,G43526,G43527,G43528,G43529,G43530,G43531,G43532,G43533,G43534,G43535,G43536,G43537,G43538,G43539,G43540,
       G43541,G43542,G43543,G43544,G43545,G43546,G43547,G43548,G43549,G43550,G43551,G43552,G43553,G43554,G43555,G43556,G43557,G43558,G43559,G43560,
       G43561,G43562,G43563,G43564,G43565,G43566,G43567,G43568,G43569,G43570,G43571,G43572,G43573,G43574,G43575,G43576,G43577,G43578,G43579,G43580,
       G43581,G43582,G43583,G43584,G43585,G43586,G43587,G43588,G43589,G43590,G43591,G43592,G43593,G43594,G43595,G43596,G43597,G43598,G43599,G43600,
       G43601,G43602,G43603,G43604,G43605,G43606,G43607,G43608,G43609,G43610,G43611,G43612,G43613,G43614,G43615,G43616,G43617,G43618,G43619,G43620,
       G43621,G43622,G43623,G43624,G43625,G43626,G43627,G43628,G43629,G43630,G43631,G43632,G43633,G43634,G43635,G43636,G43637,G43638,G43639,G43640,
       G43641,G43642,G43643,G43644,G43645,G43646,G43647,G43648,G43649,G43650,G43651,G43652,G43653,G43654,G43655,G43656,G43657,G43658,G43659,G43660,
       G43661,G43662,G43663,G43664,G43665,G43666,G43667,G43668,G43669,G43670,G43671,G43672,G43673,G43674,G43675,G43676,G43677,G43678,G43679,G43680,
       G43681,G43682,G43683,G43684,G43685,G43686,G43687,G43688,G43689,G43690,G43691,G43692,G43693,G43694,G43695,G43696,G43697,G43698,G43699,G43700,
       G43701,G43702,G43703,G43704,G43705,G43706,G43707,G43708,G43709,G43710,G43711,G43712,G43713,G43714,G43715,G43716,G43717,G43718,G43719,G43720,
       G43721,G43722,G43723,G43724,G43725,G43726,G43727,G43728,G43729,G43730,G43731,G43732,G43733,G43734,G43735,G43736,G43737,G43738,G43739,G43740,
       G43741,G43742,G43743,G43744,G43745,G43746,G43747,G43748,G43749,G43750,G43751,G43752,G43753,G43754,G43755,G43756,G43757,G43758,G43759,G43760,
       G43761,G43762,G43763,G43764,G43765,G43766,G43767,G43768,G43769,G43770,G43771,G43772,G43773,G43774,G43775,G43776,G43777,G43778,G43779,G43780,
       G43781,G43782,G43783,G43784,G43785,G43786,G43787,G43788,G43789,G43790,G43791,G43792,G43793,G43794,G43795,G43796,G43797,G43798,G43799,G43800,
       G43801,G43802,G43803,G43804,G43805,G43806,G43807,G43808,G43809,G43810,G43811,G43812,G43813,G43814,G43815,G43816,G43817,G43818,G43819,G43820,
       G43821,G43822,G43823,G43824,G43825,G43826,G43827,G43828,G43829,G43830,G43831,G43832,G43833,G43834,G43835,G43836,G43837,G43838,G43839,G43840,
       G43841,G43842,G43843,G43844,G43845,G43846,G43847,G43848,G43849,G43850,G43851,G43852,G43853,G43854,G43855,G43856,G43857,G43858,G43859,G43860,
       G43861,G43862,G43863,G43864,G43865,G43866,G43867,G43868,G43869,G43870,G43871,G43872,G43873,G43874,G43875,G43876,G43877,G43878,G43879,G43880,
       G43881,G43882,G43883,G43884,G43885,G43886,G43887,G43888,G43889,G43890,G43891,G43892,G43893,G43894,G43895,G43896,G43897,G43898,G43899,G43900,
       G43901,G43902,G43903,G43904,G43905,G43906,G43907,G43908,G43909,G43910,G43911,G43912,G43913,G43914,G43915,G43916,G43917,G43918,G43919,G43920,
       G43921,G43922,G43923,G43924,G43925,G43926,G43927,G43928,G43929,G43930,G43931,G43932,G43933,G43934,G43935,G43936,G43937,G43938,G43939,G43940,
       G43941,G43942,G43943,G43944,G43945,G43946,G43947,G43948,G43949,G43950,G43951,G43952,G43953,G43954,G43955,G43956,G43957,G43958,G43959,G43960,
       G43961,G43962,G43963,G43964,G43965,G43966,G43967,G43968,G43969,G43970,G43971,G43972,G43973,G43974,G43975,G43976,G43977,G43978,G43979,G43980,
       G43981,G43982,G43983,G43984,G43985,G43986,G43987,G43988,G43989,G43990,G43991,G43992,G43993,G43994,G43995,G43996,G43997,G43998,G43999,G44000,
       G44001,G44002,G44003,G44004,G44005,G44006,G44007,G44008,G44009,G44010,G44011,G44012,G44013,G44014,G44015,G44016,G44017,G44018,G44019,G44020,
       G44021,G44022,G44023,G44024,G44025,G44026,G44027,G44028,G44029,G44030,G44031,G44032,G44033,G44034,G44035,G44036,G44037,G44038,G44039,G44040,
       G44041,G44042,G44043,G44044,G44045,G44046,G44047,G44048,G44049,G44050,G44051,G44052,G44053,G44054,G44055,G44056,G44057,G44058,G44059,G44060,
       G44061,G44062,G44063,G44064,G44065,G44066,G44067,G44068,G44069,G44070,G44071,G44072,G44073,G44074,G44075,G44076,G44077,G44078,G44079,G44080,
       G44081,G44082,G44083,G44084,G44085,G44086,G44087,G44088,G44089,G44090,G44091,G44092,G44093,G44094,G44095,G44096,G44097,G44098,G44099,G44100,
       G44101,G44102,G44103,G44104,G44105,G44106,G44107,G44108,G44109,G44110,G44111,G44112,G44113,G44114,G44115,G44116,G44117,G44118,G44119,G44120,
       G44121,G44122,G44123,G44124,G44125,G44126,G44127,G44128,G44129,G44130,G44131,G44132,G44133,G44134,G44135,G44136,G44137,G44138,G44139,G44140,
       G44141,G44142,G44143,G44144,G44145,G44146,G44147,G44148,G44149,G44150,G44151,G44152,G44153,G44154,G44155,G44156,G44157,G44158,G44159,G44160,
       G44161,G44162,G44163,G44164,G44165,G44166,G44167,G44168,G44169,G44170,G44171,G44172,G44173,G44174,G44175,G44176,G44177,G44178,G44179,G44180,
       G44181,G44182,G44183,G44184,G44185,G44186,G44187,G44188,G44189,G44190,G44191,G44192,G44193,G44194,G44195,G44196,G44197,G44198,G44199,G44200,
       G44201,G44202,G44203,G44204,G44205,G44206,G44207,G44208,G44209,G44210,G44211,G44212,G44213,G44214,G44215,G44216,G44217,G44218,G44219,G44220,
       G44221,G44222,G44223,G44224,G44225,G44226,G44227,G44228,G44229,G44230,G44231,G44232,G44233,G44234,G44235,G44236,G44237,G44238,G44239,G44240,
       G44241,G44242,G44243,G44244,G44245,G44246,G44247,G44248,G44249,G44250,G44251,G44252,G44253,G44254,G44255,G44256,G44257,G44258,G44259,G44260,
       G44261,G44262,G44263,G44264,G44265,G44266,G44267,G44268,G44269,G44270,G44271,G44272,G44273,G44274,G44275,G44276,G44277,G44278,G44279,G44280,
       G44281,G44282,G44283,G44284,G44285,G44286,G44287,G44288,G44289,G44290,G44291,G44292,G44293,G44294,G44295,G44296,G44297,G44298,G44299,G44300,
       G44301,G44302,G44303,G44304,G44305,G44306,G44307,G44308,G44309,G44310,G44311,G44312,G44313,G44314,G44315,G44316,G44317,G44318,G44319,G44320,
       G44321,G44322,G44323,G44324,G44325,G44326,G44327,G44328,G44329,G44330,G44331,G44332,G44333,G44334,G44335,G44336,G44337,G44338,G44339,G44340,
       G44341,G44342,G44343,G44344,G44345,G44346,G44347,G44348,G44349,G44350,G44351,G44352,G44353,G44354,G44355,G44356,G44357,G44358,G44359,G44360,
       G44361,G44362,G44363,G44364,G44365,G44366,G44367,G44368,G44369,G44370,G44371,G44372,G44373,G44374,G44375,G44376,G44377,G44378,G44379,G44380,
       G44381,G44382,G44383,G44384,G44385,G44386,G44387,G44388,G44389,G44390,G44391,G44392,G44393,G44394,G44395,G44396,G44397,G44398,G44399,G44400,
       G44401,G44402,G44403,G44404,G44405,G44406,G44407,G44408,G44409,G44410,G44411,G44412,G44413,G44414,G44415,G44416,G44417,G44418,G44419,G44420,
       G44421,G44422,G44423,G44424,G44425,G44426,G44427,G44428,G44429,G44430,G44431,G44432,G44433,G44434,G44435,G44436,G44437,G44438,G44439,G44440,
       G44441,G44442,G44443,G44444,G44445,G44446,G44447,G44448,G44449,G44450,G44451,G44452,G44453,G44454,G44455,G44456,G44457,G44458,G44459,G44460,
       G44461,G44462,G44463,G44464,G44465,G44466,G44467,G44468,G44469,G44470,G44471,G44472,G44473,G44474,G44475,G44476,G44477,G44478,G44479,G44480,
       G44481,G44482,G44483,G44484,G44485,G44486,G44487,G44488,G44489,G44490,G44491,G44492,G44493,G44494,G44495,G44496,G44497,G44498,G44499,G44500,
       G44501,G44502,G44503,G44504,G44505,G44506,G44507,G44508,G44509,G44510,G44511,G44512,G44513,G44514,G44515,G44516,G44517,G44518,G44519,G44520,
       G44521,G44522,G44523,G44524,G44525,G44526,G44527,G44528,G44529,G44530,G44531,G44532,G44533,G44534,G44535,G44536,G44537,G44538,G44539,G44540,
       G44541,G44542,G44543,G44544,G44545,G44546,G44547,G44548,G44549,G44550,G44551,G44552,G44553,G44554,G44555,G44556,G44557,G44558,G44559,G44560,
       G44561,G44562,G44563,G44564,G44565,G44566,G44567,G44568,G44569,G44570,G44571,G44572,G44573,G44574,G44575,G44576,G44577,G44578,G44579,G44580,
       G44581,G44582,G44583,G44584,G44585,G44586,G44587,G44588,G44589,G44590,G44591,G44592,G44593,G44594,G44595,G44596,G44597,G44598,G44599,G44600,
       G44601,G44602,G44603,G44604,G44605,G44606,G44607,G44608,G44609,G44610,G44611,G44612,G44613,G44614,G44615,G44616,G44617,G44618,G44619,G44620,
       G44621,G44622,G44623,G44624,G44625,G44626,G44627,G44628,G44629,G44630,G44631,G44632,G44633,G44634,G44635,G44636,G44637,G44638,G44639,G44640,
       G44641,G44642,G44643,G44644,G44645,G44646,G44647,G44648,G44649,G44650,G44651,G44652,G44653,G44654,G44655,G44656,G44657,G44658,G44659,G44660,
       G44661,G44662,G44663,G44664,G44665,G44666,G44667,G44668,G44669,G44670,G44671,G44672,G44673,G44674,G44675,G44676,G44677,G44678,G44679,G44680,
       G44681,G44682,G44683,G44684,G44685,G44686,G44687,G44688,G44689,G44690,G44691,G44692,G44693,G44694,G44695,G44696,G44697,G44698,G44699,G44700,
       G44701,G44702,G44703,G44704,G44705,G44706,G44707,G44708,G44709,G44710,G44711,G44712,G44713,G44714,G44715,G44716,G44717,G44718,G44719,G44720,
       G44721,G44722,G44723,G44724,G44725,G44726,G44727,G44728,G44729,G44730,G44731,G44732,G44733,G44734,G44735,G44736,G44737,G44738,G44739,G44740,
       G44741,G44742,G44743,G44744,G44745,G44746,G44747,G44748,G44749,G44750,G44751,G44752,G44753,G44754,G44755,G44756,G44757,G44758,G44759,G44760,
       G44761,G44762,G44763,G44764,G44765,G44766,G44767,G44768,G44769,G44770,G44771,G44772,G44773,G44774,G44775,G44776,G44777,G44778,G44779,G44780,
       G44781,G44782,G44783,G44784,G44785,G44786,G44787,G44788,G44789,G44790,G44791,G44792,G44793,G44794,G44795,G44796,G44797,G44798,G44799,G44800,
       G44801,G44802,G44803,G44804,G44805,G44806,G44807,G44808,G44809,G44810,G44811,G44812,G44813,G44814,G44815,G44816,G44817,G44818,G44819,G44820,
       G44821,G44822,G44823,G44824,G44825,G44826,G44827,G44828,G44829,G44830,G44831,G44832,G44833,G44834,G44835,G44836,G44837,G44838,G44839,G44840,
       G44841,G44842,G44843,G44844,G44845,G44846,G44847,G44848,G44849,G44850,G44851,G44852,G44853,G44854,G44855,G44856,G44857,G44858,G44859,G44860,
       G44861,G44862,G44863,G44864,G44865,G44866,G44867,G44868,G44869,G44870,G44871,G44872,G44873,G44874,G44875,G44876,G44877,G44878,G44879,G44880,
       G44881,G44882,G44883,G44884,G44885,G44886,G44887,G44888,G44889,G44890,G44891,G44892,G44893,G44894,G44895,G44896,G44897,G44898,G44899,G44900,
       G44901,G44902,G44903,G44904,G44905,G44906,G44907,G44908,G44909,G44910,G44911,G44912,G44913,G44914,G44915,G44916,G44917,G44918,G44919,G44920,
       G44921,G44922,G44923,G44924,G44925,G44926,G44927,G44928,G44929,G44930,G44931,G44932,G44933,G44934,G44935,G44936,G44937,G44938,G44939,G44940,
       G44941,G44942,G44943,G44944,G44945,G44946,G44947,G44948,G44949,G44950,G44951,G44952,G44953,G44954,G44955,G44956,G44957,G44958,G44959,G44960,
       G44961,G44962,G44963,G44964,G44965,G44966,G44967,G44968,G44969,G44970,G44971,G44972,G44973,G44974,G44975,G44976,G44977,G44978,G44979,G44980,
       G44981,G44982,G44983,G44984,G44985,G44986,G44987,G44988,G44989,G44990,G44991,G44992,G44993,G44994,G44995,G44996,G44997,G44998,G44999,G45000,
       G45001,G45002,G45003,G45004,G45005,G45006,G45007,G45008,G45009,G45010,G45011,G45012,G45013,G45014,G45015,G45016,G45017,G45018,G45019,G45020,
       G45021,G45022,G45023,G45024,G45025,G45026,G45027,G45028,G45029,G45030,G45031,G45032,G45033,G45034,G45035,G45036,G45037,G45038,G45039,G45040,
       G45041,G45042,G45043,G45044,G45045,G45046,G45047,G45048,G45049,G45050,G45051,G45052,G45053,G45054,G45055,G45056,G45057,G45058,G45059,G45060,
       G45061,G45062,G45063,G45064,G45065,G45066,G45067,G45068,G45069,G45070,G45071,G45072,G45073,G45074,G45075,G45076,G45077,G45078,G45079,G45080,
       G45081,G45082,G45083,G45084,G45085,G45086,G45087,G45088,G45089,G45090,G45091,G45092,G45093,G45094,G45095,G45096,G45097,G45098,G45099,G45100,
       G45101,G45102,G45103,G45104,G45105,G45106,G45107,G45108,G45109,G45110,G45111,G45112,G45113,G45114,G45115,G45116,G45117,G45118,G45119,G45120,
       G45121,G45122,G45123,G45124,G45125,G45126,G45127,G45128,G45129,G45130,G45131,G45132,G45133,G45134,G45135,G45136,G45137,G45138,G45139,G45140,
       G45141,G45142,G45143,G45144,G45145,G45146,G45147,G45148,G45149,G45150,G45151,G45152,G45153,G45154,G45155,G45156,G45157,G45158,G45159,G45160,
       G45161,G45162,G45163,G45164,G45165,G45166,G45167,G45168,G45169,G45170,G45171,G45172,G45173,G45174,G45175,G45176,G45177,G45178,G45179,G45180,
       G45181,G45182,G45183,G45184,G45185,G45186,G45187,G45188,G45189,G45190,G45191,G45192,G45193,G45194,G45195,G45196,G45197,G45198,G45199,G45200,
       G45201,G45202,G45203,G45204,G45205,G45206,G45207,G45208,G45209,G45210,G45211,G45212,G45213,G45214,G45215,G45216,G45217,G45218,G45219,G45220,
       G45221,G45222,G45223,G45224,G45225,G45226,G45227,G45228,G45229,G45230,G45231,G45232,G45233,G45234,G45235,G45236,G45237,G45238,G45239,G45240,
       G45241,G45242,G45243,G45244,G45245,G45246,G45247,G45248,G45249,G45250,G45251,G45252,G45253,G45254,G45255,G45256,G45257,G45258,G45259,G45260,
       G45261,G45262,G45263,G45264,G45265,G45266,G45267,G45268,G45269,G45270,G45271,G45272,G45273,G45274,G45275,G45276,G45277,G45278,G45279,G45280,
       G45281,G45282,G45283,G45284,G45285,G45286,G45287,G45288,G45289,G45290,G45291,G45292,G45293,G45294,G45295,G45296,G45297,G45298,G45299,G45300,
       G45301,G45302,G45303,G45304,G45305,G45306,G45307,G45308,G45309,G45310,G45311,G45312,G45313,G45314,G45315,G45316,G45317,G45318,G45319,G45320,
       G45321,G45322,G45323,G45324,G45325,G45326,G45327,G45328,G45329,G45330,G45331,G45332,G45333,G45334,G45335,G45336,G45337,G45338,G45339,G45340,
       G45341,G45342,G45343,G45344,G45345,G45346,G45347,G45348,G45349,G45350,G45351,G45352,G45353,G45354,G45355,G45356,G45357,G45358,G45359,G45360,
       G45361,G45362,G45363,G45364,G45365,G45366,G45367,G45368,G45369,G45370,G45371,G45372,G45373,G45374,G45375,G45376,G45377,G45378,G45379,G45380,
       G45381,G45382,G45383,G45384,G45385,G45386,G45387,G45388,G45389,G45390,G45391,G45392,G45393,G45394,G45395,G45396,G45397,G45398,G45399,G45400,
       G45401,G45402,G45403,G45404,G45405,G45406,G45407,G45408,G45409,G45410,G45411,G45412,G45413,G45414,G45415,G45416,G45417,G45418,G45419,G45420,
       G45421,G45422,G45423,G45424,G45425,G45426,G45427,G45428,G45429,G45430,G45431,G45432,G45433,G45434,G45435,G45436,G45437,G45438,G45439,G45440,
       G45441,G45442,G45443,G45444,G45445,G45446,G45447,G45448,G45449,G45450,G45451,G45452,G45453,G45454,G45455,G45456,G45457,G45458,G45459,G45460,
       G45461,G45462,G45463,G45464,G45465,G45466,G45467,G45468,G45469,G45470,G45471,G45472,G45473,G45474,G45475,G45476,G45477,G45478,G45479,G45480,
       G45481,G45482,G45483,G45484,G45485,G45486,G45487,G45488,G45489,G45490,G45491,G45492,G45493,G45494,G45495,G45496,G45497,G45498,G45499,G45500,
       G45501,G45502,G45503,G45504,G45505,G45506,G45507,G45508,G45509,G45510,G45511,G45512,G45513,G45514,G45515,G45516,G45517,G45518,G45519,G45520,
       G45521,G45522,G45523,G45524,G45525,G45526,G45527,G45528,G45529,G45530,G45531,G45532,G45533,G45534,G45535,G45536,G45537,G45538,G45539,G45540,
       G45541,G45542,G45543,G45544,G45545,G45546,G45547,G45548,G45549,G45550,G45551,G45552,G45553,G45554,G45555,G45556,G45557,G45558,G45559,G45560,
       G45561,G45562,G45563,G45564,G45565,G45566,G45567,G45568,G45569,G45570,G45571,G45572,G45573,G45574,G45575,G45576,G45577,G45578,G45579,G45580,
       G45581,G45582,G45583,G45584,G45585,G45586,G45587,G45588,G45589,G45590,G45591,G45592,G45593,G45594,G45595,G45596,G45597,G45598,G45599,G45600,
       G45601,G45602,G45603,G45604,G45605,G45606,G45607,G45608,G45609,G45610,G45611,G45612,G45613,G45614,G45615,G45616,G45617,G45618,G45619,G45620,
       G45621,G45622,G45623,G45624,G45625,G45626,G45627,G45628,G45629,G45630,G45631,G45632,G45633,G45634,G45635,G45636,G45637,G45638,G45639,G45640,
       G45641,G45642,G45643,G45644,G45645,G45646,G45647,G45648,G45649,G45650,G45651,G45652,G45653,G45654,G45655,G45656,G45657,G45658,G45659,G45660,
       G45661,G45662,G45663,G45664,G45665,G45666,G45667,G45668,G45669,G45670,G45671,G45672,G45673,G45674,G45675,G45676,G45677,G45678,G45679,G45680,
       G45681,G45682,G45683,G45684,G45685,G45686,G45687,G45688,G45689,G45690,G45691,G45692,G45693,G45694,G45695,G45696,G45697,G45698,G45699,G45700,
       G45701,G45702,G45703,G45704,G45705,G45706,G45707,G45708,G45709,G45710,G45711,G45712,G45713,G45714,G45715,G45716,G45717,G45718,G45719,G45720,
       G45721,G45722,G45723,G45724,G45725,G45726,G45727,G45728,G45729,G45730,G45731,G45732,G45733,G45734,G45735,G45736,G45737,G45738,G45739,G45740,
       G45741,G45742,G45743,G45744,G45745,G45746,G45747,G45748,G45749,G45750,G45751,G45752,G45753,G45754,G45755,G45756,G45757,G45758,G45759,G45760,
       G45761,G45762,G45763,G45764,G45765,G45766,G45767,G45768,G45769,G45770,G45771,G45772,G45773,G45774,G45775,G45776,G45777,G45778,G45779,G45780,
       G45781,G45782,G45783,G45784,G45785,G45786,G45787,G45788,G45789,G45790,G45791,G45792,G45793,G45794,G45795,G45796,G45797,G45798,G45799,G45800,
       G45801,G45802,G45803,G45804,G45805,G45806,G45807,G45808,G45809,G45810,G45811,G45812,G45813,G45814,G45815,G45816,G45817,G45818,G45819,G45820,
       G45821,G45822,G45823,G45824,G45825,G45826,G45827,G45828,G45829,G45830,G45831,G45832,G45833,G45834,G45835,G45836,G45837,G45838,G45839,G45840,
       G45841,G45842,G45843,G45844,G45845,G45846,G45847,G45848,G45849,G45850,G45851,G45852,G45853,G45854,G45855,G45856,G45857,G45858,G45859,G45860,
       G45861,G45862,G45863,G45864,G45865,G45866,G45867,G45868,G45869,G45870,G45871,G45872,G45873,G45874,G45875,G45876,G45877,G45878,G45879,G45880,
       G45881,G45882,G45883,G45884,G45885,G45886,G45887,G45888,G45889,G45890,G45891,G45892,G45893,G45894,G45895,G45896,G45897,G45898,G45899,G45900,
       G45901,G45902,G45903,G45904,G45905,G45906,G45907,G45908,G45909,G45910,G45911,G45912,G45913,G45914,G45915,G45916,G45917,G45918,G45919,G45920,
       G45921,G45922,G45923,G45924,G45925,G45926,G45927,G45928,G45929,G45930,G45931,G45932,G45933,G45934,G45935,G45936,G45937,G45938,G45939,G45940,
       G45941,G45942,G45943,G45944,G45945,G45946,G45947,G45948,G45949,G45950,G45951,G45952,G45953,G45954,G45955,G45956,G45957,G45958,G45959,G45960,
       G45961,G45962,G45963,G45964,G45965,G45966,G45967,G45968,G45969,G45970,G45971,G45972,G45973,G45974,G45975,G45976,G45977,G45978,G45979,G45980,
       G45981,G45982,G45983,G45984,G45985,G45986,G45987,G45988,G45989,G45990,G45991,G45992,G45993,G45994,G45995,G45996,G45997,G45998,G45999,G46000,
       G46001,G46002,G46003,G46004,G46005,G46006,G46007,G46008,G46009,G46010,G46011,G46012,G46013,G46014,G46015,G46016,G46017,G46018,G46019,G46020,
       G46021,G46022,G46023,G46024,G46025,G46026,G46027,G46028,G46029,G46030,G46031,G46032,G46033,G46034,G46035,G46036,G46037,G46038,G46039,G46040,
       G46041,G46042,G46043,G46044,G46045,G46046,G46047,G46048,G46049,G46050,G46051,G46052,G46053,G46054,G46055,G46056,G46057,G46058,G46059,G46060,
       G46061,G46062,G46063,G46064,G46065,G46066,G46067,G46068,G46069,G46070,G46071,G46072,G46073,G46074,G46075,G46076,G46077,G46078,G46079,G46080,
       G46081,G46082,G46083,G46084,G46085,G46086,G46087,G46088,G46089,G46090,G46091,G46092,G46093,G46094,G46095,G46096,G46097,G46098,G46099,G46100,
       G46101,G46102,G46103,G46104,G46105,G46106,G46107,G46108,G46109,G46110,G46111,G46112,G46113,G46114,G46115,G46116,G46117,G46118,G46119,G46120,
       G46121,G46122,G46123,G46124,G46125,G46126,G46127,G46128,G46129,G46130,G46131,G46132,G46133,G46134,G46135,G46136,G46137,G46138,G46139,G46140,
       G46141,G46142,G46143,G46144,G46145,G46146,G46147,G46148,G46149,G46150,G46151,G46152,G46153,G46154,G46155,G46156,G46157,G46158,G46159,G46160,
       G46161,G46162,G46163,G46164,G46165,G46166,G46167,G46168,G46169,G46170,G46171,G46172,G46173,G46174,G46175,G46176,G46177,G46178,G46179,G46180,
       G46181,G46182,G46183,G46184,G46185,G46186,G46187,G46188,G46189,G46190,G46191,G46192,G46193,G46194,G46195,G46196,G46197,G46198,G46199,G46200,
       G46201,G46202,G46203,G46204,G46205,G46206,G46207,G46208,G46209,G46210,G46211,G46212,G46213,G46214,G46215,G46216,G46217,G46218,G46219,G46220,
       G46221,G46222,G46223,G46224,G46225,G46226,G46227,G46228,G46229,G46230,G46231,G46232,G46233,G46234,G46235,G46236,G46237,G46238,G46239,G46240,
       G46241,G46242,G46243,G46244,G46245,G46246,G46247,G46248,G46249,G46250,G46251,G46252,G46253,G46254,G46255,G46256,G46257,G46258,G46259,G46260,
       G46261,G46262,G46263,G46264,G46265,G46266,G46267,G46268,G46269,G46270,G46271,G46272,G46273,G46274,G46275,G46276,G46277,G46278,G46279,G46280,
       G46281,G46282,G46283,G46284,G46285,G46286,G46287,G46288,G46289,G46290,G46291,G46292,G46293,G46294,G46295,G46296,G46297,G46298,G46299,G46300,
       G46301,G46302,G46303,G46304,G46305,G46306,G46307,G46308,G46309,G46310,G46311,G46312,G46313,G46314,G46315,G46316,G46317,G46318,G46319,G46320,
       G46321,G46322,G46323,G46324,G46325,G46326,G46327,G46328,G46329,G46330,G46331,G46332,G46333,G46334,G46335,G46336,G46337,G46338,G46339,G46340,
       G46341,G46342,G46343,G46344,G46345,G46346,G46347,G46348,G46349,G46350,G46351,G46352,G46353,G46354,G46355,G46356,G46357,G46358,G46359,G46360,
       G46361,G46362,G46363,G46364,G46365,G46366,G46367,G46368,G46369,G46370,G46371,G46372,G46373,G46374,G46375,G46376,G46377,G46378,G46379,G46380,
       G46381,G46382,G46383,G46384,G46385,G46386,G46387,G46388,G46389,G46390,G46391,G46392,G46393,G46394,G46395,G46396,G46397,G46398,G46399,G46400,
       G46401,G46402,G46403,G46404,G46405,G46406,G46407,G46408,G46409,G46410,G46411,G46412,G46413,G46414,G46415,G46416,G46417,G46418,G46419,G46420,
       G46421,G46422,G46423,G46424,G46425,G46426,G46427,G46428,G46429,G46430,G46431,G46432,G46433,G46434,G46435,G46436,G46437,G46438,G46439,G46440,
       G46441,G46442,G46443,G46444,G46445,G46446,G46447,G46448,G46449,G46450,G46451,G46452,G46453,G46454,G46455,G46456,G46457,G46458,G46459,G46460,
       G46461,G46462,G46463,G46464,G46465,G46466,G46467,G46468,G46469,G46470,G46471,G46472,G46473,G46474,G46475,G46476,G46477,G46478,G46479,G46480,
       G46481,G46482,G46483,G46484,G46485,G46486,G46487,G46488,G46489,G46490,G46491,G46492,G46493,G46494,G46495,G46496,G46497,G46498,G46499,G46500,
       G46501,G46502,G46503,G46504,G46505,G46506,G46507,G46508,G46509,G46510,G46511,G46512,G46513,G46514,G46515,G46516,G46517,G46518,G46519,G46520,
       G46521,G46522,G46523,G46524,G46525,G46526,G46527,G46528,G46529,G46530,G46531,G46532,G46533,G46534,G46535,G46536,G46537,G46538,G46539,G46540,
       G46541,G46542,G46543,G46544,G46545,G46546,G46547,G46548,G46549,G46550,G46551,G46552,G46553,G46554,G46555,G46556,G46557,G46558,G46559,G46560,
       G46561,G46562,G46563,G46564,G46565,G46566,G46567,G46568,G46569,G46570,G46571,G46572,G46573,G46574,G46575,G46576,G46577,G46578,G46579,G46580,
       G46581,G46582,G46583,G46584,G46585,G46586,G46587,G46588,G46589,G46590,G46591,G46592,G46593,G46594,G46595,G46596,G46597,G46598,G46599,G46600,
       G46601,G46602,G46603,G46604,G46605,G46606,G46607,G46608,G46609,G46610,G46611,G46612,G46613,G46614,G46615,G46616,G46617,G46618,G46619,G46620,
       G46621,G46622,G46623,G46624,G46625,G46626,G46627,G46628,G46629,G46630,G46631,G46632,G46633,G46634,G46635,G46636,G46637,G46638,G46639,G46640,
       G46641,G46642,G46643,G46644,G46645,G46646,G46647,G46648,G46649,G46650,G46651,G46652,G46653,G46654,G46655,G46656,G46657,G46658,G46659,G46660,
       G46661,G46662,G46663,G46664,G46665,G46666,G46667,G46668,G46669,G46670,G46671,G46672,G46673,G46674,G46675,G46676,G46677,G46678,G46679,G46680,
       G46681,G46682,G46683,G46684,G46685,G46686,G46687,G46688,G46689,G46690,G46691,G46692,G46693,G46694,G46695,G46696,G46697,G46698,G46699,G46700,
       G46701,G46702,G46703,G46704,G46705,G46706,G46707,G46708,G46709,G46710,G46711,G46712,G46713,G46714,G46715,G46716,G46717,G46718,G46719,G46720,
       G46721,G46722,G46723,G46724,G46725,G46726,G46727,G46728,G46729,G46730,G46731,G46732,G46733,G46734,G46735,G46736,G46737,G46738,G46739,G46740,
       G46741,G46742,G46743,G46744,G46745,G46746,G46747,G46748,G46749,G46750,G46751,G46752,G46753,G46754,G46755,G46756,G46757,G46758,G46759,G46760,
       G46761,G46762,G46763,G46764,G46765,G46766,G46767,G46768,G46769,G46770,G46771,G46772,G46773,G46774,G46775,G46776,G46777,G46778,G46779,G46780,
       G46781,G46782,G46783,G46784,G46785,G46786,G46787,G46788,G46789,G46790,G46791,G46792,G46793,G46794,G46795,G46796,G46797,G46798,G46799,G46800,
       G46801,G46802,G46803,G46804,G46805,G46806,G46807,G46808,G46809,G46810,G46811,G46812,G46813,G46814,G46815,G46816,G46817,G46818,G46819,G46820,
       G46821,G46822,G46823,G46824,G46825,G46826,G46827,G46828,G46829,G46830,G46831,G46832,G46833,G46834,G46835,G46836,G46837,G46838,G46839,G46840,
       G46841,G46842,G46843,G46844,G46845,G46846,G46847,G46848,G46849,G46850,G46851,G46852,G46853,G46854,G46855,G46856,G46857,G46858,G46859,G46860,
       G46861,G46862,G46863,G46864,G46865,G46866,G46867,G46868,G46869,G46870,G46871,G46872,G46873,G46874,G46875,G46876,G46877,G46878,G46879,G46880,
       G46881,G46882,G46883,G46884,G46885,G46886,G46887,G46888,G46889,G46890,G46891,G46892,G46893,G46894,G46895,G46896,G46897,G46898,G46899,G46900,
       G46901,G46902,G46903,G46904,G46905,G46906,G46907,G46908,G46909,G46910,G46911,G46912,G46913,G46914,G46915,G46916,G46917,G46918,G46919,G46920,
       G46921,G46922,G46923,G46924,G46925,G46926,G46927,G46928,G46929,G46930,G46931,G46932,G46933,G46934,G46935,G46936,G46937,G46938,G46939,G46940,
       G46941,G46942,G46943,G46944,G46945,G46946,G46947,G46948,G46949,G46950,G46951,G46952,G46953,G46954,G46955,G46956,G46957,G46958,G46959,G46960,
       G46961,G46962,G46963,G46964,G46965,G46966,G46967,G46968,G46969,G46970,G46971,G46972,G46973,G46974,G46975,G46976,G46977,G46978,G46979,G46980,
       G46981,G46982,G46983,G46984,G46985,G46986,G46987,G46988,G46989,G46990,G46991,G46992,G46993,G46994,G46995,G46996,G46997,G46998,G46999,G47000,
       G47001,G47002,G47003,G47004,G47005,G47006,G47007,G47008,G47009,G47010,G47011,G47012,G47013,G47014,G47015,G47016,G47017,G47018,G47019,G47020,
       G47021,G47022,G47023,G47024,G47025,G47026,G47027,G47028,G47029,G47030,G47031,G47032,G47033,G47034,G47035,G47036,G47037,G47038,G47039,G47040,
       G47041,G47042,G47043,G47044,G47045,G47046,G47047,G47048,G47049,G47050,G47051,G47052,G47053,G47054,G47055,G47056,G47057,G47058,G47059,G47060,
       G47061,G47062,G47063,G47064,G47065,G47066,G47067,G47068,G47069,G47070,G47071,G47072,G47073,G47074,G47075,G47076,G47077,G47078,G47079,G47080,
       G47081,G47082,G47083,G47084,G47085,G47086,G47087,G47088,G47089,G47090,G47091,G47092,G47093,G47094,G47095,G47096,G47097,G47098,G47099,G47100,
       G47101,G47102,G47103,G47104,G47105,G47106,G47107,G47108,G47109,G47110,G47111,G47112,G47113,G47114,G47115,G47116,G47117,G47118,G47119,G47120,
       G47121,G47122,G47123,G47124,G47125,G47126,G47127,G47128,G47129,G47130,G47131,G47132,G47133,G47134,G47135,G47136,G47137,G47138,G47139,G47140,
       G47141,G47142,G47143,G47144,G47145,G47146,G47147,G47148,G47149,G47150,G47151,G47152,G47153,G47154,G47155,G47156,G47157,G47158,G47159,G47160,
       G47161,G47162,G47163,G47164,G47165,G47166,G47167,G47168,G47169,G47170,G47171,G47172,G47173,G47174,G47175,G47176,G47177,G47178,G47179,G47180,
       G47181,G47182,G47183,G47184,G47185,G47186,G47187,G47188,G47189,G47190,G47191,G47192,G47193,G47194,G47195,G47196,G47197,G47198,G47199,G47200,
       G47201,G47202,G47203,G47204,G47205,G47206,G47207,G47208,G47209,G47210,G47211,G47212,G47213,G47214,G47215,G47216,G47217,G47218,G47219,G47220,
       G47221,G47222,G47223,G47224,G47225,G47226,G47227,G47228,G47229,G47230,G47231,G47232,G47233,G47234,G47235,G47236,G47237,G47238,G47239,G47240,
       G47241,G47242,G47243,G47244,G47245,G47246,G47247,G47248,G47249,G47250,G47251,G47252,G47253,G47254,G47255,G47256,G47257,G47258,G47259,G47260,
       G47261,G47262,G47263,G47264,G47265,G47266,G47267,G47268,G47269,G47270,G47271,G47272,G47273,G47274,G47275,G47276,G47277,G47278,G47279,G47280,
       G47281,G47282,G47283,G47284,G47285,G47286,G47287,G47288,G47289,G47290,G47291,G47292,G47293,G47294,G47295,G47296,G47297,G47298,G47299,G47300,
       G47301,G47302,G47303,G47304,G47305,G47306,G47307,G47308,G47309,G47310,G47311,G47312,G47313,G47314,G47315,G47316,G47317,G47318,G47319,G47320,
       G47321,G47322,G47323,G47324,G47325,G47326,G47327,G47328,G47329,G47330,G47331,G47332,G47333,G47334,G47335,G47336,G47337,G47338,G47339,G47340,
       G47341,G47342,G47343,G47344,G47345,G47346,G47347,G47348,G47349,G47350,G47351,G47352,G47353,G47354,G47355,G47356,G47357,G47358,G47359,G47360,
       G47361,G47362,G47363,G47364,G47365,G47366,G47367,G47368,G47369,G47370,G47371,G47372,G47373,G47374,G47375,G47376,G47377,G47378,G47379,G47380,
       G47381,G47382,G47383,G47384,G47385,G47386,G47387,G47388,G47389,G47390,G47391,G47392,G47393,G47394,G47395,G47396,G47397,G47398,G47399,G47400,
       G47401,G47402,G47403,G47404,G47405,G47406,G47407,G47408,G47409,G47410,G47411,G47412,G47413,G47414,G47415,G47416,G47417,G47418,G47419,G47420,
       G47421,G47422,G47423,G47424,G47425,G47426,G47427,G47428,G47429,G47430,G47431,G47432,G47433,G47434,G47435,G47436,G47437,G47438,G47439,G47440,
       G47441,G47442,G47443,G47444,G47445,G47446,G47447,G47448,G47449,G47450,G47451,G47452,G47453,G47454,G47455,G47456,G47457,G47458,G47459,G47460,
       G47461,G47462,G47463,G47464,G47465,G47466,G47467,G47468,G47469,G47470,G47471,G47472,G47473,G47474,G47475,G47476,G47477,G47478,G47479,G47480,
       G47481,G47482,G47483,G47484,G47485,G47486,G47487,G47488,G47489,G47490,G47491,G47492,G47493,G47494,G47495,G47496,G47497,G47498,G47499,G47500,
       G47501,G47502,G47503,G47504,G47505,G47506,G47507,G47508,G47509,G47510,G47511,G47512,G47513,G47514,G47515,G47516,G47517,G47518,G47519,G47520,
       G47521,G47522,G47523,G47524,G47525,G47526,G47527,G47528,G47529,G47530,G47531,G47532,G47533,G47534,G47535,G47536,G47537,G47538,G47539,G47540,
       G47541,G47542,G47543,G47544,G47545,G47546,G47547,G47548,G47549,G47550,G47551,G47552,G47553,G47554,G47555,G47556,G47557,G47558,G47559,G47560,
       G47561,G47562,G47563,G47564,G47565,G47566,G47567,G47568,G47569,G47570,G47571,G47572,G47573,G47574,G47575,G47576,G47577,G47578,G47579,G47580,
       G47581,G47582,G47583,G47584,G47585,G47586,G47587,G47588,G47589,G47590,G47591,G47592,G47593,G47594,G47595,G47596,G47597,G47598,G47599,G47600,
       G47601,G47602,G47603,G47604,G47605,G47606,G47607,G47608,G47609,G47610,G47611,G47612,G47613,G47614,G47615,G47616,G47617,G47618,G47619,G47620,
       G47621,G47622,G47623,G47624,G47625,G47626,G47627,G47628,G47629,G47630,G47631,G47632,G47633,G47634,G47635,G47636,G47637,G47638,G47639,G47640,
       G47641,G47642,G47643,G47644,G47645,G47646,G47647,G47648,G47649,G47650,G47651,G47652,G47653,G47654,G47655,G47656,G47657,G47658,G47659,G47660,
       G47661,G47662,G47663,G47664,G47665,G47666,G47667,G47668,G47669,G47670,G47671,G47672,G47673,G47674,G47675,G47676,G47677,G47678,G47679,G47680,
       G47681,G47682,G47683,G47684,G47685,G47686,G47687,G47688,G47689,G47690,G47691,G47692,G47693,G47694,G47695,G47696,G47697,G47698,G47699,G47700,
       G47701,G47702,G47703,G47704,G47705,G47706,G47707,G47708,G47709,G47710,G47711,G47712,G47713,G47714,G47715,G47716,G47717,G47718,G47719,G47720,
       G47721,G47722,G47723,G47724,G47725,G47726,G47727,G47728,G47729,G47730,G47731,G47732,G47733,G47734,G47735,G47736,G47737,G47738,G47739,G47740,
       G47741,G47742,G47743,G47744,G47745,G47746,G47747,G47748,G47749,G47750,G47751,G47752,G47753,G47754,G47755,G47756,G47757,G47758,G47759,G47760,
       G47761,G47762,G47763,G47764,G47765,G47766,G47767,G47768,G47769,G47770,G47771,G47772,G47773,G47774,G47775,G47776,G47777,G47778,G47779,G47780,
       G47781,G47782,G47783,G47784,G47785,G47786,G47787,G47788,G47789,G47790,G47791,G47792,G47793,G47794,G47795,G47796,G47797,G47798,G47799,G47800,
       G47801,G47802,G47803,G47804,G47805,G47806,G47807,G47808,G47809,G47810,G47811,G47812,G47813,G47814,G47815,G47816,G47817,G47818,G47819,G47820,
       G47821,G47822,G47823,G47824,G47825,G47826,G47827,G47828,G47829,G47830,G47831,G47832,G47833,G47834,G47835,G47836,G47837,G47838,G47839,G47840,
       G47841,G47842,G47843,G47844,G47845,G47846,G47847,G47848,G47849,G47850,G47851,G47852,G47853,G47854,G47855,G47856,G47857,G47858,G47859,G47860,
       G47861,G47862,G47863,G47864,G47865,G47866,G47867,G47868,G47869,G47870,G47871,G47872,G47873,G47874,G47875,G47876,G47877,G47878,G47879,G47880,
       G47881,G47882,G47883,G47884,G47885,G47886,G47887,G47888,G47889,G47890,G47891,G47892,G47893,G47894,G47895,G47896,G47897,G47898,G47899,G47900,
       G47901,G47902,G47903,G47904,G47905,G47906,G47907,G47908,G47909,G47910,G47911,G47912,G47913,G47914,G47915,G47916,G47917,G47918,G47919,G47920,
       G47921,G47922,G47923,G47924,G47925,G47926,G47927,G47928,G47929,G47930,G47931,G47932,G47933,G47934,G47935,G47936,G47937,G47938,G47939,G47940,
       G47941,G47942,G47943,G47944,G47945,G47946,G47947,G47948,G47949,G47950,G47951,G47952,G47953,G47954,G47955,G47956,G47957,G47958,G47959,G47960,
       G47961,G47962,G47963,G47964,G47965,G47966,G47967,G47968,G47969,G47970,G47971,G47972,G47973,G47974,G47975,G47976,G47977,G47978,G47979,G47980,
       G47981,G47982,G47983,G47984,G47985,G47986,G47987,G47988,G47989,G47990,G47991,G47992,G47993,G47994,G47995,G47996,G47997,G47998,G47999,G48000,
       G48001,G48002,G48003,G48004,G48005,G48006,G48007,G48008,G48009,G48010,G48011,G48012,G48013,G48014,G48015,G48016,G48017,G48018,G48019,G48020,
       G48021,G48022,G48023,G48024,G48025,G48026,G48027,G48028,G48029,G48030,G48031,G48032,G48033,G48034,G48035,G48036,G48037,G48038,G48039,G48040,
       G48041,G48042,G48043,G48044,G48045,G48046,G48047,G48048,G48049,G48050,G48051,G48052,G48053,G48054,G48055,G48056,G48057,G48058,G48059,G48060,
       G48061,G48062,G48063,G48064,G48065,G48066,G48067,G48068,G48069,G48070,G48071,G48072,G48073,G48074,G48075,G48076,G48077,G48078,G48079,G48080,
       G48081,G48082,G48083,G48084,G48085,G48086,G48087,G48088,G48089,G48090,G48091,G48092,G48093,G48094,G48095,G48096,G48097,G48098,G48099,G48100,
       G48101,G48102,G48103,G48104,G48105,G48106,G48107,G48108,G48109,G48110,G48111,G48112,G48113,G48114,G48115,G48116,G48117,G48118,G48119,G48120,
       G48121,G48122,G48123,G48124,G48125,G48126,G48127,G48128,G48129,G48130,G48131,G48132,G48133,G48134,G48135,G48136,G48137,G48138,G48139,G48140,
       G48141,G48142,G48143,G48144,G48145,G48146,G48147,G48148,G48149,G48150,G48151,G48152,G48153,G48154,G48155,G48156,G48157,G48158,G48159,G48160,
       G48161,G48162,G48163,G48164,G48165,G48166,G48167,G48168,G48169,G48170,G48171,G48172,G48173,G48174,G48175,G48176,G48177,G48178,G48179,G48180,
       G48181,G48182,G48183,G48184,G48185,G48186,G48187,G48188,G48189,G48190,G48191,G48192,G48193,G48194,G48195,G48196,G48197,G48198,G48199,G48200,
       G48201,G48202,G48203,G48204,G48205,G48206,G48207,G48208,G48209,G48210,G48211,G48212,G48213,G48214,G48215,G48216,G48217,G48218,G48219,G48220,
       G48221,G48222,G48223,G48224,G48225,G48226,G48227,G48228,G48229,G48230,G48231,G48232,G48233,G48234,G48235,G48236,G48237,G48238,G48239,G48240,
       G48241,G48242,G48243,G48244,G48245,G48246,G48247,G48248,G48249,G48250,G48251,G48252,G48253,G48254,G48255,G48256,G48257,G48258,G48259,G48260,
       G48261,G48262,G48263,G48264,G48265,G48266,G48267,G48268,G48269,G48270,G48271,G48272,G48273,G48274,G48275,G48276,G48277,G48278,G48279,G48280,
       G48281,G48282,G48283,G48284,G48285,G48286,G48287,G48288,G48289,G48290,G48291,G48292,G48293,G48294,G48295,G48296,G48297,G48298,G48299,G48300,
       G48301,G48302,G48303,G48304,G48305,G48306,G48307,G48308,G48309,G48310,G48311,G48312,G48313,G48314,G48315,G48316,G48317,G48318,G48319,G48320,
       G48321,G48322,G48323,G48324,G48325,G48326,G48327,G48328,G48329,G48330,G48331,G48332,G48333,G48334,G48335,G48336,G48337,G48338,G48339,G48340,
       G48341,G48342,G48343,G48344,G48345,G48346,G48347,G48348,G48349,G48350,G48351,G48352,G48353,G48354,G48355,G48356,G48357,G48358,G48359,G48360,
       G48361,G48362,G48363,G48364,G48365,G48366,G48367,G48368,G48369,G48370,G48371,G48372,G48373,G48374,G48375,G48376,G48377,G48378,G48379,G48380,
       G48381,G48382,G48383,G48384,G48385,G48386,G48387,G48388,G48389,G48390,G48391,G48392,G48393,G48394,G48395,G48396,G48397,G48398,G48399,G48400,
       G48401,G48402,G48403,G48404,G48405,G48406,G48407,G48408,G48409,G48410,G48411,G48412,G48413,G48414,G48415,G48416,G48417,G48418,G48419,G48420,
       G48421,G48422,G48423,G48424,G48425,G48426,G48427,G48428,G48429,G48430,G48431,G48432,G48433,G48434,G48435,G48436,G48437,G48438,G48439,G48440,
       G48441,G48442,G48443,G48444,G48445,G48446,G48447,G48448,G48449,G48450,G48451,G48452,G48453,G48454,G48455,G48456,G48457,G48458,G48459,G48460,
       G48461,G48462,G48463,G48464,G48465,G48466,G48467,G48468,G48469,G48470,G48471,G48472,G48473,G48474,G48475,G48476,G48477,G48478,G48479,G48480,
       G48481,G48482,G48483,G48484,G48485,G48486,G48487,G48488,G48489,G48490,G48491,G48492,G48493,G48494,G48495,G48496,G48497,G48498,G48499,G48500,
       G48501,G48502,G48503,G48504,G48505,G48506,G48507,G48508,G48509,G48510,G48511,G48512,G48513,G48514,G48515,G48516,G48517,G48518,G48519,G48520,
       G48521,G48522,G48523,G48524,G48525,G48526,G48527,G48528,G48529,G48530,G48531,G48532,G48533,G48534,G48535,G48536,G48537,G48538,G48539,G48540,
       G48541,G48542,G48543,G48544,G48545,G48546,G48547,G48548,G48549,G48550,G48551,G48552,G48553,G48554,G48555,G48556,G48557,G48558,G48559,G48560,
       G48561,G48562,G48563,G48564,G48565,G48566,G48567,G48568,G48569,G48570,G48571,G48572,G48573,G48574,G48575,G48576,G48577,G48578,G48579,G48580,
       G48581,G48582,G48583,G48584,G48585,G48586,G48587,G48588,G48589,G48590,G48591,G48592,G48593,G48594,G48595,G48596,G48597,G48598,G48599,G48600,
       G48601,G48602,G48603,G48604,G48605,G48606,G48607,G48608,G48609,G48610,G48611,G48612,G48613,G48614,G48615,G48616,G48617,G48618,G48619,G48620,
       G48621,G48622,G48623,G48624,G48625,G48626,G48627,G48628,G48629,G48630,G48631,G48632,G48633,G48634,G48635,G48636,G48637,G48638,G48639,G48640,
       G48641,G48642,G48643,G48644,G48645,G48646,G48647,G48648,G48649,G48650,G48651,G48652,G48653,G48654,G48655,G48656,G48657,G48658,G48659,G48660,
       G48661,G48662,G48663,G48664,G48665,G48666,G48667,G48668,G48669,G48670,G48671,G48672,G48673,G48674,G48675,G48676,G48677,G48678,G48679,G48680,
       G48681,G48682,G48683,G48684,G48685,G48686,G48687,G48688,G48689,G48690,G48691,G48692,G48693,G48694,G48695,G48696,G48697,G48698,G48699,G48700,
       G48701,G48702,G48703,G48704,G48705,G48706,G48707,G48708,G48709,G48710,G48711,G48712,G48713,G48714,G48715,G48716,G48717,G48718,G48719,G48720,
       G48721,G48722,G48723,G48724,G48725,G48726,G48727,G48728,G48729,G48730,G48731,G48732,G48733,G48734,G48735,G48736,G48737,G48738,G48739,G48740,
       G48741,G48742,G48743,G48744,G48745,G48746,G48747,G48748,G48749,G48750,G48751,G48752,G48753,G48754,G48755,G48756,G48757,G48758,G48759,G48760,
       G48761,G48762,G48763,G48764,G48765,G48766,G48767,G48768,G48769,G48770,G48771,G48772,G48773,G48774,G48775,G48776,G48777,G48778,G48779,G48780,
       G48781,G48782,G48783,G48784,G48785,G48786,G48787,G48788,G48789,G48790,G48791,G48792,G48793,G48794,G48795,G48796,G48797,G48798,G48799,G48800,
       G48801,G48802,G48803,G48804,G48805,G48806,G48807,G48808,G48809,G48810,G48811,G48812,G48813,G48814,G48815,G48816,G48817,G48818,G48819,G48820,
       G48821,G48822,G48823,G48824,G48825,G48826,G48827,G48828,G48829,G48830,G48831,G48832,G48833,G48834,G48835,G48836,G48837,G48838,G48839,G48840,
       G48841,G48842,G48843,G48844,G48845,G48846,G48847,G48848,G48849,G48850,G48851,G48852,G48853,G48854,G48855,G48856,G48857,G48858,G48859,G48860,
       G48861,G48862,G48863,G48864,G48865,G48866,G48867,G48868,G48869,G48870,G48871,G48872,G48873,G48874,G48875,G48876,G48877,G48878,G48879,G48880,
       G48881,G48882,G48883,G48884,G48885,G48886,G48887,G48888,G48889,G48890,G48891,G48892,G48893,G48894,G48895,G48896,G48897,G48898,G48899,G48900,
       G48901,G48902,G48903,G48904,G48905,G48906,G48907,G48908,G48909,G48910,G48911,G48912,G48913,G48914,G48915,G48916,G48917,G48918,G48919,G48920,
       G48921,G48922,G48923,G48924,G48925,G48926,G48927,G48928,G48929,G48930,G48931,G48932,G48933,G48934,G48935,G48936,G48937,G48938,G48939,G48940,
       G48941,G48942,G48943,G48944,G48945,G48946,G48947,G48948,G48949,G48950,G48951,G48952,G48953,G48954,G48955,G48956,G48957,G48958,G48959,G48960,
       G48961,G48962,G48963,G48964,G48965,G48966,G48967,G48968,G48969,G48970,G48971,G48972,G48973,G48974,G48975,G48976,G48977,G48978,G48979,G48980,
       G48981,G48982,G48983,G48984,G48985,G48986,G48987,G48988,G48989,G48990,G48991,G48992,G48993,G48994,G48995,G48996,G48997,G48998,G48999,G49000,
       G49001,G49002,G49003,G49004,G49005,G49006,G49007,G49008,G49009,G49010,G49011,G49012,G49013,G49014,G49015,G49016,G49017,G49018,G49019,G49020,
       G49021,G49022,G49023,G49024,G49025,G49026,G49027,G49028,G49029,G49030,G49031,G49032,G49033,G49034,G49035,G49036,G49037,G49038,G49039,G49040,
       G49041,G49042,G49043,G49044,G49045,G49046,G49047,G49048,G49049,G49050,G49051,G49052,G49053,G49054,G49055,G49056,G49057,G49058,G49059,G49060,
       G49061,G49062,G49063,G49064,G49065,G49066,G49067,G49068,G49069,G49070,G49071,G49072,G49073,G49074,G49075,G49076,G49077,G49078,G49079,G49080,
       G49081,G49082,G49083,G49084,G49085,G49086,G49087,G49088,G49089,G49090,G49091,G49092,G49093,G49094,G49095,G49096,G49097,G49098,G49099,G49100,
       G49101,G49102,G49103,G49104,G49105,G49106,G49107,G49108,G49109,G49110,G49111,G49112,G49113,G49114,G49115,G49116,G49117,G49118,G49119,G49120,
       G49121,G49122,G49123,G49124,G49125,G49126,G49127,G49128,G49129,G49130,G49131,G49132,G49133,G49134,G49135,G49136,G49137,G49138,G49139,G49140,
       G49141,G49142,G49143,G49144,G49145,G49146,G49147,G49148,G49149,G49150,G49151,G49152,G49153,G49154,G49155,G49156,G49157,G49158,G49159,G49160,
       G49161,G49162,G49163,G49164,G49165,G49166,G49167,G49168,G49169,G49170,G49171,G49172,G49173,G49174,G49175,G49176,G49177,G49178,G49179,G49180,
       G49181,G49182,G49183,G49184,G49185,G49186,G49187,G49188,G49189,G49190,G49191,G49192,G49193,G49194,G49195,G49196,G49197,G49198,G49199,G49200,
       G49201,G49202,G49203,G49204,G49205,G49206,G49207,G49208,G49209,G49210,G49211,G49212,G49213,G49214,G49215,G49216,G49217,G49218,G49219,G49220,
       G49221,G49222,G49223,G49224,G49225,G49226,G49227,G49228,G49229,G49230,G49231,G49232,G49233,G49234,G49235,G49236,G49237,G49238,G49239,G49240,
       G49241,G49242,G49243,G49244,G49245,G49246,G49247,G49248,G49249,G49250,G49251,G49252,G49253,G49254,G49255,G49256,G49257,G49258,G49259,G49260,
       G49261,G49262,G49263,G49264,G49265,G49266,G49267,G49268,G49269,G49270,G49271,G49272,G49273,G49274,G49275,G49276,G49277,G49278,G49279,G49280,
       G49281,G49282,G49283,G49284,G49285,G49286,G49287,G49288,G49289,G49290,G49291,G49292,G49293,G49294,G49295,G49296,G49297,G49298,G49299,G49300,
       G49301,G49302,G49303,G49304,G49305,G49306,G49307,G49308,G49309,G49310,G49311,G49312,G49313,G49314,G49315,G49316,G49317,G49318,G49319,G49320,
       G49321,G49322,G49323,G49324,G49325,G49326,G49327,G49328,G49329,G49330,G49331,G49332,G49333,G49334,G49335,G49336,G49337,G49338,G49339,G49340,
       G49341,G49342,G49343,G49344,G49345,G49346,G49347,G49348,G49349,G49350,G49351,G49352,G49353,G49354,G49355,G49356,G49357,G49358,G49359,G49360,
       G49361,G49362,G49363,G49364,G49365,G49366,G49367,G49368,G49369,G49370,G49371,G49372,G49373,G49374,G49375,G49376,G49377,G49378,G49379,G49380,
       G49381,G49382,G49383,G49384,G49385,G49386,G49387,G49388,G49389,G49390,G49391,G49392,G49393,G49394,G49395,G49396,G49397,G49398,G49399,G49400,
       G49401,G49402,G49403,G49404,G49405,G49406,G49407,G49408,G49409,G49410,G49411,G49412,G49413,G49414,G49415,G49416,G49417,G49418,G49419,G49420,
       G49421,G49422,G49423,G49424,G49425,G49426,G49427,G49428,G49429,G49430,G49431,G49432,G49433,G49434,G49435,G49436,G49437,G49438,G49439,G49440,
       G49441,G49442,G49443,G49444,G49445,G49446,G49447,G49448,G49449,G49450,G49451,G49452,G49453,G49454,G49455,G49456,G49457,G49458,G49459,G49460,
       G49461,G49462,G49463,G49464,G49465,G49466,G49467,G49468,G49469,G49470,G49471,G49472,G49473,G49474,G49475,G49476,G49477,G49478,G49479,G49480,
       G49481,G49482,G49483,G49484,G49485,G49486,G49487,G49488,G49489,G49490,G49491,G49492,G49493,G49494,G49495,G49496,G49497,G49498,G49499,G49500,
       G49501,G49502,G49503,G49504,G49505,G49506,G49507,G49508,G49509,G49510,G49511,G49512,G49513,G49514,G49515,G49516,G49517,G49518,G49519,G49520,
       G49521,G49522,G49523,G49524,G49525,G49526,G49527,G49528,G49529,G49530,G49531,G49532,G49533,G49534,G49535,G49536,G49537,G49538,G49539,G49540,
       G49541,G49542,G49543,G49544,G49545,G49546,G49547,G49548,G49549,G49550,G49551,G49552,G49553,G49554,G49555,G49556,G49557,G49558,G49559,G49560,
       G49561,G49562,G49563,G49564,G49565,G49566,G49567,G49568,G49569,G49570,G49571,G49572,G49573,G49574,G49575,G49576,G49577,G49578,G49579,G49580,
       G49581,G49582,G49583,G49584,G49585,G49586,G49587,G49588,G49589,G49590,G49591,G49592,G49593,G49594,G49595,G49596,G49597,G49598,G49599,G49600,
       G49601,G49602,G49603,G49604,G49605,G49606,G49607,G49608,G49609,G49610,G49611,G49612,G49613,G49614,G49615,G49616,G49617,G49618,G49619,G49620,
       G49621,G49622,G49623,G49624,G49625,G49626,G49627,G49628,G49629,G49630,G49631,G49632,G49633,G49634,G49635,G49636,G49637,G49638,G49639,G49640,
       G49641,G49642,G49643,G49644,G49645,G49646,G49647,G49648,G49649,G49650,G49651,G49652,G49653,G49654,G49655,G49656,G49657,G49658,G49659,G49660,
       G49661,G49662,G49663,G49664,G49665,G49666,G49667,G49668,G49669,G49670,G49671,G49672,G49673,G49674,G49675,G49676,G49677,G49678,G49679,G49680,
       G49681,G49682,G49683,G49684,G49685,G49686,G49687,G49688,G49689,G49690,G49691,G49692,G49693,G49694,G49695,G49696,G49697,G49698,G49699,G49700,
       G49701,G49702,G49703,G49704,G49705,G49706,G49707,G49708,G49709,G49710,G49711,G49712,G49713,G49714,G49715,G49716,G49717,G49718,G49719,G49720,
       G49721,G49722,G49723,G49724,G49725,G49726,G49727,G49728,G49729,G49730,G49731,G49732,G49733,G49734,G49735,G49736,G49737,G49738,G49739,G49740,
       G49741,G49742,G49743,G49744,G49745,G49746,G49747,G49748,G49749,G49750,G49751,G49752,G49753,G49754,G49755,G49756,G49757,G49758,G49759,G49760,
       G49761,G49762,G49763,G49764,G49765,G49766,G49767,G49768,G49769,G49770,G49771,G49772,G49773,G49774,G49775,G49776,G49777,G49778,G49779,G49780,
       G49781,G49782,G49783,G49784,G49785,G49786,G49787,G49788,G49789,G49790,G49791,G49792,G49793,G49794,G49795,G49796,G49797,G49798,G49799,G49800,
       G49801,G49802,G49803,G49804,G49805,G49806,G49807,G49808,G49809,G49810,G49811,G49812,G49813,G49814,G49815,G49816,G49817,G49818,G49819,G49820,
       G49821,G49822,G49823,G49824,G49825,G49826,G49827,G49828,G49829,G49830,G49831,G49832,G49833,G49834,G49835,G49836,G49837,G49838,G49839,G49840,
       G49841,G49842,G49843,G49844,G49845,G49846,G49847,G49848,G49849,G49850,G49851,G49852,G49853,G49854,G49855,G49856,G49857,G49858,G49859,G49860,
       G49861,G49862,G49863,G49864,G49865,G49866,G49867,G49868,G49869,G49870,G49871,G49872,G49873,G49874,G49875,G49876,G49877,G49878,G49879,G49880,
       G49881,G49882,G49883,G49884,G49885,G49886,G49887,G49888,G49889,G49890,G49891,G49892,G49893,G49894,G49895,G49896,G49897,G49898,G49899,G49900,
       G49901,G49902,G49903,G49904,G49905,G49906,G49907,G49908,G49909,G49910,G49911,G49912,G49913,G49914,G49915,G49916,G49917,G49918,G49919,G49920,
       G49921,G49922,G49923,G49924,G49925,G49926,G49927,G49928,G49929,G49930,G49931,G49932,G49933,G49934,G49935,G49936,G49937,G49938,G49939,G49940,
       G49941,G49942,G49943,G49944,G49945,G49946,G49947,G49948,G49949,G49950,G49951,G49952,G49953,G49954,G49955,G49956,G49957,G49958,G49959,G49960,
       G49961,G49962,G49963,G49964,G49965,G49966,G49967,G49968,G49969,G49970,G49971,G49972,G49973,G49974,G49975,G49976,G49977,G49978,G49979,G49980,
       G49981,G49982,G49983,G49984,G49985,G49986,G49987,G49988,G49989,G49990,G49991,G49992,G49993,G49994,G49995,G49996,G49997,G49998,G49999,G50000,
       G50001,G50002,G50003,G50004,G50005,G50006,G50007,G50008,G50009,G50010,G50011,G50012,G50013,G50014,G50015,G50016,G50017,G50018,G50019,G50020,
       G50021,G50022,G50023,G50024,G50025,G50026,G50027,G50028,G50029,G50030,G50031,G50032,G50033,G50034,G50035,G50036,G50037,G50038,G50039,G50040,
       G50041,G50042,G50043,G50044,G50045,G50046,G50047,G50048,G50049,G50050,G50051,G50052,G50053,G50054,G50055,G50056,G50057,G50058,G50059,G50060,
       G50061,G50062,G50063,G50064,G50065,G50066,G50067,G50068,G50069,G50070,G50071,G50072,G50073,G50074,G50075,G50076,G50077,G50078,G50079,G50080,
       G50081,G50082,G50083,G50084,G50085,G50086,G50087,G50088,G50089,G50090,G50091,G50092,G50093,G50094,G50095,G50096,G50097,G50098,G50099,G50100,
       G50101,G50102,G50103,G50104,G50105,G50106,G50107,G50108,G50109,G50110,G50111,G50112,G50113,G50114,G50115,G50116,G50117,G50118,G50119,G50120,
       G50121,G50122,G50123,G50124,G50125,G50126,G50127,G50128,G50129,G50130,G50131,G50132,G50133,G50134,G50135,G50136,G50137,G50138,G50139,G50140,
       G50141,G50142,G50143,G50144,G50145,G50146,G50147,G50148,G50149,G50150,G50151,G50152,G50153,G50154,G50155,G50156,G50157,G50158,G50159,G50160,
       G50161,G50162,G50163,G50164,G50165,G50166,G50167,G50168,G50169,G50170,G50171,G50172,G50173,G50174,G50175,G50176,G50177,G50178,G50179,G50180,
       G50181,G50182,G50183,G50184,G50185,G50186,G50187,G50188,G50189,G50190,G50191,G50192,G50193,G50194,G50195,G50196,G50197,G50198,G50199,G50200,
       G50201,G50202,G50203,G50204,G50205,G50206,G50207,G50208,G50209,G50210,G50211,G50212,G50213,G50214,G50215,G50216,G50217,G50218,G50219,G50220,
       G50221,G50222,G50223,G50224,G50225,G50226,G50227,G50228,G50229,G50230,G50231,G50232,G50233,G50234,G50235,G50236,G50237,G50238,G50239,G50240,
       G50241,G50242,G50243,G50244,G50245,G50246,G50247,G50248,G50249,G50250,G50251,G50252,G50253,G50254,G50255,G50256,G50257,G50258,G50259,G50260,
       G50261,G50262,G50263,G50264,G50265,G50266,G50267,G50268,G50269,G50270,G50271,G50272,G50273,G50274,G50275,G50276,G50277,G50278,G50279,G50280,
       G50281,G50282,G50283,G50284,G50285,G50286,G50287,G50288,G50289,G50290,G50291,G50292,G50293,G50294,G50295,G50296,G50297,G50298,G50299,G50300,
       G50301,G50302,G50303,G50304,G50305,G50306,G50307,G50308,G50309,G50310,G50311,G50312,G50313,G50314,G50315,G50316,G50317,G50318,G50319,G50320,
       G50321,G50322,G50323,G50324,G50325,G50326,G50327,G50328,G50329,G50330,G50331,G50332,G50333,G50334,G50335,G50336,G50337,G50338,G50339,G50340,
       G50341,G50342,G50343,G50344,G50345,G50346,G50347,G50348,G50349,G50350,G50351,G50352,G50353,G50354,G50355,G50356,G50357,G50358,G50359,G50360,
       G50361,G50362,G50363,G50364,G50365,G50366,G50367,G50368,G50369,G50370,G50371,G50372,G50373,G50374,G50375,G50376,G50377,G50378,G50379,G50380,
       G50381,G50382,G50383,G50384,G50385,G50386,G50387,G50388,G50389,G50390,G50391,G50392,G50393,G50394,G50395,G50396,G50397,G50398,G50399,G50400,
       G50401,G50402,G50403,G50404,G50405,G50406,G50407,G50408,G50409,G50410,G50411,G50412,G50413,G50414,G50415,G50416,G50417,G50418,G50419,G50420,
       G50421,G50422,G50423,G50424,G50425,G50426,G50427,G50428,G50429,G50430,G50431,G50432,G50433,G50434,G50435,G50436,G50437,G50438,G50439,G50440,
       G50441,G50442,G50443,G50444,G50445,G50446,G50447,G50448,G50449,G50450,G50451,G50452,G50453,G50454,G50455,G50456,G50457,G50458,G50459,G50460,
       G50461,G50462,G50463,G50464,G50465,G50466,G50467,G50468,G50469,G50470,G50471,G50472,G50473,G50474,G50475,G50476,G50477,G50478,G50479,G50480,
       G50481,G50482,G50483,G50484,G50485,G50486,G50487,G50488,G50489,G50490,G50491,G50492,G50493,G50494,G50495,G50496,G50497,G50498,G50499,G50500,
       G50501,G50502,G50503,G50504,G50505,G50506,G50507,G50508,G50509,G50510,G50511,G50512,G50513,G50514,G50515,G50516,G50517,G50518,G50519,G50520,
       G50521,G50522,G50523,G50524,G50525,G50526,G50527,G50528,G50529,G50530,G50531,G50532,G50533,G50534,G50535,G50536,G50537,G50538,G50539,G50540,
       G50541,G50542,G50543,G50544,G50545,G50546,G50547,G50548,G50549,G50550,G50551,G50552,G50553,G50554,G50555,G50556,G50557,G50558,G50559,G50560,
       G50561,G50562,G50563,G50564,G50565,G50566,G50567,G50568,G50569,G50570,G50571,G50572,G50573,G50574,G50575,G50576,G50577,G50578,G50579,G50580,
       G50581,G50582,G50583,G50584,G50585,G50586,G50587,G50588,G50589,G50590,G50591,G50592,G50593,G50594,G50595,G50596,G50597,G50598,G50599,G50600,
       G50601,G50602,G50603,G50604,G50605,G50606,G50607,G50608,G50609,G50610,G50611,G50612,G50613,G50614,G50615,G50616,G50617,G50618,G50619,G50620,
       G50621,G50622,G50623,G50624,G50625,G50626,G50627,G50628,G50629,G50630,G50631,G50632,G50633,G50634,G50635,G50636,G50637,G50638,G50639,G50640,
       G50641,G50642,G50643,G50644,G50645,G50646,G50647,G50648,G50649,G50650,G50651,G50652,G50653,G50654,G50655,G50656,G50657,G50658,G50659,G50660,
       G50661,G50662,G50663,G50664,G50665,G50666,G50667,G50668,G50669,G50670,G50671,G50672,G50673,G50674,G50675,G50676,G50677,G50678,G50679,G50680,
       G50681,G50682,G50683,G50684,G50685,G50686,G50687,G50688,G50689,G50690,G50691,G50692,G50693,G50694,G50695,G50696,G50697,G50698,G50699,G50700,
       G50701,G50702,G50703,G50704,G50705,G50706,G50707,G50708,G50709,G50710,G50711,G50712,G50713,G50714,G50715,G50716,G50717,G50718,G50719,G50720,
       G50721,G50722,G50723,G50724,G50725,G50726,G50727,G50728,G50729,G50730,G50731,G50732,G50733,G50734,G50735,G50736,G50737,G50738,G50739,G50740,
       G50741,G50742,G50743,G50744,G50745,G50746,G50747,G50748,G50749,G50750,G50751,G50752,G50753,G50754,G50755,G50756,G50757,G50758,G50759,G50760,
       G50761,G50762,G50763,G50764,G50765,G50766,G50767,G50768,G50769,G50770,G50771,G50772,G50773,G50774,G50775,G50776,G50777,G50778,G50779,G50780,
       G50781,G50782,G50783,G50784,G50785,G50786,G50787,G50788,G50789,G50790,G50791,G50792,G50793,G50794,G50795,G50796,G50797,G50798,G50799,G50800,
       G50801,G50802,G50803,G50804,G50805,G50806,G50807,G50808,G50809,G50810,G50811,G50812,G50813,G50814,G50815,G50816,G50817,G50818,G50819,G50820,
       G50821,G50822,G50823,G50824,G50825,G50826,G50827,G50828,G50829,G50830,G50831,G50832,G50833,G50834,G50835,G50836,G50837,G50838,G50839,G50840,
       G50841,G50842,G50843,G50844,G50845,G50846,G50847,G50848,G50849,G50850,G50851,G50852,G50853,G50854,G50855,G50856,G50857,G50858,G50859,G50860,
       G50861,G50862,G50863,G50864,G50865,G50866,G50867,G50868,G50869,G50870,G50871,G50872,G50873,G50874,G50875,G50876,G50877,G50878,G50879,G50880,
       G50881,G50882,G50883,G50884,G50885,G50886,G50887,G50888,G50889,G50890,G50891,G50892,G50893,G50894,G50895,G50896,G50897,G50898,G50899,G50900,
       G50901,G50902,G50903,G50904,G50905,G50906,G50907,G50908,G50909,G50910,G50911,G50912,G50913,G50914,G50915,G50916,G50917,G50918,G50919,G50920,
       G50921,G50922,G50923,G50924,G50925,G50926,G50927,G50928,G50929,G50930,G50931,G50932,G50933,G50934,G50935,G50936,G50937,G50938,G50939,G50940,
       G50941,G50942,G50943,G50944,G50945,G50946,G50947,G50948,G50949,G50950,G50951,G50952,G50953,G50954,G50955,G50956,G50957,G50958,G50959,G50960,
       G50961,G50962,G50963,G50964,G50965,G50966,G50967,G50968,G50969,G50970,G50971,G50972,G50973,G50974,G50975,G50976,G50977,G50978,G50979,G50980,
       G50981,G50982,G50983,G50984,G50985,G50986,G50987,G50988,G50989,G50990,G50991,G50992,G50993,G50994,G50995,G50996,G50997,G50998,G50999,G51000,
       G51001,G51002,G51003,G51004,G51005,G51006,G51007,G51008,G51009,G51010,G51011,G51012,G51013,G51014,G51015,G51016,G51017,G51018,G51019,G51020,
       G51021,G51022,G51023,G51024,G51025,G51026,G51027,G51028,G51029,G51030,G51031,G51032,G51033,G51034,G51035,G51036,G51037,G51038,G51039,G51040,
       G51041,G51042,G51043,G51044,G51045,G51046,G51047,G51048,G51049,G51050,G51051,G51052,G51053,G51054,G51055,G51056,G51057,G51058,G51059,G51060,
       G51061,G51062,G51063,G51064,G51065,G51066,G51067,G51068,G51069,G51070,G51071,G51072,G51073,G51074,G51075,G51076,G51077,G51078,G51079,G51080,
       G51081,G51082,G51083,G51084,G51085,G51086,G51087,G51088,G51089,G51090,G51091,G51092,G51093,G51094,G51095,G51096,G51097,G51098,G51099,G51100,
       G51101,G51102,G51103,G51104,G51105,G51106,G51107,G51108,G51109,G51110,G51111,G51112,G51113,G51114,G51115,G51116,G51117,G51118,G51119,G51120,
       G51121,G51122,G51123,G51124,G51125,G51126,G51127,G51128,G51129,G51130,G51131,G51132,G51133,G51134,G51135,G51136,G51137,G51138,G51139,G51140,
       G51141,G51142,G51143,G51144,G51145,G51146,G51147,G51148,G51149,G51150,G51151,G51152,G51153,G51154,G51155,G51156,G51157,G51158,G51159,G51160,
       G51161,G51162,G51163,G51164,G51165,G51166,G51167,G51168,G51169,G51170,G51171,G51172,G51173,G51174,G51175,G51176,G51177,G51178,G51179,G51180,
       G51181,G51182,G51183,G51184,G51185,G51186,G51187,G51188,G51189,G51190,G51191,G51192,G51193,G51194,G51195,G51196,G51197,G51198,G51199,G51200,
       G51201,G51202,G51203,G51204,G51205,G51206,G51207,G51208,G51209,G51210,G51211,G51212,G51213,G51214,G51215,G51216,G51217,G51218,G51219,G51220,
       G51221,G51222,G51223,G51224,G51225,G51226,G51227,G51228,G51229,G51230,G51231,G51232,G51233,G51234,G51235,G51236,G51237,G51238,G51239,G51240,
       G51241,G51242,G51243,G51244,G51245,G51246,G51247,G51248,G51249,G51250,G51251,G51252,G51253,G51254,G51255,G51256,G51257,G51258,G51259,G51260,
       G51261,G51262,G51263,G51264,G51265,G51266,G51267,G51268,G51269,G51270,G51271,G51272,G51273,G51274,G51275,G51276,G51277,G51278,G51279,G51280,
       G51281,G51282,G51283,G51284,G51285,G51286,G51287,G51288,G51289,G51290,G51291,G51292,G51293,G51294,G51295,G51296,G51297,G51298,G51299,G51300,
       G51301,G51302,G51303,G51304,G51305,G51306,G51307,G51308,G51309,G51310,G51311,G51312,G51313,G51314,G51315,G51316,G51317,G51318,G51319,G51320,
       G51321,G51322,G51323,G51324,G51325,G51326,G51327,G51328,G51329,G51330,G51331,G51332,G51333,G51334,G51335,G51336,G51337,G51338,G51339,G51340,
       G51341,G51342,G51343,G51344,G51345,G51346,G51347,G51348,G51349,G51350,G51351,G51352,G51353,G51354,G51355,G51356,G51357,G51358,G51359,G51360,
       G51361,G51362,G51363,G51364,G51365,G51366,G51367,G51368,G51369,G51370,G51371,G51372,G51373,G51374,G51375,G51376,G51377,G51378,G51379,G51380,
       G51381,G51382,G51383,G51384,G51385,G51386,G51387,G51388,G51389,G51390,G51391,G51392,G51393,G51394,G51395,G51396,G51397,G51398,G51399,G51400,
       G51401,G51402,G51403,G51404,G51405,G51406,G51407,G51408,G51409,G51410,G51411,G51412,G51413,G51414,G51415,G51416,G51417,G51418,G51419,G51420,
       G51421,G51422,G51423,G51424,G51425,G51426,G51427,G51428,G51429,G51430,G51431,G51432,G51433,G51434,G51435,G51436,G51437,G51438,G51439,G51440,
       G51441,G51442,G51443,G51444,G51445,G51446,G51447,G51448,G51449,G51450,G51451,G51452,G51453,G51454,G51455,G51456,G51457,G51458,G51459,G51460,
       G51461,G51462,G51463,G51464,G51465,G51466,G51467,G51468,G51469,G51470,G51471,G51472,G51473,G51474,G51475,G51476,G51477,G51478,G51479,G51480,
       G51481,G51482,G51483,G51484,G51485,G51486,G51487,G51488,G51489,G51490,G51491,G51492,G51493,G51494,G51495,G51496,G51497,G51498,G51499,G51500,
       G51501,G51502,G51503,G51504,G51505,G51506,G51507,G51508,G51509,G51510,G51511,G51512,G51513,G51514,G51515,G51516,G51517,G51518,G51519,G51520,
       G51521,G51522,G51523,G51524,G51525,G51526,G51527,G51528,G51529,G51530,G51531,G51532,G51533,G51534,G51535,G51536,G51537,G51538,G51539,G51540,
       G51541,G51542,G51543,G51544,G51545,G51546,G51547,G51548,G51549,G51550,G51551,G51552,G51553,G51554,G51555,G51556,G51557,G51558,G51559,G51560,
       G51561,G51562,G51563,G51564,G51565,G51566,G51567,G51568,G51569,G51570,G51571,G51572,G51573,G51574,G51575,G51576,G51577,G51578,G51579,G51580,
       G51581,G51582,G51583,G51584,G51585,G51586,G51587,G51588,G51589,G51590,G51591,G51592,G51593,G51594,G51595,G51596,G51597,G51598,G51599,G51600,
       G51601,G51602,G51603,G51604,G51605,G51606,G51607,G51608,G51609,G51610,G51611,G51612,G51613,G51614,G51615,G51616,G51617,G51618,G51619,G51620,
       G51621,G51622,G51623,G51624,G51625,G51626,G51627,G51628,G51629,G51630,G51631,G51632,G51633,G51634,G51635,G51636,G51637,G51638,G51639,G51640,
       G51641,G51642,G51643,G51644,G51645,G51646,G51647,G51648,G51649,G51650,G51651,G51652,G51653,G51654,G51655,G51656,G51657,G51658,G51659,G51660,
       G51661,G51662,G51663,G51664,G51665,G51666,G51667,G51668,G51669,G51670,G51671,G51672,G51673,G51674,G51675,G51676,G51677,G51678,G51679,G51680,
       G51681,G51682,G51683,G51684,G51685,G51686,G51687,G51688,G51689,G51690,G51691,G51692,G51693,G51694,G51695,G51696,G51697,G51698,G51699,G51700,
       G51701,G51702,G51703,G51704,G51705,G51706,G51707,G51708,G51709,G51710,G51711,G51712,G51713,G51714,G51715,G51716,G51717,G51718,G51719,G51720,
       G51721,G51722,G51723,G51724,G51725,G51726,G51727,G51728,G51729,G51730,G51731,G51732,G51733,G51734,G51735,G51736,G51737,G51738,G51739,G51740,
       G51741,G51742,G51743,G51744,G51745,G51746,G51747,G51748,G51749,G51750,G51751,G51752,G51753,G51754,G51755,G51756,G51757,G51758,G51759,G51760,
       G51761,G51762,G51763,G51764,G51765,G51766,G51767,G51768,G51769,G51770,G51771,G51772,G51773,G51774,G51775,G51776,G51777,G51778,G51779,G51780,
       G51781,G51782,G51783,G51784,G51785,G51786,G51787,G51788,G51789,G51790,G51791,G51792,G51793,G51794,G51795,G51796,G51797,G51798,G51799,G51800,
       G51801,G51802,G51803,G51804,G51805,G51806,G51807,G51808,G51809,G51810,G51811,G51812,G51813,G51814,G51815,G51816,G51817,G51818,G51819,G51820,
       G51821,G51822,G51823,G51824,G51825,G51826,G51827,G51828,G51829,G51830,G51831,G51832,G51833,G51834,G51835,G51836,G51837,G51838,G51839,G51840,
       G51841,G51842,G51843,G51844,G51845,G51846,G51847,G51848,G51849,G51850,G51851,G51852,G51853,G51854,G51855,G51856,G51857,G51858,G51859,G51860,
       G51861,G51862,G51863,G51864,G51865,G51866,G51867,G51868,G51869,G51870,G51871,G51872,G51873,G51874,G51875,G51876,G51877,G51878,G51879,G51880,
       G51881,G51882,G51883,G51884,G51885,G51886,G51887,G51888,G51889,G51890,G51891,G51892,G51893,G51894,G51895,G51896,G51897,G51898,G51899,G51900,
       G51901,G51902,G51903,G51904,G51905,G51906,G51907,G51908,G51909,G51910,G51911,G51912,G51913,G51914,G51915,G51916,G51917,G51918,G51919,G51920,
       G51921,G51922,G51923,G51924,G51925,G51926,G51927,G51928,G51929,G51930,G51931,G51932,G51933,G51934,G51935,G51936,G51937,G51938,G51939,G51940,
       G51941,G51942,G51943,G51944,G51945,G51946,G51947,G51948,G51949,G51950,G51951,G51952,G51953,G51954,G51955,G51956,G51957,G51958,G51959,G51960,
       G51961,G51962,G51963,G51964,G51965,G51966,G51967,G51968,G51969,G51970,G51971,G51972,G51973,G51974,G51975,G51976,G51977,G51978,G51979,G51980,
       G51981,G51982,G51983,G51984,G51985,G51986,G51987,G51988,G51989,G51990,G51991,G51992,G51993,G51994,G51995,G51996,G51997,G51998,G51999,G52000,
       G52001,G52002,G52003,G52004,G52005,G52006,G52007,G52008,G52009,G52010,G52011,G52012,G52013,G52014,G52015,G52016,G52017,G52018,G52019,G52020,
       G52021,G52022,G52023,G52024,G52025,G52026,G52027,G52028,G52029,G52030,G52031,G52032,G52033,G52034,G52035,G52036,G52037,G52038,G52039,G52040,
       G52041,G52042,G52043,G52044,G52045,G52046,G52047,G52048,G52049,G52050,G52051,G52052,G52053,G52054,G52055,G52056,G52057,G52058,G52059,G52060,
       G52061,G52062,G52063,G52064,G52065,G52066,G52067,G52068,G52069,G52070,G52071,G52072,G52073,G52074,G52075,G52076,G52077,G52078,G52079,G52080,
       G52081,G52082,G52083,G52084,G52085,G52086,G52087,G52088,G52089,G52090,G52091,G52092,G52093,G52094,G52095,G52096,G52097,G52098,G52099,G52100,
       G52101,G52102,G52103,G52104,G52105,G52106,G52107,G52108,G52109,G52110,G52111,G52112,G52113,G52114,G52115,G52116,G52117,G52118,G52119,G52120,
       G52121,G52122,G52123,G52124,G52125,G52126,G52127,G52128,G52129,G52130,G52131,G52132,G52133,G52134,G52135,G52136,G52137,G52138,G52139,G52140,
       G52141,G52142,G52143,G52144,G52145,G52146,G52147,G52148,G52149,G52150,G52151,G52152,G52153,G52154,G52155,G52156,G52157,G52158,G52159,G52160,
       G52161,G52162,G52163,G52164,G52165,G52166,G52167,G52168,G52169,G52170,G52171,G52172,G52173,G52174,G52175,G52176,G52177,G52178,G52179,G52180,
       G52181,G52182,G52183,G52184,G52185,G52186,G52187,G52188,G52189,G52190,G52191,G52192,G52193,G52194,G52195,G52196,G52197,G52198,G52199,G52200,
       G52201,G52202,G52203,G52204,G52205,G52206,G52207,G52208,G52209,G52210,G52211,G52212,G52213,G52214,G52215,G52216,G52217,G52218,G52219,G52220,
       G52221,G52222,G52223,G52224,G52225,G52226,G52227,G52228,G52229,G52230,G52231,G52232,G52233,G52234,G52235,G52236,G52237,G52238,G52239,G52240,
       G52241,G52242,G52243,G52244,G52245,G52246,G52247,G52248,G52249,G52250,G52251,G52252,G52253,G52254,G52255,G52256,G52257,G52258,G52259,G52260,
       G52261,G52262,G52263,G52264,G52265,G52266,G52267,G52268,G52269,G52270,G52271,G52272,G52273,G52274,G52275,G52276,G52277,G52278,G52279,G52280,
       G52281,G52282,G52283,G52284,G52285,G52286,G52287,G52288,G52289,G52290,G52291,G52292,G52293,G52294,G52295,G52296,G52297,G52298,G52299,G52300,
       G52301,G52302,G52303,G52304,G52305,G52306,G52307,G52308,G52309,G52310,G52311,G52312,G52313,G52314,G52315,G52316,G52317,G52318,G52319,G52320,
       G52321,G52322,G52323,G52324,G52325,G52326,G52327,G52328,G52329,G52330,G52331,G52332,G52333,G52334,G52335,G52336,G52337,G52338,G52339,G52340,
       G52341,G52342,G52343,G52344,G52345,G52346,G52347,G52348,G52349,G52350,G52351,G52352,G52353,G52354,G52355,G52356,G52357,G52358,G52359,G52360,
       G52361,G52362,G52363,G52364,G52365,G52366,G52367,G52368,G52369,G52370,G52371,G52372,G52373,G52374,G52375,G52376,G52377,G52378,G52379,G52380,
       G52381,G52382,G52383,G52384,G52385,G52386,G52387,G52388,G52389,G52390,G52391,G52392,G52393,G52394,G52395,G52396,G52397,G52398,G52399,G52400,
       G52401,G52402,G52403,G52404,G52405,G52406,G52407,G52408,G52409,G52410,G52411,G52412,G52413,G52414,G52415,G52416,G52417,G52418,G52419,G52420,
       G52421,G52422,G52423,G52424,G52425,G52426,G52427,G52428,G52429,G52430,G52431,G52432,G52433,G52434,G52435,G52436,G52437,G52438,G52439,G52440,
       G52441,G52442,G52443,G52444,G52445,G52446,G52447,G52448,G52449,G52450,G52451,G52452,G52453,G52454,G52455,G52456,G52457,G52458,G52459,G52460,
       G52461,G52462,G52463,G52464,G52465,G52466,G52467,G52468,G52469,G52470,G52471,G52472,G52473,G52474,G52475,G52476,G52477,G52478,G52479,G52480,
       G52481,G52482,G52483,G52484,G52485,G52486,G52487,G52488,G52489,G52490,G52491,G52492,G52493,G52494,G52495,G52496,G52497,G52498,G52499,G52500,
       G52501,G52502,G52503,G52504,G52505,G52506,G52507,G52508,G52509,G52510,G52511,G52512,G52513,G52514,G52515,G52516,G52517,G52518,G52519,G52520,
       G52521,G52522,G52523,G52524,G52525,G52526,G52527,G52528,G52529,G52530,G52531,G52532,G52533,G52534,G52535,G52536,G52537,G52538,G52539,G52540,
       G52541,G52542,G52543,G52544,G52545,G52546,G52547,G52548,G52549,G52550,G52551,G52552,G52553,G52554,G52555,G52556,G52557,G52558,G52559,G52560,
       G52561,G52562,G52563,G52564,G52565,G52566,G52567,G52568,G52569,G52570,G52571,G52572,G52573,G52574,G52575,G52576,G52577,G52578,G52579,G52580,
       G52581,G52582,G52583,G52584,G52585,G52586,G52587,G52588,G52589,G52590,G52591,G52592,G52593,G52594,G52595,G52596,G52597,G52598,G52599,G52600,
       G52601,G52602,G52603,G52604,G52605,G52606,G52607,G52608,G52609,G52610,G52611,G52612,G52613,G52614,G52615,G52616,G52617,G52618,G52619,G52620,
       G52621,G52622,G52623,G52624,G52625,G52626,G52627,G52628,G52629,G52630,G52631,G52632,G52633,G52634,G52635,G52636,G52637,G52638,G52639,G52640,
       G52641,G52642,G52643,G52644,G52645,G52646,G52647,G52648,G52649,G52650,G52651,G52652,G52653,G52654,G52655,G52656,G52657,G52658,G52659,G52660,
       G52661,G52662,G52663,G52664,G52665,G52666,G52667,G52668,G52669,G52670,G52671,G52672,G52673,G52674,G52675,G52676,G52677,G52678,G52679,G52680,
       G52681,G52682,G52683,G52684,G52685,G52686,G52687,G52688,G52689,G52690,G52691,G52692,G52693,G52694,G52695,G52696,G52697,G52698,G52699,G52700,
       G52701,G52702,G52703,G52704,G52705,G52706,G52707,G52708,G52709,G52710,G52711,G52712,G52713,G52714,G52715,G52716,G52717,G52718,G52719,G52720,
       G52721,G52722,G52723,G52724,G52725,G52726,G52727,G52728,G52729,G52730,G52731,G52732,G52733,G52734,G52735,G52736,G52737,G52738,G52739,G52740,
       G52741,G52742,G52743,G52744,G52745,G52746,G52747,G52748,G52749,G52750,G52751,G52752,G52753,G52754,G52755,G52756,G52757,G52758,G52759,G52760,
       G52761,G52762,G52763,G52764,G52765,G52766,G52767,G52768,G52769,G52770,G52771,G52772,G52773,G52774,G52775,G52776,G52777,G52778,G52779,G52780,
       G52781,G52782,G52783,G52784,G52785,G52786,G52787,G52788,G52789,G52790,G52791,G52792,G52793,G52794,G52795,G52796,G52797,G52798,G52799,G52800,
       G52801,G52802,G52803,G52804,G52805,G52806,G52807,G52808,G52809,G52810,G52811,G52812,G52813,G52814,G52815,G52816,G52817,G52818,G52819,G52820,
       G52821,G52822,G52823,G52824,G52825,G52826,G52827,G52828,G52829,G52830,G52831,G52832,G52833,G52834,G52835,G52836,G52837,G52838,G52839,G52840,
       G52841,G52842,G52843,G52844,G52845,G52846,G52847,G52848,G52849,G52850,G52851,G52852,G52853,G52854,G52855,G52856,G52857,G52858,G52859,G52860,
       G52861,G52862,G52863,G52864,G52865,G52866,G52867,G52868,G52869,G52870,G52871,G52872,G52873,G52874,G52875,G52876,G52877,G52878,G52879,G52880,
       G52881,G52882,G52883,G52884,G52885,G52886,G52887,G52888,G52889,G52890,G52891,G52892,G52893,G52894,G52895,G52896,G52897,G52898,G52899,G52900,
       G52901,G52902,G52903,G52904,G52905,G52906,G52907,G52908,G52909,G52910,G52911,G52912,G52913,G52914,G52915,G52916,G52917,G52918,G52919,G52920,
       G52921,G52922,G52923,G52924,G52925,G52926,G52927,G52928,G52929,G52930,G52931,G52932,G52933,G52934,G52935,G52936,G52937,G52938,G52939,G52940,
       G52941,G52942,G52943,G52944,G52945,G52946,G52947,G52948,G52949,G52950,G52951,G52952,G52953,G52954,G52955,G52956,G52957,G52958,G52959,G52960,
       G52961,G52962,G52963,G52964,G52965,G52966,G52967,G52968,G52969,G52970,G52971,G52972,G52973,G52974,G52975,G52976,G52977,G52978,G52979,G52980,
       G52981,G52982,G52983,G52984,G52985,G52986,G52987,G52988,G52989,G52990,G52991,G52992,G52993,G52994,G52995,G52996,G52997,G52998,G52999,G53000,
       G53001,G53002,G53003,G53004,G53005,G53006,G53007,G53008,G53009,G53010,G53011,G53012,G53013,G53014,G53015,G53016,G53017,G53018,G53019,G53020,
       G53021,G53022,G53023,G53024,G53025,G53026,G53027,G53028,G53029,G53030,G53031,G53032,G53033,G53034,G53035,G53036,G53037,G53038,G53039,G53040,
       G53041,G53042,G53043,G53044,G53045,G53046,G53047,G53048,G53049,G53050,G53051,G53052,G53053,G53054,G53055,G53056,G53057,G53058,G53059,G53060,
       G53061,G53062,G53063,G53064,G53065,G53066,G53067,G53068,G53069,G53070,G53071,G53072,G53073,G53074,G53075,G53076,G53077,G53078,G53079,G53080,
       G53081,G53082,G53083,G53084,G53085,G53086,G53087,G53088,G53089,G53090,G53091,G53092,G53093,G53094,G53095,G53096,G53097,G53098,G53099,G53100,
       G53101,G53102,G53103,G53104,G53105,G53106,G53107,G53108,G53109,G53110,G53111,G53112,G53113,G53114,G53115,G53116,G53117,G53118,G53119,G53120,
       G53121,G53122,G53123,G53124,G53125,G53126,G53127,G53128,G53129,G53130,G53131,G53132,G53133,G53134,G53135,G53136,G53137,G53138,G53139,G53140,
       G53141,G53142,G53143,G53144,G53145,G53146,G53147,G53148,G53149,G53150,G53151,G53152,G53153,G53154,G53155,G53156,G53157,G53158,G53159,G53160,
       G53161,G53162,G53163,G53164,G53165,G53166,G53167,G53168,G53169,G53170,G53171,G53172,G53173,G53174,G53175,G53176,G53177,G53178,G53179,G53180,
       G53181,G53182,G53183,G53184,G53185,G53186,G53187,G53188,G53189,G53190,G53191,G53192,G53193,G53194,G53195,G53196,G53197,G53198,G53199,G53200,
       G53201,G53202,G53203,G53204,G53205,G53206,G53207,G53208,G53209,G53210,G53211,G53212,G53213,G53214,G53215,G53216,G53217,G53218,G53219,G53220,
       G53221,G53222,G53223,G53224,G53225,G53226,G53227,G53228,G53229,G53230,G53231,G53232,G53233,G53234,G53235,G53236,G53237,G53238,G53239,G53240,
       G53241,G53242,G53243,G53244,G53245,G53246,G53247,G53248,G53249,G53250,G53251,G53252,G53253,G53254,G53255,G53256,G53257,G53258,G53259,G53260,
       G53261,G53262,G53263,G53264,G53265,G53266,G53267,G53268,G53269,G53270,G53271,G53272,G53273,G53274,G53275,G53276,G53277,G53278,G53279,G53280,
       G53281,G53282,G53283,G53284,G53285,G53286,G53287,G53288,G53289,G53290,G53291,G53292,G53293,G53294,G53295,G53296,G53297,G53298,G53299,G53300,
       G53301,G53302,G53303,G53304,G53305,G53306,G53307,G53308,G53309,G53310,G53311,G53312,G53313,G53314,G53315,G53316,G53317,G53318,G53319,G53320,
       G53321,G53322,G53323,G53324,G53325,G53326,G53327,G53328,G53329,G53330,G53331,G53332,G53333,G53334,G53335,G53336,G53337,G53338,G53339,G53340,
       G53341,G53342,G53343,G53344,G53345,G53346,G53347,G53348,G53349,G53350,G53351,G53352,G53353,G53354,G53355,G53356,G53357,G53358,G53359,G53360,
       G53361,G53362,G53363,G53364,G53365,G53366,G53367,G53368,G53369,G53370,G53371,G53372,G53373,G53374,G53375,G53376,G53377,G53378,G53379,G53380,
       G53381,G53382,G53383,G53384,G53385,G53386,G53387,G53388,G53389,G53390,G53391,G53392,G53393,G53394,G53395,G53396,G53397,G53398,G53399,G53400,
       G53401,G53402,G53403,G53404,G53405,G53406,G53407,G53408,G53409,G53410,G53411,G53412,G53413,G53414,G53415,G53416,G53417,G53418,G53419,G53420,
       G53421,G53422,G53423,G53424,G53425,G53426,G53427,G53428,G53429,G53430,G53431,G53432,G53433,G53434,G53435,G53436,G53437,G53438,G53439,G53440,
       G53441,G53442,G53443,G53444,G53445,G53446,G53447,G53448,G53449,G53450,G53451,G53452,G53453,G53454,G53455,G53456,G53457,G53458,G53459,G53460,
       G53461,G53462,G53463,G53464,G53465,G53466,G53467,G53468,G53469,G53470,G53471,G53472,G53473,G53474,G53475,G53476,G53477,G53478,G53479,G53480,
       G53481,G53482,G53483,G53484,G53485,G53486,G53487,G53488,G53489,G53490,G53491,G53492,G53493,G53494,G53495,G53496,G53497,G53498,G53499,G53500,
       G53501,G53502,G53503,G53504,G53505,G53506,G53507,G53508,G53509,G53510,G53511,G53512,G53513,G53514,G53515,G53516,G53517,G53518,G53519,G53520,
       G53521,G53522,G53523,G53524,G53525,G53526,G53527,G53528,G53529,G53530,G53531,G53532,G53533,G53534,G53535,G53536,G53537,G53538,G53539,G53540,
       G53541,G53542,G53543,G53544,G53545,G53546,G53547,G53548,G53549,G53550,G53551,G53552,G53553,G53554,G53555,G53556,G53557,G53558,G53559,G53560,
       G53561,G53562,G53563,G53564,G53565,G53566,G53567,G53568,G53569,G53570,G53571,G53572,G53573,G53574,G53575,G53576,G53577,G53578,G53579,G53580,
       G53581,G53582,G53583,G53584,G53585,G53586,G53587,G53588,G53589,G53590,G53591,G53592,G53593,G53594,G53595,G53596,G53597,G53598,G53599,G53600,
       G53601,G53602,G53603,G53604,G53605,G53606,G53607,G53608,G53609,G53610,G53611,G53612,G53613,G53614,G53615,G53616,G53617,G53618,G53619,G53620,
       G53621,G53622,G53623,G53624,G53625,G53626,G53627,G53628,G53629,G53630,G53631,G53632,G53633,G53634,G53635,G53636,G53637,G53638,G53639,G53640,
       G53641,G53642,G53643,G53644,G53645,G53646,G53647,G53648,G53649,G53650,G53651,G53652,G53653,G53654,G53655,G53656,G53657,G53658,G53659,G53660,
       G53661,G53662,G53663,G53664,G53665,G53666,G53667,G53668,G53669,G53670,G53671,G53672,G53673,G53674,G53675,G53676,G53677,G53678,G53679,G53680,
       G53681,G53682,G53683,G53684,G53685,G53686,G53687,G53688,G53689,G53690,G53691,G53692,G53693,G53694,G53695,G53696,G53697,G53698,G53699,G53700,
       G53701,G53702,G53703,G53704,G53705,G53706,G53707,G53708,G53709,G53710,G53711,G53712,G53713,G53714,G53715,G53716,G53717,G53718,G53719,G53720,
       G53721,G53722,G53723,G53724,G53725,G53726,G53727,G53728,G53729,G53730,G53731,G53732,G53733,G53734,G53735,G53736,G53737,G53738,G53739,G53740,
       G53741,G53742,G53743,G53744,G53745,G53746,G53747,G53748,G53749,G53750,G53751,G53752,G53753,G53754,G53755,G53756,G53757,G53758,G53759,G53760,
       G53761,G53762,G53763,G53764,G53765,G53766,G53767,G53768,G53769,G53770,G53771,G53772,G53773,G53774,G53775,G53776,G53777,G53778,G53779,G53780,
       G53781,G53782,G53783,G53784,G53785,G53786,G53787,G53788,G53789,G53790,G53791,G53792,G53793,G53794,G53795,G53796,G53797,G53798,G53799,G53800,
       G53801,G53802,G53803,G53804,G53805,G53806,G53807,G53808,G53809,G53810,G53811,G53812,G53813,G53814,G53815,G53816,G53817,G53818,G53819,G53820,
       G53821,G53822,G53823,G53824,G53825,G53826,G53827,G53828,G53829,G53830,G53831,G53832,G53833,G53834,G53835,G53836,G53837,G53838,G53839,G53840,
       G53841,G53842,G53843,G53844,G53845,G53846,G53847,G53848,G53849,G53850,G53851,G53852,G53853,G53854,G53855,G53856,G53857,G53858,G53859,G53860,
       G53861,G53862,G53863,G53864,G53865,G53866,G53867,G53868,G53869,G53870,G53871,G53872,G53873,G53874,G53875,G53876,G53877,G53878,G53879,G53880,
       G53881,G53882,G53883,G53884,G53885,G53886,G53887,G53888,G53889,G53890,G53891,G53892,G53893,G53894,G53895,G53896,G53897,G53898,G53899,G53900,
       G53901,G53902,G53903,G53904,G53905,G53906,G53907,G53908,G53909,G53910,G53911,G53912,G53913,G53914,G53915,G53916,G53917,G53918,G53919,G53920,
       G53921,G53922,G53923,G53924,G53925,G53926,G53927,G53928,G53929,G53930,G53931,G53932,G53933,G53934,G53935,G53936,G53937,G53938,G53939,G53940,
       G53941,G53942,G53943,G53944,G53945,G53946,G53947,G53948,G53949,G53950,G53951,G53952,G53953,G53954,G53955,G53956,G53957,G53958,G53959,G53960,
       G53961,G53962,G53963,G53964,G53965,G53966,G53967,G53968,G53969,G53970,G53971,G53972,G53973,G53974,G53975,G53976,G53977,G53978,G53979,G53980,
       G53981,G53982,G53983,G53984,G53985,G53986,G53987,G53988,G53989,G53990,G53991,G53992,G53993,G53994,G53995,G53996,G53997,G53998,G53999,G54000,
       G54001,G54002,G54003,G54004,G54005,G54006,G54007,G54008,G54009,G54010,G54011,G54012,G54013,G54014,G54015,G54016,G54017,G54018,G54019,G54020,
       G54021,G54022,G54023,G54024,G54025,G54026,G54027,G54028,G54029,G54030,G54031,G54032,G54033,G54034,G54035,G54036,G54037,G54038,G54039,G54040,
       G54041,G54042,G54043,G54044,G54045,G54046,G54047,G54048,G54049,G54050,G54051,G54052,G54053,G54054,G54055,G54056,G54057,G54058,G54059,G54060,
       G54061,G54062,G54063,G54064,G54065,G54066,G54067,G54068,G54069,G54070,G54071,G54072,G54073,G54074,G54075,G54076,G54077,G54078,G54079,G54080,
       G54081,G54082,G54083,G54084,G54085,G54086,G54087,G54088,G54089,G54090,G54091,G54092,G54093,G54094,G54095,G54096,G54097,G54098,G54099,G54100,
       G54101,G54102,G54103,G54104,G54105,G54106,G54107,G54108,G54109,G54110,G54111,G54112,G54113,G54114,G54115,G54116,G54117,G54118,G54119,G54120,
       G54121,G54122,G54123,G54124,G54125,G54126,G54127,G54128,G54129,G54130,G54131,G54132,G54133,G54134,G54135,G54136,G54137,G54138,G54139,G54140,
       G54141,G54142,G54143,G54144,G54145,G54146,G54147,G54148,G54149,G54150,G54151,G54152,G54153,G54154,G54155,G54156,G54157,G54158,G54159,G54160,
       G54161,G54162,G54163,G54164,G54165,G54166,G54167,G54168,G54169,G54170,G54171,G54172,G54173,G54174,G54175,G54176,G54177,G54178,G54179,G54180,
       G54181,G54182,G54183,G54184,G54185,G54186,G54187,G54188,G54189,G54190,G54191,G54192,G54193,G54194,G54195,G54196,G54197,G54198,G54199,G54200,
       G54201,G54202,G54203,G54204,G54205,G54206,G54207,G54208,G54209,G54210,G54211,G54212,G54213,G54214,G54215,G54216,G54217,G54218,G54219,G54220,
       G54221,G54222,G54223,G54224,G54225,G54226,G54227,G54228,G54229,G54230,G54231,G54232,G54233,G54234,G54235,G54236,G54237,G54238,G54239,G54240,
       G54241,G54242,G54243,G54244,G54245,G54246,G54247,G54248,G54249,G54250,G54251,G54252,G54253,G54254,G54255,G54256,G54257,G54258,G54259,G54260,
       G54261,G54262,G54263,G54264,G54265,G54266,G54267,G54268,G54269,G54270,G54271,G54272,G54273,G54274,G54275,G54276,G54277,G54278,G54279,G54280,
       G54281,G54282,G54283,G54284,G54285,G54286,G54287,G54288,G54289,G54290,G54291,G54292,G54293,G54294,G54295,G54296,G54297,G54298,G54299,G54300,
       G54301,G54302,G54303,G54304,G54305,G54306,G54307,G54308,G54309,G54310,G54311,G54312,G54313,G54314,G54315,G54316,G54317,G54318,G54319,G54320,
       G54321,G54322,G54323,G54324,G54325,G54326,G54327,G54328,G54329,G54330,G54331,G54332,G54333,G54334,G54335,G54336,G54337,G54338,G54339,G54340,
       G54341,G54342,G54343,G54344,G54345,G54346,G54347,G54348,G54349,G54350,G54351,G54352,G54353,G54354,G54355,G54356,G54357,G54358,G54359,G54360,
       G54361,G54362,G54363,G54364,G54365,G54366,G54367,G54368,G54369,G54370,G54371,G54372,G54373,G54374,G54375,G54376,G54377,G54378,G54379,G54380,
       G54381,G54382,G54383,G54384,G54385,G54386,G54387,G54388,G54389,G54390,G54391,G54392,G54393,G54394,G54395,G54396,G54397,G54398,G54399,G54400,
       G54401,G54402,G54403,G54404,G54405,G54406,G54407,G54408,G54409,G54410,G54411,G54412,G54413,G54414,G54415,G54416,G54417,G54418,G54419,G54420,
       G54421,G54422,G54423,G54424,G54425,G54426,G54427,G54428,G54429,G54430,G54431,G54432,G54433,G54434,G54435,G54436,G54437,G54438,G54439,G54440,
       G54441,G54442,G54443,G54444,G54445,G54446,G54447,G54448,G54449,G54450,G54451,G54452,G54453,G54454,G54455,G54456,G54457,G54458,G54459,G54460,
       G54461,G54462,G54463,G54464,G54465,G54466,G54467,G54468,G54469,G54470,G54471,G54472,G54473,G54474,G54475,G54476,G54477,G54478,G54479,G54480,
       G54481,G54482,G54483,G54484,G54485,G54486,G54487,G54488,G54489,G54490,G54491,G54492,G54493,G54494,G54495,G54496,G54497,G54498,G54499,G54500,
       G54501,G54502,G54503,G54504,G54505,G54506,G54507,G54508,G54509,G54510,G54511,G54512,G54513,G54514,G54515,G54516,G54517,G54518,G54519,G54520,
       G54521,G54522,G54523,G54524,G54525,G54526,G54527,G54528,G54529,G54530,G54531,G54532,G54533,G54534,G54535,G54536,G54537,G54538,G54539,G54540,
       G54541,G54542,G54543,G54544,G54545,G54546,G54547,G54548,G54549,G54550,G54551,G54552,G54553,G54554,G54555,G54556,G54557,G54558,G54559,G54560,
       G54561,G54562,G54563,G54564,G54565,G54566,G54567,G54568,G54569,G54570,G54571,G54572,G54573,G54574,G54575,G54576,G54577,G54578,G54579,G54580,
       G54581,G54582,G54583,G54584,G54585,G54586,G54587,G54588,G54589,G54590,G54591,G54592,G54593,G54594,G54595,G54596,G54597,G54598,G54599,G54600,
       G54601,G54602,G54603,G54604,G54605,G54606,G54607,G54608,G54609,G54610,G54611,G54612,G54613,G54614,G54615,G54616,G54617,G54618,G54619,G54620,
       G54621,G54622,G54623,G54624,G54625,G54626,G54627,G54628,G54629,G54630,G54631,G54632,G54633,G54634,G54635,G54636,G54637,G54638,G54639,G54640,
       G54641,G54642,G54643,G54644,G54645,G54646,G54647,G54648,G54649,G54650,G54651,G54652,G54653,G54654,G54655,G54656,G54657,G54658,G54659,G54660,
       G54661,G54662,G54663,G54664,G54665,G54666,G54667,G54668,G54669,G54670,G54671,G54672,G54673,G54674,G54675,G54676,G54677,G54678,G54679,G54680,
       G54681,G54682,G54683,G54684,G54685,G54686,G54687,G54688,G54689,G54690,G54691,G54692,G54693,G54694,G54695,G54696,G54697,G54698,G54699,G54700,
       G54701,G54702,G54703,G54704,G54705,G54706,G54707,G54708,G54709,G54710,G54711,G54712,G54713,G54714,G54715,G54716,G54717,G54718,G54719,G54720,
       G54721,G54722,G54723,G54724,G54725,G54726,G54727,G54728,G54729,G54730,G54731,G54732,G54733,G54734,G54735,G54736,G54737,G54738,G54739,G54740,
       G54741,G54742,G54743,G54744,G54745,G54746,G54747,G54748,G54749,G54750,G54751,G54752,G54753,G54754,G54755,G54756,G54757,G54758,G54759,G54760,
       G54761,G54762,G54763,G54764,G54765,G54766,G54767,G54768,G54769,G54770,G54771,G54772,G54773,G54774,G54775,G54776,G54777,G54778,G54779,G54780,
       G54781,G54782,G54783,G54784,G54785,G54786,G54787,G54788,G54789,G54790,G54791,G54792,G54793,G54794,G54795,G54796,G54797,G54798,G54799,G54800,
       G54801,G54802,G54803,G54804,G54805,G54806,G54807,G54808,G54809,G54810,G54811,G54812,G54813,G54814,G54815,G54816,G54817,G54818,G54819,G54820,
       G54821,G54822,G54823,G54824,G54825,G54826,G54827,G54828,G54829,G54830,G54831,G54832,G54833,G54834,G54835,G54836,G54837,G54838,G54839,G54840,
       G54841,G54842,G54843,G54844,G54845,G54846,G54847,G54848,G54849,G54850,G54851,G54852,G54853,G54854,G54855,G54856,G54857,G54858,G54859,G54860,
       G54861,G54862,G54863,G54864,G54865,G54866,G54867,G54868,G54869,G54870,G54871,G54872,G54873,G54874,G54875,G54876,G54877,G54878,G54879,G54880,
       G54881,G54882,G54883,G54884,G54885,G54886,G54887,G54888,G54889,G54890,G54891,G54892,G54893,G54894,G54895,G54896,G54897,G54898,G54899,G54900,
       G54901,G54902,G54903,G54904,G54905,G54906,G54907,G54908,G54909,G54910,G54911,G54912,G54913,G54914,G54915,G54916,G54917,G54918,G54919,G54920,
       G54921,G54922,G54923,G54924,G54925,G54926,G54927,G54928,G54929,G54930,G54931,G54932,G54933,G54934,G54935,G54936,G54937,G54938,G54939,G54940,
       G54941,G54942,G54943,G54944,G54945,G54946,G54947,G54948,G54949,G54950,G54951,G54952,G54953,G54954,G54955,G54956,G54957,G54958,G54959,G54960,
       G54961,G54962,G54963,G54964,G54965,G54966,G54967,G54968,G54969,G54970,G54971,G54972,G54973,G54974,G54975,G54976,G54977,G54978,G54979,G54980,
       G54981,G54982,G54983,G54984,G54985,G54986,G54987,G54988,G54989,G54990,G54991,G54992,G54993,G54994,G54995,G54996,G54997,G54998,G54999,G55000,
       G55001,G55002,G55003,G55004,G55005,G55006,G55007,G55008,G55009,G55010,G55011,G55012,G55013,G55014,G55015,G55016,G55017,G55018,G55019,G55020,
       G55021,G55022,G55023,G55024,G55025,G55026,G55027,G55028,G55029,G55030,G55031,G55032,G55033,G55034,G55035,G55036,G55037,G55038,G55039,G55040,
       G55041,G55042,G55043,G55044,G55045,G55046,G55047,G55048,G55049,G55050,G55051,G55052,G55053,G55054,G55055,G55056,G55057,G55058,G55059,G55060,
       G55061,G55062,G55063,G55064,G55065,G55066,G55067,G55068,G55069,G55070,G55071,G55072,G55073,G55074,G55075,G55076,G55077,G55078,G55079,G55080,
       G55081,G55082,G55083,G55084,G55085,G55086,G55087,G55088,G55089,G55090,G55091,G55092,G55093,G55094,G55095,G55096,G55097,G55098,G55099,G55100,
       G55101,G55102,G55103,G55104,G55105,G55106,G55107,G55108,G55109,G55110,G55111,G55112,G55113,G55114,G55115,G55116,G55117,G55118,G55119,G55120,
       G55121,G55122,G55123,G55124,G55125,G55126,G55127,G55128,G55129,G55130,G55131,G55132,G55133,G55134,G55135,G55136,G55137,G55138,G55139,G55140,
       G55141,G55142,G55143,G55144,G55145,G55146,G55147,G55148,G55149,G55150,G55151,G55152,G55153,G55154,G55155,G55156,G55157,G55158,G55159,G55160,
       G55161,G55162,G55163,G55164,G55165,G55166,G55167,G55168,G55169,G55170,G55171,G55172,G55173,G55174,G55175,G55176,G55177,G55178,G55179,G55180,
       G55181,G55182,G55183,G55184,G55185,G55186,G55187,G55188,G55189,G55190,G55191,G55192,G55193,G55194,G55195,G55196,G55197,G55198,G55199,G55200,
       G55201,G55202,G55203,G55204,G55205,G55206,G55207,G55208,G55209,G55210,G55211,G55212,G55213,G55214,G55215,G55216,G55217,G55218,G55219,G55220,
       G55221,G55222,G55223,G55224,G55225,G55226,G55227,G55228,G55229,G55230,G55231,G55232,G55233,G55234,G55235,G55236,G55237,G55238,G55239,G55240,
       G55241,G55242,G55243,G55244,G55245,G55246,G55247,G55248,G55249,G55250,G55251,G55252,G55253,G55254,G55255,G55256,G55257,G55258,G55259,G55260,
       G55261,G55262,G55263,G55264,G55265,G55266,G55267,G55268,G55269,G55270,G55271,G55272,G55273,G55274,G55275,G55276,G55277,G55278,G55279,G55280,
       G55281,G55282,G55283,G55284,G55285,G55286,G55287,G55288,G55289,G55290,G55291,G55292,G55293,G55294,G55295,G55296,G55297,G55298,G55299,G55300,
       G55301,G55302,G55303,G55304,G55305,G55306,G55307,G55308,G55309,G55310,G55311,G55312,G55313,G55314,G55315,G55316,G55317,G55318,G55319,G55320,
       G55321,G55322,G55323,G55324,G55325,G55326,G55327,G55328,G55329,G55330,G55331,G55332,G55333,G55334,G55335,G55336,G55337,G55338,G55339,G55340,
       G55341,G55342,G55343,G55344,G55345,G55346,G55347,G55348,G55349,G55350,G55351,G55352,G55353,G55354,G55355,G55356,G55357,G55358,G55359,G55360,
       G55361,G55362,G55363,G55364,G55365,G55366,G55367,G55368,G55369,G55370,G55371,G55372,G55373,G55374,G55375,G55376,G55377,G55378,G55379,G55380,
       G55381,G55382,G55383,G55384,G55385,G55386,G55387,G55388,G55389,G55390,G55391,G55392,G55393,G55394,G55395,G55396,G55397,G55398,G55399,G55400,
       G55401,G55402,G55403,G55404,G55405,G55406,G55407,G55408,G55409,G55410,G55411,G55412,G55413,G55414,G55415,G55416,G55417,G55418,G55419,G55420,
       G55421,G55422,G55423,G55424,G55425,G55426,G55427,G55428,G55429,G55430,G55431,G55432,G55433,G55434,G55435,G55436,G55437,G55438,G55439,G55440,
       G55441,G55442,G55443,G55444,G55445,G55446,G55447,G55448,G55449,G55450,G55451,G55452,G55453,G55454,G55455,G55456,G55457,G55458,G55459,G55460,
       G55461,G55462,G55463,G55464,G55465,G55466,G55467,G55468,G55469,G55470,G55471,G55472,G55473,G55474,G55475,G55476,G55477,G55478,G55479,G55480,
       G55481,G55482,G55483,G55484,G55485,G55486,G55487,G55488,G55489,G55490,G55491,G55492,G55493,G55494,G55495,G55496,G55497,G55498,G55499,G55500,
       G55501,G55502,G55503,G55504,G55505,G55506,G55507,G55508,G55509,G55510,G55511,G55512,G55513,G55514,G55515,G55516,G55517,G55518,G55519,G55520,
       G55521,G55522,G55523,G55524,G55525,G55526,G55527,G55528,G55529,G55530,G55531,G55532,G55533,G55534,G55535,G55536,G55537,G55538,G55539,G55540,
       G55541,G55542,G55543,G55544,G55545,G55546,G55547,G55548,G55549,G55550,G55551,G55552,G55553,G55554,G55555,G55556,G55557,G55558,G55559,G55560,
       G55561,G55562,G55563,G55564,G55565,G55566,G55567,G55568,G55569,G55570,G55571,G55572,G55573,G55574,G55575,G55576,G55577,G55578,G55579,G55580,
       G55581,G55582,G55583,G55584,G55585,G55586,G55587,G55588,G55589,G55590,G55591,G55592,G55593,G55594,G55595,G55596,G55597,G55598,G55599,G55600,
       G55601,G55602,G55603,G55604,G55605,G55606,G55607,G55608,G55609,G55610,G55611,G55612,G55613,G55614,G55615,G55616,G55617,G55618,G55619,G55620,
       G55621,G55622,G55623,G55624,G55625,G55626,G55627,G55628,G55629,G55630,G55631,G55632,G55633,G55634,G55635,G55636,G55637,G55638,G55639,G55640,
       G55641,G55642,G55643,G55644,G55645,G55646,G55647,G55648,G55649,G55650,G55651,G55652,G55653,G55654,G55655,G55656,G55657,G55658,G55659,G55660,
       G55661,G55662,G55663,G55664,G55665,G55666,G55667,G55668,G55669,G55670,G55671,G55672,G55673,G55674,G55675,G55676,G55677,G55678,G55679,G55680,
       G55681,G55682,G55683,G55684,G55685,G55686,G55687,G55688,G55689,G55690,G55691,G55692,G55693,G55694,G55695,G55696,G55697,G55698,G55699,G55700,
       G55701,G55702,G55703,G55704,G55705,G55706,G55707,G55708,G55709,G55710,G55711,G55712,G55713,G55714,G55715,G55716,G55717,G55718,G55719,G55720,
       G55721,G55722,G55723,G55724,G55725,G55726,G55727,G55728,G55729,G55730,G55731,G55732,G55733,G55734,G55735,G55736,G55737,G55738,G55739,G55740,
       G55741,G55742,G55743,G55744,G55745,G55746,G55747,G55748,G55749,G55750,G55751,G55752,G55753,G55754,G55755,G55756,G55757,G55758,G55759,G55760,
       G55761,G55762,G55763,G55764,G55765,G55766,G55767,G55768,G55769,G55770,G55771,G55772,G55773,G55774,G55775,G55776,G55777,G55778,G55779,G55780,
       G55781,G55782,G55783,G55784,G55785,G55786,G55787,G55788,G55789,G55790,G55791,G55792,G55793,G55794,G55795,G55796,G55797,G55798,G55799,G55800,
       G55801,G55802,G55803,G55804,G55805,G55806,G55807,G55808,G55809,G55810,G55811,G55812,G55813,G55814,G55815,G55816,G55817,G55818,G55819,G55820,
       G55821,G55822,G55823,G55824,G55825,G55826,G55827,G55828,G55829,G55830,G55831,G55832,G55833,G55834,G55835,G55836,G55837,G55838,G55839,G55840,
       G55841,G55842,G55843,G55844,G55845,G55846,G55847,G55848,G55849,G55850,G55851,G55852,G55853,G55854,G55855,G55856,G55857,G55858,G55859,G55860,
       G55861,G55862,G55863,G55864,G55865,G55866,G55867,G55868,G55869,G55870,G55871,G55872,G55873,G55874,G55875,G55876,G55877,G55878,G55879,G55880,
       G55881,G55882,G55883,G55884,G55885,G55886,G55887,G55888,G55889,G55890,G55891,G55892,G55893,G55894,G55895,G55896,G55897,G55898,G55899,G55900,
       G55901,G55902,G55903,G55904,G55905,G55906,G55907,G55908,G55909,G55910,G55911,G55912,G55913,G55914,G55915,G55916,G55917,G55918,G55919,G55920,
       G55921,G55922,G55923,G55924,G55925,G55926,G55927,G55928,G55929,G55930,G55931,G55932,G55933,G55934,G55935,G55936,G55937,G55938,G55939,G55940,
       G55941,G55942,G55943,G55944,G55945,G55946,G55947,G55948,G55949,G55950,G55951,G55952,G55953,G55954,G55955,G55956,G55957,G55958,G55959,G55960,
       G55961,G55962,G55963,G55964,G55965,G55966,G55967,G55968,G55969,G55970,G55971,G55972,G55973,G55974,G55975,G55976,G55977,G55978,G55979,G55980,
       G55981,G55982,G55983,G55984,G55985,G55986,G55987,G55988,G55989,G55990,G55991,G55992,G55993,G55994,G55995,G55996,G55997,G55998,G55999,G56000,
       G56001,G56002,G56003,G56004,G56005,G56006,G56007,G56008,G56009,G56010,G56011,G56012,G56013,G56014,G56015,G56016,G56017,G56018,G56019,G56020,
       G56021,G56022,G56023,G56024,G56025,G56026,G56027,G56028,G56029,G56030,G56031,G56032,G56033,G56034,G56035,G56036,G56037,G56038,G56039,G56040,
       G56041,G56042,G56043,G56044,G56045,G56046,G56047,G56048,G56049,G56050,G56051,G56052,G56053,G56054,G56055,G56056,G56057,G56058,G56059,G56060,
       G56061,G56062,G56063,G56064,G56065,G56066,G56067,G56068,G56069,G56070,G56071,G56072,G56073,G56074,G56075,G56076,G56077,G56078,G56079,G56080,
       G56081,G56082,G56083,G56084,G56085,G56086,G56087,G56088,G56089,G56090,G56091,G56092,G56093,G56094,G56095,G56096,G56097,G56098,G56099,G56100,
       G56101,G56102,G56103,G56104,G56105,G56106,G56107,G56108,G56109,G56110,G56111,G56112,G56113,G56114,G56115,G56116,G56117,G56118,G56119,G56120,
       G56121,G56122,G56123,G56124,G56125,G56126,G56127,G56128,G56129,G56130,G56131,G56132,G56133,G56134,G56135,G56136,G56137,G56138,G56139,G56140,
       G56141,G56142,G56143,G56144,G56145,G56146,G56147,G56148,G56149,G56150,G56151,G56152,G56153,G56154,G56155,G56156,G56157,G56158,G56159,G56160,
       G56161,G56162,G56163,G56164,G56165,G56166,G56167,G56168,G56169,G56170,G56171,G56172,G56173,G56174,G56175,G56176,G56177,G56178,G56179,G56180,
       G56181,G56182,G56183,G56184,G56185,G56186,G56187,G56188,G56189,G56190,G56191,G56192,G56193,G56194,G56195,G56196,G56197,G56198,G56199,G56200,
       G56201,G56202,G56203,G56204,G56205,G56206,G56207,G56208,G56209,G56210,G56211,G56212,G56213,G56214,G56215,G56216,G56217,G56218,G56219,G56220,
       G56221,G56222,G56223,G56224,G56225,G56226,G56227,G56228,G56229,G56230,G56231,G56232,G56233,G56234,G56235,G56236,G56237,G56238,G56239,G56240,
       G56241,G56242,G56243,G56244,G56245,G56246,G56247,G56248,G56249,G56250,G56251,G56252,G56253,G56254,G56255,G56256,G56257,G56258,G56259,G56260,
       G56261,G56262,G56263,G56264,G56265,G56266,G56267,G56268,G56269,G56270,G56271,G56272,G56273,G56274,G56275,G56276,G56277,G56278,G56279,G56280,
       G56281,G56282,G56283,G56284,G56285,G56286,G56287,G56288,G56289,G56290,G56291,G56292,G56293,G56294,G56295,G56296,G56297,G56298,G56299,G56300,
       G56301,G56302,G56303,G56304,G56305,G56306,G56307,G56308,G56309,G56310,G56311,G56312,G56313,G56314,G56315,G56316,G56317,G56318,G56319,G56320,
       G56321,G56322,G56323,G56324,G56325,G56326,G56327,G56328,G56329,G56330,G56331,G56332,G56333,G56334,G56335,G56336,G56337,G56338,G56339,G56340,
       G56341,G56342,G56343,G56344,G56345,G56346,G56347,G56348,G56349,G56350,G56351,G56352,G56353,G56354,G56355,G56356,G56357,G56358,G56359,G56360,
       G56361,G56362,G56363,G56364,G56365,G56366,G56367,G56368,G56369,G56370,G56371,G56372,G56373,G56374,G56375,G56376,G56377,G56378,G56379,G56380,
       G56381,G56382,G56383,G56384,G56385,G56386,G56387,G56388,G56389,G56390,G56391,G56392,G56393,G56394,G56395,G56396,G56397,G56398,G56399,G56400,
       G56401,G56402,G56403,G56404,G56405,G56406,G56407,G56408,G56409,G56410,G56411,G56412,G56413,G56414,G56415,G56416,G56417,G56418,G56419,G56420,
       G56421,G56422,G56423,G56424,G56425,G56426,G56427,G56428,G56429,G56430,G56431,G56432,G56433,G56434,G56435,G56436,G56437,G56438,G56439,G56440,
       G56441,G56442,G56443,G56444,G56445,G56446,G56447,G56448,G56449,G56450,G56451,G56452,G56453,G56454,G56455,G56456,G56457,G56458,G56459,G56460,
       G56461,G56462,G56463,G56464,G56465,G56466,G56467,G56468,G56469,G56470,G56471,G56472,G56473,G56474,G56475,G56476,G56477,G56478,G56479,G56480,
       G56481,G56482,G56483,G56484,G56485,G56486,G56487,G56488,G56489,G56490,G56491,G56492,G56493,G56494,G56495,G56496,G56497,G56498,G56499,G56500,
       G56501,G56502,G56503,G56504,G56505,G56506,G56507,G56508,G56509,G56510,G56511,G56512,G56513,G56514,G56515,G56516,G56517,G56518,G56519,G56520,
       G56521,G56522,G56523,G56524,G56525,G56526,G56527,G56528,G56529,G56530,G56531,G56532,G56533,G56534,G56535,G56536,G56537,G56538,G56539,G56540,
       G56541,G56542,G56543,G56544,G56545,G56546,G56547,G56548,G56549,G56550,G56551,G56552,G56553,G56554,G56555,G56556,G56557,G56558,G56559,G56560,
       G56561,G56562,G56563,G56564,G56565,G56566,G56567,G56568,G56569,G56570,G56571,G56572,G56573,G56574,G56575,G56576,G56577,G56578,G56579,G56580,
       G56581,G56582,G56583,G56584,G56585,G56586,G56587,G56588,G56589,G56590,G56591,G56592,G56593,G56594,G56595,G56596,G56597,G56598,G56599,G56600,
       G56601,G56602,G56603,G56604,G56605,G56606,G56607,G56608,G56609,G56610,G56611,G56612,G56613,G56614,G56615,G56616,G56617,G56618,G56619,G56620,
       G56621,G56622,G56623,G56624,G56625,G56626,G56627,G56628,G56629,G56630,G56631,G56632,G56633,G56634,G56635,G56636,G56637,G56638,G56639,G56640,
       G56641,G56642,G56643,G56644,G56645,G56646,G56647,G56648,G56649,G56650,G56651,G56652,G56653,G56654,G56655,G56656,G56657,G56658,G56659,G56660,
       G56661,G56662,G56663,G56664,G56665,G56666,G56667,G56668,G56669,G56670,G56671,G56672,G56673,G56674,G56675,G56676,G56677,G56678,G56679,G56680,
       G56681,G56682,G56683,G56684,G56685,G56686,G56687,G56688,G56689,G56690,G56691,G56692,G56693,G56694,G56695,G56696,G56697,G56698,G56699,G56700,
       G56701,G56702,G56703,G56704,G56705,G56706,G56707,G56708,G56709,G56710,G56711,G56712,G56713,G56714,G56715,G56716,G56717,G56718,G56719,G56720,
       G56721,G56722,G56723,G56724,G56725,G56726,G56727,G56728,G56729,G56730,G56731,G56732,G56733,G56734,G56735,G56736,G56737,G56738,G56739,G56740,
       G56741,G56742,G56743,G56744,G56745,G56746,G56747,G56748,G56749,G56750,G56751,G56752,G56753,G56754,G56755,G56756,G56757,G56758,G56759,G56760,
       G56761,G56762,G56763,G56764,G56765,G56766,G56767,G56768,G56769,G56770,G56771,G56772,G56773,G56774,G56775,G56776,G56777,G56778,G56779,G56780,
       G56781,G56782,G56783,G56784,G56785,G56786,G56787,G56788,G56789,G56790,G56791,G56792,G56793,G56794,G56795,G56796,G56797,G56798,G56799,G56800,
       G56801,G56802,G56803,G56804,G56805,G56806,G56807,G56808,G56809,G56810,G56811,G56812,G56813,G56814,G56815,G56816,G56817,G56818,G56819,G56820,
       G56821,G56822,G56823,G56824,G56825,G56826,G56827,G56828,G56829,G56830,G56831,G56832,G56833,G56834,G56835,G56836,G56837,G56838,G56839,G56840,
       G56841,G56842,G56843,G56844,G56845,G56846,G56847,G56848,G56849,G56850,G56851,G56852,G56853,G56854,G56855,G56856,G56857,G56858,G56859,G56860,
       G56861,G56862,G56863,G56864,G56865,G56866,G56867,G56868,G56869,G56870,G56871,G56872,G56873,G56874,G56875,G56876,G56877,G56878,G56879,G56880,
       G56881,G56882,G56883,G56884,G56885,G56886,G56887,G56888,G56889,G56890,G56891,G56892,G56893,G56894,G56895,G56896,G56897,G56898,G56899,G56900,
       G56901,G56902,G56903,G56904,G56905,G56906,G56907,G56908,G56909,G56910,G56911,G56912,G56913,G56914,G56915,G56916,G56917,G56918,G56919,G56920,
       G56921,G56922,G56923,G56924,G56925,G56926,G56927,G56928,G56929,G56930,G56931,G56932,G56933,G56934,G56935,G56936,G56937,G56938,G56939,G56940,
       G56941,G56942,G56943,G56944,G56945,G56946,G56947,G56948,G56949,G56950,G56951,G56952,G56953,G56954,G56955,G56956,G56957,G56958,G56959,G56960,
       G56961,G56962,G56963,G56964,G56965,G56966,G56967,G56968,G56969,G56970,G56971,G56972,G56973,G56974,G56975,G56976,G56977,G56978,G56979,G56980,
       G56981,G56982,G56983,G56984,G56985,G56986,G56987,G56988,G56989,G56990,G56991,G56992,G56993,G56994,G56995,G56996,G56997,G56998,G56999,G57000,
       G57001,G57002,G57003,G57004,G57005,G57006,G57007,G57008,G57009,G57010,G57011,G57012,G57013,G57014,G57015,G57016,G57017,G57018,G57019,G57020,
       G57021,G57022,G57023,G57024,G57025,G57026,G57027,G57028,G57029,G57030,G57031,G57032,G57033,G57034,G57035,G57036,G57037,G57038,G57039,G57040,
       G57041,G57042,G57043,G57044,G57045,G57046,G57047,G57048,G57049,G57050,G57051,G57052,G57053,G57054,G57055,G57056,G57057,G57058,G57059,G57060,
       G57061,G57062,G57063,G57064,G57065,G57066,G57067,G57068,G57069,G57070,G57071,G57072,G57073,G57074,G57075,G57076,G57077,G57078,G57079,G57080,
       G57081,G57082,G57083,G57084,G57085,G57086,G57087,G57088,G57089,G57090,G57091,G57092,G57093,G57094,G57095,G57096,G57097,G57098,G57099,G57100,
       G57101,G57102,G57103,G57104,G57105,G57106,G57107,G57108,G57109,G57110,G57111,G57112,G57113,G57114,G57115,G57116,G57117,G57118,G57119,G57120,
       G57121,G57122,G57123,G57124,G57125,G57126,G57127,G57128,G57129,G57130,G57131,G57132,G57133,G57134,G57135,G57136,G57137,G57138,G57139,G57140,
       G57141,G57142,G57143,G57144,G57145,G57146,G57147,G57148,G57149,G57150,G57151,G57152,G57153,G57154,G57155,G57156,G57157,G57158,G57159,G57160,
       G57161,G57162,G57163,G57164,G57165,G57166,G57167,G57168,G57169,G57170,G57171,G57172,G57173,G57174,G57175,G57176,G57177,G57178,G57179,G57180,
       G57181,G57182,G57183,G57184,G57185,G57186,G57187,G57188,G57189,G57190,G57191,G57192,G57193,G57194,G57195,G57196,G57197,G57198,G57199,G57200,
       G57201,G57202,G57203,G57204,G57205,G57206,G57207,G57208,G57209,G57210,G57211,G57212,G57213,G57214,G57215,G57216,G57217,G57218,G57219,G57220,
       G57221,G57222,G57223,G57224,G57225,G57226,G57227,G57228,G57229,G57230,G57231,G57232,G57233,G57234,G57235,G57236,G57237,G57238,G57239,G57240,
       G57241,G57242,G57243,G57244,G57245,G57246,G57247,G57248,G57249,G57250,G57251,G57252,G57253,G57254,G57255,G57256,G57257,G57258,G57259,G57260,
       G57261,G57262,G57263,G57264,G57265,G57266,G57267,G57268,G57269,G57270,G57271,G57272,G57273,G57274,G57275,G57276,G57277,G57278,G57279,G57280,
       G57281,G57282,G57283,G57284,G57285,G57286,G57287,G57288,G57289,G57290,G57291,G57292,G57293,G57294,G57295,G57296,G57297,G57298,G57299,G57300,
       G57301,G57302,G57303,G57304,G57305,G57306,G57307,G57308,G57309,G57310,G57311,G57312,G57313,G57314,G57315,G57316,G57317,G57318,G57319,G57320,
       G57321,G57322,G57323,G57324,G57325,G57326,G57327,G57328,G57329,G57330,G57331,G57332,G57333,G57334,G57335,G57336,G57337,G57338,G57339,G57340,
       G57341,G57342,G57343,G57344,G57345,G57346,G57347,G57348,G57349,G57350,G57351,G57352,G57353,G57354,G57355,G57356,G57357,G57358,G57359,G57360,
       G57361,G57362,G57363,G57364,G57365,G57366,G57367,G57368,G57369,G57370,G57371,G57372,G57373,G57374,G57375,G57376,G57377,G57378,G57379,G57380,
       G57381,G57382,G57383,G57384,G57385,G57386,G57387,G57388,G57389,G57390,G57391,G57392,G57393,G57394,G57395,G57396,G57397,G57398,G57399,G57400,
       G57401,G57402,G57403,G57404,G57405,G57406,G57407,G57408,G57409,G57410,G57411,G57412,G57413,G57414,G57415,G57416,G57417,G57418,G57419,G57420,
       G57421,G57422,G57423,G57424,G57425,G57426,G57427,G57428,G57429,G57430,G57431,G57432,G57433,G57434,G57435,G57436,G57437,G57438,G57439,G57440,
       G57441,G57442,G57443,G57444,G57445,G57446,G57447,G57448,G57449,G57450,G57451,G57452,G57453,G57454,G57455,G57456,G57457,G57458,G57459,G57460,
       G57461,G57462,G57463,G57464,G57465,G57466,G57467,G57468,G57469,G57470,G57471,G57472,G57473,G57474,G57475,G57476,G57477,G57478,G57479,G57480,
       G57481,G57482,G57483,G57484,G57485,G57486,G57487,G57488,G57489,G57490,G57491,G57492,G57493,G57494,G57495,G57496,G57497,G57498,G57499,G57500,
       G57501,G57502,G57503,G57504,G57505,G57506,G57507,G57508,G57509,G57510,G57511,G57512,G57513,G57514,G57515,G57516,G57517,G57518,G57519,G57520,
       G57521,G57522,G57523,G57524,G57525,G57526,G57527,G57528,G57529,G57530,G57531,G57532,G57533,G57534,G57535,G57536,G57537,G57538,G57539,G57540,
       G57541,G57542,G57543,G57544,G57545,G57546,G57547,G57548,G57549,G57550,G57551,G57552,G57553,G57554,G57555,G57556,G57557,G57558,G57559,G57560,
       G57561,G57562,G57563,G57564,G57565,G57566,G57567,G57568,G57569,G57570,G57571,G57572,G57573,G57574,G57575,G57576,G57577,G57578,G57579,G57580,
       G57581,G57582,G57583,G57584,G57585,G57586,G57587,G57588,G57589,G57590,G57591,G57592,G57593,G57594,G57595,G57596,G57597,G57598,G57599,G57600,
       G57601,G57602,G57603,G57604,G57605,G57606,G57607,G57608,G57609,G57610,G57611,G57612,G57613,G57614,G57615,G57616,G57617,G57618,G57619,G57620,
       G57621,G57622,G57623,G57624,G57625,G57626,G57627,G57628,G57629,G57630,G57631,G57632,G57633,G57634,G57635,G57636,G57637,G57638,G57639,G57640,
       G57641,G57642,G57643,G57644,G57645,G57646,G57647,G57648,G57649,G57650,G57651,G57652,G57653,G57654,G57655,G57656,G57657,G57658,G57659,G57660,
       G57661,G57662,G57663,G57664,G57665,G57666,G57667,G57668,G57669,G57670,G57671,G57672,G57673,G57674,G57675,G57676,G57677,G57678,G57679,G57680,
       G57681,G57682,G57683,G57684,G57685,G57686,G57687,G57688,G57689,G57690,G57691,G57692,G57693,G57694,G57695,G57696,G57697,G57698,G57699,G57700,
       G57701,G57702,G57703,G57704,G57705,G57706,G57707,G57708,G57709,G57710,G57711,G57712,G57713,G57714,G57715,G57716,G57717,G57718,G57719,G57720,
       G57721,G57722,G57723,G57724,G57725,G57726,G57727,G57728,G57729,G57730,G57731,G57732,G57733,G57734,G57735,G57736,G57737,G57738,G57739,G57740,
       G57741,G57742,G57743,G57744,G57745,G57746,G57747,G57748,G57749,G57750,G57751,G57752,G57753,G57754,G57755,G57756,G57757,G57758,G57759,G57760,
       G57761,G57762,G57763,G57764,G57765,G57766,G57767,G57768,G57769,G57770,G57771,G57772,G57773,G57774,G57775,G57776,G57777,G57778,G57779,G57780,
       G57781,G57782,G57783,G57784,G57785,G57786,G57787,G57788,G57789,G57790,G57791,G57792,G57793,G57794,G57795,G57796,G57797,G57798,G57799,G57800,
       G57801,G57802,G57803,G57804,G57805,G57806,G57807,G57808,G57809,G57810,G57811,G57812,G57813,G57814,G57815,G57816,G57817,G57818,G57819,G57820,
       G57821,G57822,G57823,G57824,G57825,G57826,G57827,G57828,G57829,G57830,G57831,G57832,G57833,G57834,G57835,G57836,G57837,G57838,G57839,G57840,
       G57841,G57842,G57843,G57844,G57845,G57846,G57847,G57848,G57849,G57850,G57851,G57852,G57853,G57854,G57855,G57856,G57857,G57858,G57859,G57860,
       G57861,G57862,G57863,G57864,G57865,G57866,G57867,G57868,G57869,G57870,G57871,G57872,G57873,G57874,G57875,G57876,G57877,G57878,G57879,G57880,
       G57881,G57882,G57883,G57884,G57885,G57886,G57887,G57888,G57889,G57890,G57891,G57892,G57893,G57894,G57895,G57896,G57897,G57898,G57899,G57900,
       G57901,G57902,G57903,G57904,G57905,G57906,G57907,G57908,G57909,G57910,G57911,G57912,G57913,G57914,G57915,G57916,G57917,G57918,G57919,G57920,
       G57921,G57922,G57923,G57924,G57925,G57926,G57927,G57928,G57929,G57930,G57931,G57932,G57933,G57934,G57935,G57936,G57937,G57938,G57939,G57940,
       G57941,G57942,G57943,G57944,G57945,G57946,G57947,G57948,G57949,G57950,G57951,G57952,G57953,G57954,G57955,G57956,G57957,G57958,G57959,G57960,
       G57961,G57962,G57963,G57964,G57965,G57966,G57967,G57968,G57969,G57970,G57971,G57972,G57973,G57974,G57975,G57976,G57977,G57978,G57979,G57980,
       G57981,G57982,G57983,G57984,G57985,G57986,G57987,G57988,G57989,G57990,G57991,G57992,G57993,G57994,G57995,G57996,G57997,G57998,G57999,G58000,
       G58001,G58002,G58003,G58004,G58005,G58006,G58007,G58008,G58009,G58010,G58011,G58012,G58013,G58014,G58015,G58016,G58017,G58018,G58019,G58020,
       G58021,G58022,G58023,G58024,G58025,G58026,G58027,G58028,G58029,G58030,G58031,G58032,G58033,G58034,G58035,G58036,G58037,G58038,G58039,G58040,
       G58041,G58042,G58043,G58044,G58045,G58046,G58047,G58048,G58049,G58050,G58051,G58052,G58053,G58054,G58055,G58056,G58057,G58058,G58059,G58060,
       G58061,G58062,G58063,G58064,G58065,G58066,G58067,G58068,G58069,G58070,G58071,G58072,G58073,G58074,G58075,G58076,G58077,G58078,G58079,G58080,
       G58081,G58082,G58083,G58084,G58085,G58086,G58087,G58088,G58089,G58090,G58091,G58092,G58093,G58094,G58095,G58096,G58097,G58098,G58099,G58100,
       G58101,G58102,G58103,G58104,G58105,G58106,G58107,G58108,G58109,G58110,G58111,G58112,G58113,G58114,G58115,G58116,G58117,G58118,G58119,G58120,
       G58121,G58122,G58123,G58124,G58125,G58126,G58127,G58128,G58129,G58130,G58131,G58132,G58133,G58134,G58135,G58136,G58137,G58138,G58139,G58140,
       G58141,G58142,G58143,G58144,G58145,G58146,G58147,G58148,G58149,G58150,G58151,G58152,G58153,G58154,G58155,G58156,G58157,G58158,G58159,G58160,
       G58161,G58162,G58163,G58164,G58165,G58166,G58167,G58168,G58169,G58170,G58171,G58172,G58173,G58174,G58175,G58176,G58177,G58178,G58179,G58180,
       G58181,G58182,G58183,G58184,G58185,G58186,G58187,G58188,G58189,G58190,G58191,G58192,G58193,G58194,G58195,G58196,G58197,G58198,G58199,G58200,
       G58201,G58202,G58203,G58204,G58205,G58206,G58207,G58208,G58209,G58210,G58211,G58212,G58213,G58214,G58215,G58216,G58217,G58218,G58219,G58220,
       G58221,G58222,G58223,G58224,G58225,G58226,G58227,G58228,G58229,G58230,G58231,G58232,G58233,G58234,G58235,G58236,G58237,G58238,G58239,G58240,
       G58241,G58242,G58243,G58244,G58245,G58246,G58247,G58248,G58249,G58250,G58251,G58252,G58253,G58254,G58255,G58256,G58257,G58258,G58259,G58260,
       G58261,G58262,G58263,G58264,G58265,G58266,G58267,G58268,G58269,G58270,G58271,G58272,G58273,G58274,G58275,G58276,G58277,G58278,G58279,G58280,
       G58281,G58282,G58283,G58284,G58285,G58286,G58287,G58288,G58289,G58290,G58291,G58292,G58293,G58294,G58295,G58296,G58297,G58298,G58299,G58300,
       G58301,G58302,G58303,G58304,G58305,G58306,G58307,G58308,G58309,G58310,G58311,G58312,G58313,G58314,G58315,G58316,G58317,G58318,G58319,G58320,
       G58321,G58322,G58323,G58324,G58325,G58326,G58327,G58328,G58329,G58330,G58331,G58332,G58333,G58334,G58335,G58336,G58337,G58338,G58339,G58340,
       G58341,G58342,G58343,G58344,G58345,G58346,G58347,G58348,G58349,G58350,G58351,G58352,G58353,G58354,G58355,G58356,G58357,G58358,G58359,G58360,
       G58361,G58362,G58363,G58364,G58365,G58366,G58367,G58368,G58369,G58370,G58371,G58372,G58373,G58374,G58375,G58376,G58377,G58378,G58379,G58380,
       G58381,G58382,G58383,G58384,G58385,G58386,G58387,G58388,G58389,G58390,G58391,G58392,G58393,G58394,G58395,G58396,G58397,G58398,G58399,G58400,
       G58401,G58402,G58403,G58404,G58405,G58406,G58407,G58408,G58409,G58410,G58411,G58412,G58413,G58414,G58415,G58416,G58417,G58418,G58419,G58420,
       G58421,G58422,G58423,G58424,G58425,G58426,G58427,G58428,G58429,G58430,G58431,G58432,G58433,G58434,G58435,G58436,G58437,G58438,G58439,G58440,
       G58441,G58442,G58443,G58444,G58445,G58446,G58447,G58448,G58449,G58450,G58451,G58452,G58453,G58454,G58455,G58456,G58457,G58458,G58459,G58460,
       G58461,G58462,G58463,G58464,G58465,G58466,G58467,G58468,G58469,G58470,G58471,G58472,G58473,G58474,G58475,G58476,G58477,G58478,G58479,G58480,
       G58481,G58482,G58483,G58484,G58485,G58486,G58487,G58488,G58489,G58490,G58491,G58492,G58493,G58494,G58495,G58496,G58497,G58498,G58499,G58500,
       G58501,G58502,G58503,G58504,G58505,G58506,G58507,G58508,G58509,G58510,G58511,G58512,G58513,G58514,G58515,G58516,G58517,G58518,G58519,G58520,
       G58521,G58522,G58523,G58524,G58525,G58526,G58527,G58528,G58529,G58530,G58531,G58532,G58533,G58534,G58535,G58536,G58537,G58538,G58539,G58540,
       G58541,G58542,G58543,G58544,G58545,G58546,G58547,G58548,G58549,G58550,G58551,G58552,G58553,G58554,G58555,G58556,G58557,G58558,G58559,G58560,
       G58561,G58562,G58563,G58564,G58565,G58566,G58567,G58568,G58569,G58570,G58571,G58572,G58573,G58574,G58575,G58576,G58577,G58578,G58579,G58580,
       G58581,G58582,G58583,G58584,G58585,G58586,G58587,G58588,G58589,G58590,G58591,G58592,G58593,G58594,G58595,G58596,G58597,G58598,G58599,G58600,
       G58601,G58602,G58603,G58604,G58605,G58606,G58607,G58608,G58609,G58610,G58611,G58612,G58613,G58614,G58615,G58616,G58617,G58618,G58619,G58620,
       G58621,G58622,G58623,G58624,G58625,G58626,G58627,G58628,G58629,G58630,G58631,G58632,G58633,G58634,G58635,G58636,G58637,G58638,G58639,G58640,
       G58641,G58642,G58643,G58644,G58645,G58646,G58647,G58648,G58649,G58650,G58651,G58652,G58653,G58654,G58655,G58656,G58657,G58658,G58659,G58660,
       G58661,G58662,G58663,G58664,G58665,G58666,G58667,G58668,G58669,G58670,G58671,G58672,G58673,G58674,G58675,G58676,G58677,G58678,G58679,G58680,
       G58681,G58682,G58683,G58684,G58685,G58686,G58687,G58688,G58689,G58690,G58691,G58692,G58693,G58694,G58695,G58696,G58697,G58698,G58699,G58700,
       G58701,G58702,G58703,G58704,G58705,G58706,G58707,G58708,G58709,G58710,G58711,G58712,G58713,G58714,G58715,G58716,G58717,G58718,G58719,G58720,
       G58721,G58722,G58723,G58724,G58725,G58726,G58727,G58728,G58729,G58730,G58731,G58732,G58733,G58734,G58735,G58736,G58737,G58738,G58739,G58740,
       G58741,G58742,G58743,G58744,G58745,G58746,G58747,G58748,G58749,G58750,G58751,G58752,G58753,G58754,G58755,G58756,G58757,G58758,G58759,G58760,
       G58761,G58762,G58763,G58764,G58765,G58766,G58767,G58768,G58769,G58770,G58771,G58772,G58773,G58774,G58775,G58776,G58777,G58778,G58779,G58780,
       G58781,G58782,G58783,G58784,G58785,G58786,G58787,G58788,G58789,G58790,G58791,G58792,G58793,G58794,G58795,G58796,G58797,G58798,G58799,G58800,
       G58801,G58802,G58803,G58804,G58805,G58806,G58807,G58808,G58809,G58810,G58811,G58812,G58813,G58814,G58815,G58816,G58817,G58818,G58819,G58820,
       G58821,G58822,G58823,G58824,G58825,G58826,G58827,G58828,G58829,G58830,G58831,G58832,G58833,G58834,G58835,G58836,G58837,G58838,G58839,G58840,
       G58841,G58842,G58843,G58844,G58845,G58846,G58847,G58848,G58849,G58850,G58851,G58852,G58853,G58854,G58855,G58856,G58857,G58858,G58859,G58860,
       G58861,G58862,G58863,G58864,G58865,G58866,G58867,G58868,G58869,G58870,G58871,G58872,G58873,G58874,G58875,G58876,G58877,G58878,G58879,G58880,
       G58881,G58882,G58883,G58884,G58885,G58886,G58887,G58888,G58889,G58890,G58891,G58892,G58893,G58894,G58895,G58896,G58897,G58898,G58899,G58900,
       G58901,G58902,G58903,G58904,G58905,G58906,G58907,G58908,G58909,G58910,G58911,G58912,G58913,G58914,G58915,G58916,G58917,G58918,G58919,G58920,
       G58921,G58922,G58923,G58924,G58925,G58926,G58927,G58928,G58929,G58930,G58931,G58932,G58933,G58934,G58935,G58936,G58937,G58938,G58939,G58940,
       G58941,G58942,G58943,G58944,G58945,G58946,G58947,G58948,G58949,G58950,G58951,G58952,G58953,G58954,G58955,G58956,G58957,G58958,G58959,G58960,
       G58961,G58962,G58963,G58964,G58965,G58966,G58967,G58968,G58969,G58970,G58971,G58972,G58973,G58974,G58975,G58976,G58977,G58978,G58979,G58980,
       G58981,G58982,G58983,G58984,G58985,G58986,G58987,G58988,G58989,G58990,G58991,G58992,G58993,G58994,G58995,G58996,G58997,G58998,G58999,G59000,
       G59001,G59002,G59003,G59004,G59005,G59006,G59007,G59008,G59009,G59010,G59011,G59012,G59013,G59014,G59015,G59016,G59017,G59018,G59019,G59020,
       G59021,G59022,G59023,G59024,G59025,G59026,G59027,G59028,G59029,G59030,G59031,G59032,G59033,G59034,G59035,G59036,G59037,G59038,G59039,G59040,
       G59041,G59042,G59043,G59044,G59045,G59046,G59047,G59048,G59049,G59050,G59051,G59052,G59053,G59054,G59055,G59056,G59057,G59058,G59059,G59060,
       G59061,G59062,G59063,G59064,G59065,G59066,G59067,G59068,G59069,G59070,G59071,G59072,G59073,G59074,G59075,G59076,G59077,G59078,G59079,G59080,
       G59081,G59082,G59083,G59084,G59085,G59086,G59087,G59088,G59089,G59090,G59091,G59092,G59093,G59094,G59095,G59096,G59097,G59098,G59099,G59100,
       G59101,G59102,G59103,G59104,G59105,G59106,G59107,G59108,G59109,G59110,G59111,G59112,G59113,G59114,G59115,G59116,G59117,G59118,G59119,G59120,
       G59121,G59122,G59123,G59124,G59125,G59126,G59127,G59128,G59129,G59130,G59131,G59132,G59133,G59134,G59135,G59136,G59137,G59138,G59139,G59140,
       G59141,G59142,G59143,G59144,G59145,G59146,G59147,G59148,G59149,G59150,G59151,G59152,G59153,G59154,G59155,G59156,G59157,G59158,G59159,G59160,
       G59161,G59162,G59163,G59164,G59165,G59166,G59167,G59168,G59169,G59170,G59171,G59172,G59173,G59174,G59175,G59176,G59177,G59178,G59179,G59180,
       G59181,G59182,G59183,G59184,G59185,G59186,G59187,G59188,G59189,G59190,G59191,G59192,G59193,G59194,G59195,G59196,G59197,G59198,G59199,G59200,
       G59201,G59202,G59203,G59204,G59205,G59206,G59207,G59208,G59209,G59210,G59211,G59212,G59213,G59214,G59215,G59216,G59217,G59218,G59219,G59220,
       G59221,G59222,G59223,G59224,G59225,G59226,G59227,G59228,G59229,G59230,G59231,G59232,G59233,G59234,G59235,G59236,G59237,G59238,G59239,G59240,
       G59241,G59242,G59243,G59244,G59245,G59246,G59247,G59248,G59249,G59250,G59251,G59252,G59253,G59254,G59255,G59256,G59257,G59258,G59259,G59260,
       G59261,G59262,G59263,G59264,G59265,G59266,G59267,G59268,G59269,G59270,G59271,G59272,G59273,G59274,G59275,G59276,G59277,G59278,G59279,G59280,
       G59281,G59282,G59283,G59284,G59285,G59286,G59287,G59288,G59289,G59290,G59291,G59292,G59293,G59294,G59295,G59296,G59297,G59298,G59299,G59300,
       G59301,G59302,G59303,G59304,G59305,G59306,G59307,G59308,G59309,G59310,G59311,G59312,G59313,G59314,G59315,G59316,G59317,G59318,G59319,G59320,
       G59321,G59322,G59323,G59324,G59325,G59326,G59327,G59328,G59329,G59330,G59331,G59332,G59333,G59334,G59335,G59336,G59337,G59338,G59339,G59340,
       G59341,G59342,G59343,G59344,G59345,G59346,G59347,G59348,G59349,G59350,G59351,G59352,G59353,G59354,G59355,G59356,G59357,G59358,G59359,G59360,
       G59361,G59362,G59363,G59364,G59365,G59366,G59367,G59368,G59369,G59370,G59371,G59372,G59373,G59374,G59375,G59376,G59377,G59378,G59379,G59380,
       G59381,G59382,G59383,G59384,G59385,G59386,G59387,G59388,G59389,G59390,G59391,G59392,G59393,G59394,G59395,G59396,G59397,G59398,G59399,G59400,
       G59401,G59402,G59403,G59404,G59405,G59406,G59407,G59408,G59409,G59410,G59411,G59412,G59413,G59414,G59415,G59416,G59417,G59418,G59419,G59420,
       G59421,G59422,G59423,G59424,G59425,G59426,G59427,G59428,G59429,G59430,G59431,G59432,G59433,G59434,G59435,G59436,G59437,G59438,G59439,G59440,
       G59441,G59442,G59443,G59444,G59445,G59446,G59447,G59448,G59449,G59450,G59451,G59452,G59453,G59454,G59455,G59456,G59457,G59458,G59459,G59460,
       G59461,G59462,G59463,G59464,G59465,G59466,G59467,G59468,G59469,G59470,G59471,G59472,G59473,G59474,G59475,G59476,G59477,G59478,G59479,G59480,
       G59481,G59482,G59483,G59484,G59485,G59486,G59487,G59488,G59489,G59490,G59491,G59492,G59493,G59494,G59495,G59496,G59497,G59498,G59499,G59500,
       G59501,G59502,G59503,G59504,G59505,G59506,G59507,G59508,G59509,G59510,G59511,G59512,G59513,G59514,G59515,G59516,G59517,G59518,G59519,G59520,
       G59521,G59522,G59523,G59524,G59525,G59526,G59527,G59528,G59529,G59530,G59531,G59532,G59533,G59534,G59535,G59536,G59537,G59538,G59539,G59540,
       G59541,G59542,G59543,G59544,G59545,G59546,G59547,G59548,G59549,G59550,G59551,G59552,G59553,G59554,G59555,G59556,G59557,G59558,G59559,G59560,
       G59561,G59562,G59563,G59564,G59565,G59566,G59567,G59568,G59569,G59570,G59571,G59572,G59573,G59574,G59575,G59576,G59577,G59578,G59579,G59580,
       G59581,G59582,G59583,G59584,G59585,G59586,G59587,G59588,G59589,G59590,G59591,G59592,G59593,G59594,G59595,G59596,G59597,G59598,G59599,G59600,
       G59601,G59602,G59603,G59604,G59605,G59606,G59607,G59608,G59609,G59610,G59611,G59612,G59613,G59614,G59615,G59616,G59617,G59618,G59619,G59620,
       G59621,G59622,G59623,G59624,G59625,G59626,G59627,G59628,G59629,G59630,G59631,G59632,G59633,G59634,G59635,G59636,G59637,G59638,G59639,G59640,
       G59641,G59642,G59643,G59644,G59645,G59646,G59647,G59648,G59649,G59650,G59651,G59652,G59653,G59654,G59655,G59656,G59657,G59658,G59659,G59660,
       G59661,G59662,G59663,G59664,G59665,G59666,G59667,G59668,G59669,G59670,G59671,G59672,G59673,G59674,G59675,G59676,G59677,G59678,G59679,G59680,
       G59681,G59682,G59683,G59684,G59685,G59686,G59687,G59688,G59689,G59690,G59691,G59692,G59693,G59694,G59695,G59696,G59697,G59698,G59699,G59700,
       G59701,G59702,G59703,G59704,G59705,G59706,G59707,G59708,G59709,G59710,G59711,G59712,G59713,G59714,G59715,G59716,G59717,G59718,G59719,G59720,
       G59721,G59722,G59723,G59724,G59725,G59726,G59727,G59728,G59729,G59730,G59731,G59732,G59733,G59734,G59735,G59736,G59737,G59738,G59739,G59740,
       G59741,G59742,G59743,G59744,G59745,G59746,G59747,G59748,G59749,G59750,G59751,G59752,G59753,G59754,G59755,G59756,G59757,G59758,G59759,G59760,
       G59761,G59762,G59763,G59764,G59765,G59766,G59767,G59768,G59769,G59770,G59771,G59772,G59773,G59774,G59775,G59776,G59777,G59778,G59779,G59780,
       G59781,G59782,G59783,G59784,G59785,G59786,G59787,G59788,G59789,G59790,G59791,G59792,G59793,G59794,G59795,G59796,G59797,G59798,G59799,G59800,
       G59801,G59802,G59803,G59804,G59805,G59806,G59807,G59808,G59809,G59810,G59811,G59812,G59813,G59814,G59815,G59816,G59817,G59818,G59819,G59820,
       G59821,G59822,G59823,G59824,G59825,G59826,G59827,G59828,G59829,G59830,G59831,G59832,G59833,G59834,G59835,G59836,G59837,G59838,G59839,G59840,
       G59841,G59842,G59843,G59844,G59845,G59846,G59847,G59848,G59849,G59850,G59851,G59852,G59853,G59854,G59855,G59856,G59857,G59858,G59859,G59860,
       G59861,G59862,G59863,G59864,G59865,G59866,G59867,G59868,G59869,G59870,G59871,G59872,G59873,G59874,G59875,G59876,G59877,G59878,G59879,G59880,
       G59881,G59882,G59883,G59884,G59885,G59886,G59887,G59888,G59889,G59890,G59891,G59892,G59893,G59894,G59895,G59896,G59897,G59898,G59899,G59900,
       G59901,G59902,G59903,G59904,G59905,G59906,G59907,G59908,G59909,G59910,G59911,G59912,G59913,G59914,G59915,G59916,G59917,G59918,G59919,G59920,
       G59921,G59922,G59923,G59924,G59925,G59926,G59927,G59928,G59929,G59930,G59931,G59932,G59933,G59934,G59935,G59936,G59937,G59938,G59939,G59940,
       G59941,G59942,G59943,G59944,G59945,G59946,G59947,G59948,G59949,G59950,G59951,G59952,G59953,G59954,G59955,G59956,G59957,G59958,G59959,G59960,
       G59961,G59962,G59963,G59964,G59965,G59966,G59967,G59968,G59969,G59970,G59971,G59972,G59973,G59974,G59975,G59976,G59977,G59978,G59979,G59980,
       G59981,G59982,G59983,G59984,G59985,G59986,G59987,G59988,G59989,G59990,G59991,G59992,G59993,G59994,G59995,G59996,G59997,G59998,G59999,G60000,
       G60001,G60002,G60003,G60004,G60005,G60006,G60007,G60008,G60009,G60010,G60011,G60012,G60013,G60014,G60015,G60016,G60017,G60018,G60019,G60020,
       G60021,G60022,G60023,G60024,G60025,G60026,G60027,G60028,G60029,G60030,G60031,G60032,G60033,G60034,G60035,G60036,G60037,G60038,G60039,G60040,
       G60041,G60042,G60043,G60044,G60045,G60046,G60047,G60048,G60049,G60050,G60051,G60052,G60053,G60054,G60055,G60056,G60057,G60058,G60059,G60060,
       G60061,G60062,G60063,G60064,G60065,G60066,G60067,G60068,G60069,G60070,G60071,G60072,G60073,G60074,G60075,G60076,G60077,G60078,G60079,G60080,
       G60081,G60082,G60083,G60084,G60085,G60086,G60087,G60088,G60089,G60090,G60091,G60092,G60093,G60094,G60095,G60096,G60097,G60098,G60099,G60100,
       G60101,G60102,G60103,G60104,G60105,G60106,G60107,G60108,G60109,G60110,G60111,G60112,G60113,G60114,G60115,G60116,G60117,G60118,G60119,G60120,
       G60121,G60122,G60123,G60124,G60125,G60126,G60127,G60128,G60129,G60130,G60131,G60132,G60133,G60134,G60135,G60136,G60137,G60138,G60139,G60140,
       G60141,G60142,G60143,G60144,G60145,G60146,G60147,G60148,G60149,G60150,G60151,G60152,G60153,G60154,G60155,G60156,G60157,G60158,G60159,G60160,
       G60161,G60162,G60163,G60164,G60165,G60166,G60167,G60168,G60169,G60170,G60171,G60172,G60173,G60174,G60175,G60176,G60177,G60178,G60179,G60180,
       G60181,G60182,G60183,G60184,G60185,G60186,G60187,G60188,G60189,G60190,G60191,G60192,G60193,G60194,G60195,G60196,G60197,G60198,G60199,G60200,
       G60201,G60202,G60203,G60204,G60205,G60206,G60207,G60208,G60209,G60210,G60211,G60212,G60213,G60214,G60215,G60216,G60217,G60218,G60219,G60220,
       G60221,G60222,G60223,G60224,G60225,G60226,G60227,G60228,G60229,G60230,G60231,G60232,G60233,G60234,G60235,G60236,G60237,G60238,G60239,G60240,
       G60241,G60242,G60243,G60244,G60245,G60246,G60247,G60248,G60249,G60250,G60251,G60252,G60253,G60254,G60255,G60256,G60257,G60258,G60259,G60260,
       G60261,G60262,G60263,G60264,G60265,G60266,G60267,G60268,G60269,G60270,G60271,G60272,G60273,G60274,G60275,G60276,G60277,G60278,G60279,G60280,
       G60281,G60282,G60283,G60284,G60285,G60286,G60287,G60288,G60289,G60290,G60291,G60292,G60293,G60294,G60295,G60296,G60297,G60298,G60299,G60300,
       G60301,G60302,G60303,G60304,G60305,G60306,G60307,G60308,G60309,G60310,G60311,G60312,G60313,G60314,G60315,G60316,G60317,G60318,G60319,G60320,
       G60321,G60322,G60323,G60324,G60325,G60326,G60327,G60328,G60329,G60330,G60331,G60332,G60333,G60334,G60335,G60336,G60337,G60338,G60339,G60340,
       G60341,G60342,G60343,G60344,G60345,G60346,G60347,G60348,G60349,G60350,G60351,G60352,G60353,G60354,G60355,G60356,G60357,G60358,G60359,G60360,
       G60361,G60362,G60363,G60364,G60365,G60366,G60367,G60368,G60369,G60370,G60371,G60372,G60373,G60374,G60375,G60376,G60377,G60378,G60379,G60380,
       G60381,G60382,G60383,G60384,G60385,G60386,G60387,G60388,G60389,G60390,G60391,G60392,G60393,G60394,G60395,G60396,G60397,G60398,G60399,G60400,
       G60401,G60402,G60403,G60404,G60405,G60406,G60407,G60408,G60409,G60410,G60411,G60412,G60413,G60414,G60415,G60416,G60417,G60418,G60419,G60420,
       G60421,G60422,G60423,G60424,G60425,G60426,G60427,G60428,G60429,G60430,G60431,G60432,G60433,G60434,G60435,G60436,G60437,G60438,G60439,G60440,
       G60441,G60442,G60443,G60444,G60445,G60446,G60447,G60448,G60449,G60450,G60451,G60452,G60453,G60454,G60455,G60456,G60457,G60458,G60459,G60460,
       G60461,G60462,G60463,G60464,G60465,G60466,G60467,G60468,G60469,G60470,G60471,G60472,G60473,G60474,G60475,G60476,G60477,G60478,G60479,G60480,
       G60481,G60482,G60483,G60484,G60485,G60486,G60487,G60488,G60489,G60490,G60491,G60492,G60493,G60494,G60495,G60496,G60497,G60498,G60499,G60500,
       G60501,G60502,G60503,G60504,G60505,G60506,G60507,G60508,G60509,G60510,G60511,G60512,G60513,G60514,G60515,G60516,G60517,G60518,G60519,G60520,
       G60521,G60522,G60523,G60524,G60525,G60526,G60527,G60528,G60529,G60530,G60531,G60532,G60533,G60534,G60535,G60536,G60537,G60538,G60539,G60540,
       G60541,G60542,G60543,G60544,G60545,G60546,G60547,G60548,G60549,G60550,G60551,G60552,G60553,G60554,G60555,G60556,G60557,G60558,G60559,G60560,
       G60561,G60562,G60563,G60564,G60565,G60566,G60567,G60568,G60569,G60570,G60571,G60572,G60573,G60574,G60575,G60576,G60577,G60578,G60579,G60580,
       G60581,G60582,G60583,G60584,G60585,G60586,G60587,G60588,G60589,G60590,G60591,G60592,G60593,G60594,G60595,G60596,G60597,G60598,G60599,G60600,
       G60601,G60602,G60603,G60604,G60605,G60606,G60607,G60608,G60609,G60610,G60611,G60612,G60613,G60614,G60615,G60616,G60617,G60618,G60619,G60620,
       G60621,G60622,G60623,G60624,G60625,G60626,G60627,G60628,G60629,G60630,G60631,G60632,G60633,G60634,G60635,G60636,G60637,G60638,G60639,G60640,
       G60641,G60642,G60643,G60644,G60645,G60646,G60647,G60648,G60649,G60650,G60651,G60652,G60653,G60654,G60655,G60656,G60657,G60658,G60659,G60660,
       G60661,G60662,G60663,G60664,G60665,G60666,G60667,G60668,G60669,G60670,G60671,G60672,G60673,G60674,G60675,G60676,G60677,G60678,G60679,G60680,
       G60681,G60682,G60683,G60684,G60685,G60686,G60687,G60688,G60689,G60690,G60691,G60692,G60693,G60694,G60695,G60696,G60697,G60698,G60699,G60700,
       G60701,G60702,G60703,G60704,G60705,G60706,G60707,G60708,G60709,G60710,G60711,G60712,G60713,G60714,G60715,G60716,G60717,G60718,G60719,G60720,
       G60721,G60722,G60723,G60724,G60725,G60726,G60727,G60728,G60729,G60730,G60731,G60732,G60733,G60734,G60735,G60736,G60737,G60738,G60739,G60740,
       G60741,G60742,G60743,G60744,G60745,G60746,G60747,G60748,G60749,G60750,G60751,G60752,G60753,G60754,G60755,G60756,G60757,G60758,G60759,G60760,
       G60761,G60762,G60763,G60764,G60765,G60766,G60767,G60768,G60769,G60770,G60771,G60772,G60773,G60774,G60775,G60776,G60777,G60778,G60779,G60780,
       G60781,G60782,G60783,G60784,G60785,G60786,G60787,G60788,G60789,G60790,G60791,G60792,G60793,G60794,G60795,G60796,G60797,G60798,G60799,G60800,
       G60801,G60802,G60803,G60804,G60805,G60806,G60807,G60808,G60809,G60810,G60811,G60812,G60813,G60814,G60815,G60816,G60817,G60818,G60819,G60820,
       G60821,G60822,G60823,G60824,G60825,G60826,G60827,G60828,G60829,G60830,G60831,G60832,G60833,G60834,G60835,G60836,G60837,G60838,G60839,G60840,
       G60841,G60842,G60843,G60844,G60845,G60846,G60847,G60848,G60849,G60850,G60851,G60852,G60853,G60854,G60855,G60856,G60857,G60858,G60859,G60860,
       G60861,G60862,G60863,G60864,G60865,G60866,G60867,G60868,G60869,G60870,G60871,G60872,G60873,G60874,G60875,G60876,G60877,G60878,G60879,G60880,
       G60881,G60882,G60883,G60884,G60885,G60886,G60887,G60888,G60889,G60890,G60891,G60892,G60893,G60894,G60895,G60896,G60897,G60898,G60899,G60900,
       G60901,G60902,G60903,G60904,G60905,G60906,G60907,G60908,G60909,G60910,G60911,G60912,G60913,G60914,G60915,G60916,G60917,G60918,G60919,G60920,
       G60921,G60922,G60923,G60924,G60925,G60926,G60927,G60928,G60929,G60930,G60931,G60932,G60933,G60934,G60935,G60936,G60937,G60938,G60939,G60940,
       G60941,G60942,G60943,G60944,G60945,G60946,G60947,G60948,G60949,G60950,G60951,G60952,G60953,G60954,G60955,G60956,G60957,G60958,G60959,G60960,
       G60961,G60962,G60963,G60964,G60965,G60966,G60967,G60968,G60969,G60970,G60971,G60972,G60973,G60974,G60975,G60976,G60977,G60978,G60979,G60980,
       G60981,G60982,G60983,G60984,G60985,G60986,G60987,G60988,G60989,G60990,G60991,G60992,G60993,G60994,G60995,G60996,G60997,G60998,G60999,G61000,
       G61001,G61002,G61003,G61004,G61005,G61006,G61007,G61008,G61009,G61010,G61011,G61012,G61013,G61014,G61015,G61016,G61017,G61018,G61019,G61020,
       G61021,G61022,G61023,G61024,G61025,G61026,G61027,G61028,G61029,G61030,G61031,G61032,G61033,G61034,G61035,G61036,G61037,G61038,G61039,G61040,
       G61041,G61042,G61043,G61044,G61045,G61046,G61047,G61048,G61049,G61050,G61051,G61052,G61053,G61054,G61055,G61056,G61057,G61058,G61059,G61060,
       G61061,G61062,G61063,G61064,G61065,G61066,G61067,G61068,G61069,G61070,G61071,G61072,G61073,G61074,G61075,G61076,G61077,G61078,G61079,G61080,
       G61081,G61082,G61083,G61084,G61085,G61086,G61087,G61088,G61089,G61090,G61091,G61092,G61093,G61094,G61095,G61096,G61097,G61098,G61099,G61100,
       G61101,G61102,G61103,G61104,G61105,G61106,G61107,G61108,G61109,G61110,G61111,G61112,G61113,G61114,G61115,G61116,G61117,G61118,G61119,G61120,
       G61121,G61122,G61123,G61124,G61125,G61126,G61127,G61128,G61129,G61130,G61131,G61132,G61133,G61134,G61135,G61136,G61137,G61138,G61139,G61140,
       G61141,G61142,G61143,G61144,G61145,G61146,G61147,G61148,G61149,G61150,G61151,G61152,G61153,G61154,G61155,G61156,G61157,G61158,G61159,G61160,
       G61161,G61162,G61163,G61164,G61165,G61166,G61167,G61168,G61169,G61170,G61171,G61172,G61173,G61174,G61175,G61176,G61177,G61178,G61179,G61180,
       G61181,G61182,G61183,G61184,G61185,G61186,G61187,G61188,G61189,G61190,G61191,G61192,G61193,G61194,G61195,G61196,G61197,G61198,G61199,G61200,
       G61201,G61202,G61203,G61204,G61205,G61206,G61207,G61208,G61209,G61210,G61211,G61212,G61213,G61214,G61215,G61216,G61217,G61218,G61219,G61220,
       G61221,G61222,G61223,G61224,G61225,G61226,G61227,G61228,G61229,G61230,G61231,G61232,G61233,G61234,G61235,G61236,G61237,G61238,G61239,G61240,
       G61241,G61242,G61243,G61244,G61245,G61246,G61247,G61248,G61249,G61250,G61251,G61252,G61253,G61254,G61255,G61256,G61257,G61258,G61259,G61260,
       G61261,G61262,G61263,G61264,G61265,G61266,G61267,G61268,G61269,G61270,G61271,G61272,G61273,G61274,G61275,G61276,G61277,G61278,G61279,G61280,
       G61281,G61282,G61283,G61284,G61285,G61286,G61287,G61288,G61289,G61290,G61291,G61292,G61293,G61294,G61295,G61296,G61297,G61298,G61299,G61300,
       G61301,G61302,G61303,G61304,G61305,G61306,G61307,G61308,G61309,G61310,G61311,G61312,G61313,G61314,G61315,G61316,G61317,G61318,G61319,G61320,
       G61321,G61322,G61323,G61324,G61325,G61326,G61327,G61328,G61329,G61330,G61331,G61332,G61333,G61334,G61335,G61336,G61337,G61338,G61339,G61340,
       G61341,G61342,G61343,G61344,G61345,G61346,G61347,G61348,G61349,G61350,G61351,G61352,G61353,G61354,G61355,G61356,G61357,G61358,G61359,G61360,
       G61361,G61362,G61363,G61364,G61365,G61366,G61367,G61368,G61369,G61370,G61371,G61372,G61373,G61374,G61375,G61376,G61377,G61378,G61379,G61380,
       G61381,G61382,G61383,G61384,G61385,G61386,G61387,G61388,G61389,G61390,G61391,G61392,G61393,G61394,G61395,G61396,G61397,G61398,G61399,G61400,
       G61401,G61402,G61403,G61404,G61405,G61406,G61407,G61408,G61409,G61410,G61411,G61412,G61413,G61414,G61415,G61416,G61417,G61418,G61419,G61420,
       G61421,G61422,G61423,G61424,G61425,G61426,G61427,G61428,G61429,G61430,G61431,G61432,G61433,G61434,G61435,G61436,G61437,G61438,G61439,G61440,
       G61441,G61442,G61443,G61444,G61445,G61446,G61447,G61448,G61449,G61450,G61451,G61452,G61453,G61454,G61455,G61456,G61457,G61458,G61459,G61460,
       G61461,G61462,G61463,G61464,G61465,G61466,G61467,G61468,G61469,G61470,G61471,G61472,G61473,G61474,G61475,G61476,G61477,G61478,G61479,G61480,
       G61481,G61482,G61483,G61484,G61485,G61486,G61487,G61488,G61489,G61490,G61491,G61492,G61493,G61494,G61495,G61496,G61497,G61498,G61499,G61500,
       G61501,G61502,G61503,G61504,G61505,G61506,G61507,G61508,G61509,G61510,G61511,G61512,G61513,G61514,G61515,G61516,G61517,G61518,G61519,G61520,
       G61521,G61522,G61523,G61524,G61525,G61526,G61527,G61528,G61529,G61530,G61531,G61532,G61533,G61534,G61535,G61536,G61537,G61538,G61539,G61540,
       G61541,G61542,G61543,G61544,G61545,G61546,G61547,G61548,G61549,G61550,G61551,G61552,G61553,G61554,G61555,G61556,G61557,G61558,G61559,G61560,
       G61561,G61562,G61563,G61564,G61565,G61566,G61567,G61568,G61569,G61570,G61571,G61572,G61573,G61574,G61575,G61576,G61577,G61578,G61579,G61580,
       G61581,G61582,G61583,G61584,G61585,G61586,G61587,G61588,G61589,G61590,G61591,G61592,G61593,G61594,G61595,G61596,G61597,G61598,G61599,G61600,
       G61601,G61602,G61603,G61604,G61605,G61606,G61607,G61608,G61609,G61610,G61611,G61612,G61613,G61614,G61615,G61616,G61617,G61618,G61619,G61620,
       G61621,G61622,G61623,G61624,G61625,G61626,G61627,G61628,G61629,G61630,G61631,G61632,G61633,G61634,G61635,G61636,G61637,G61638,G61639,G61640,
       G61641,G61642,G61643,G61644,G61645,G61646,G61647,G61648,G61649,G61650,G61651,G61652,G61653,G61654,G61655,G61656,G61657,G61658,G61659,G61660,
       G61661,G61662,G61663,G61664,G61665,G61666,G61667,G61668,G61669,G61670,G61671,G61672,G61673,G61674,G61675,G61676,G61677,G61678,G61679,G61680,
       G61681,G61682,G61683,G61684,G61685,G61686,G61687,G61688,G61689,G61690,G61691,G61692,G61693,G61694,G61695,G61696,G61697,G61698,G61699,G61700,
       G61701,G61702,G61703,G61704,G61705,G61706,G61707,G61708,G61709,G61710,G61711,G61712,G61713,G61714,G61715,G61716,G61717,G61718,G61719,G61720,
       G61721,G61722,G61723,G61724,G61725,G61726,G61727,G61728,G61729,G61730,G61731,G61732,G61733,G61734,G61735,G61736,G61737,G61738,G61739,G61740,
       G61741,G61742,G61743,G61744,G61745,G61746,G61747,G61748,G61749,G61750,G61751,G61752,G61753,G61754,G61755,G61756,G61757,G61758,G61759,G61760,
       G61761,G61762,G61763,G61764,G61765,G61766,G61767,G61768,G61769,G61770,G61771,G61772,G61773,G61774,G61775,G61776,G61777,G61778,G61779,G61780,
       G61781,G61782,G61783,G61784,G61785,G61786,G61787,G61788,G61789,G61790,G61791,G61792,G61793,G61794,G61795,G61796,G61797,G61798,G61799,G61800,
       G61801,G61802,G61803,G61804,G61805,G61806,G61807,G61808,G61809,G61810,G61811,G61812,G61813,G61814,G61815,G61816,G61817,G61818,G61819,G61820,
       G61821,G61822,G61823,G61824,G61825,G61826,G61827,G61828,G61829,G61830,G61831,G61832,G61833,G61834,G61835,G61836,G61837,G61838,G61839,G61840,
       G61841,G61842,G61843,G61844,G61845,G61846,G61847,G61848,G61849,G61850,G61851,G61852,G61853,G61854,G61855,G61856,G61857,G61858,G61859,G61860,
       G61861,G61862,G61863,G61864,G61865,G61866,G61867,G61868,G61869,G61870,G61871,G61872,G61873,G61874,G61875,G61876,G61877,G61878,G61879,G61880,
       G61881,G61882,G61883,G61884,G61885,G61886,G61887,G61888,G61889,G61890,G61891,G61892,G61893,G61894,G61895,G61896,G61897,G61898,G61899,G61900,
       G61901,G61902,G61903,G61904,G61905,G61906,G61907,G61908,G61909,G61910,G61911,G61912,G61913,G61914,G61915,G61916,G61917,G61918,G61919,G61920,
       G61921,G61922,G61923,G61924,G61925,G61926,G61927,G61928,G61929,G61930,G61931,G61932,G61933,G61934,G61935,G61936,G61937,G61938,G61939,G61940,
       G61941,G61942,G61943,G61944,G61945,G61946,G61947,G61948,G61949,G61950,G61951,G61952,G61953,G61954,G61955,G61956,G61957,G61958,G61959,G61960,
       G61961,G61962,G61963,G61964,G61965,G61966,G61967,G61968,G61969,G61970,G61971,G61972,G61973,G61974,G61975,G61976,G61977,G61978,G61979,G61980,
       G61981,G61982,G61983,G61984,G61985,G61986,G61987,G61988,G61989,G61990,G61991,G61992,G61993,G61994,G61995,G61996,G61997,G61998,G61999,G62000,
       G62001,G62002,G62003,G62004,G62005,G62006,G62007,G62008,G62009,G62010,G62011,G62012,G62013,G62014,G62015,G62016,G62017,G62018,G62019,G62020,
       G62021,G62022,G62023,G62024,G62025,G62026,G62027,G62028,G62029,G62030,G62031,G62032,G62033,G62034,G62035,G62036,G62037,G62038,G62039,G62040,
       G62041,G62042,G62043,G62044,G62045,G62046,G62047,G62048,G62049,G62050,G62051,G62052,G62053,G62054,G62055,G62056,G62057,G62058,G62059,G62060,
       G62061,G62062,G62063,G62064,G62065,G62066,G62067,G62068,G62069,G62070,G62071,G62072,G62073,G62074,G62075,G62076,G62077,G62078,G62079,G62080,
       G62081,G62082,G62083,G62084,G62085,G62086,G62087,G62088,G62089,G62090,G62091,G62092,G62093,G62094,G62095,G62096,G62097,G62098,G62099,G62100,
       G62101,G62102,G62103,G62104,G62105,G62106,G62107,G62108,G62109,G62110,G62111,G62112,G62113,G62114,G62115,G62116,G62117,G62118,G62119,G62120,
       G62121,G62122,G62123,G62124,G62125,G62126,G62127,G62128,G62129,G62130,G62131,G62132,G62133,G62134,G62135,G62136,G62137,G62138,G62139,G62140,
       G62141,G62142,G62143,G62144,G62145,G62146,G62147,G62148,G62149,G62150,G62151,G62152,G62153,G62154,G62155,G62156,G62157,G62158,G62159,G62160,
       G62161,G62162,G62163,G62164,G62165,G62166,G62167,G62168,G62169,G62170,G62171,G62172,G62173,G62174,G62175,G62176,G62177,G62178,G62179,G62180,
       G62181,G62182,G62183,G62184,G62185,G62186,G62187,G62188,G62189,G62190,G62191,G62192,G62193,G62194,G62195,G62196,G62197,G62198,G62199,G62200,
       G62201,G62202,G62203,G62204,G62205,G62206,G62207,G62208,G62209,G62210,G62211,G62212,G62213,G62214,G62215,G62216,G62217,G62218,G62219,G62220,
       G62221,G62222,G62223,G62224,G62225,G62226,G62227,G62228,G62229,G62230,G62231,G62232,G62233,G62234,G62235,G62236,G62237,G62238,G62239,G62240,
       G62241,G62242,G62243,G62244,G62245,G62246,G62247,G62248,G62249,G62250,G62251,G62252,G62253,G62254,G62255,G62256,G62257,G62258,G62259,G62260,
       G62261,G62262,G62263,G62264,G62265,G62266,G62267,G62268,G62269,G62270,G62271,G62272,G62273,G62274,G62275,G62276,G62277,G62278,G62279,G62280,
       G62281,G62282,G62283,G62284,G62285,G62286,G62287,G62288,G62289,G62290,G62291,G62292,G62293,G62294,G62295,G62296,G62297,G62298,G62299,G62300,
       G62301,G62302,G62303,G62304,G62305,G62306,G62307,G62308,G62309,G62310,G62311,G62312,G62313,G62314,G62315,G62316,G62317,G62318,G62319,G62320,
       G62321,G62322,G62323,G62324,G62325,G62326,G62327,G62328,G62329,G62330,G62331,G62332,G62333,G62334,G62335,G62336,G62337,G62338,G62339,G62340,
       G62341,G62342,G62343,G62344,G62345,G62346,G62347,G62348,G62349,G62350,G62351,G62352,G62353,G62354,G62355,G62356,G62357,G62358,G62359,G62360,
       G62361,G62362,G62363,G62364,G62365,G62366,G62367,G62368,G62369,G62370,G62371,G62372,G62373,G62374,G62375,G62376,G62377,G62378,G62379,G62380,
       G62381,G62382,G62383,G62384,G62385,G62386,G62387,G62388,G62389,G62390,G62391,G62392,G62393,G62394,G62395,G62396,G62397,G62398,G62399,G62400,
       G62401,G62402,G62403,G62404,G62405,G62406,G62407,G62408,G62409,G62410,G62411,G62412,G62413,G62414,G62415,G62416,G62417,G62418,G62419,G62420,
       G62421,G62422,G62423,G62424,G62425,G62426,G62427,G62428,G62429,G62430,G62431,G62432,G62433,G62434,G62435,G62436,G62437,G62438,G62439,G62440,
       G62441,G62442,G62443,G62444,G62445,G62446,G62447,G62448,G62449,G62450,G62451,G62452,G62453,G62454,G62455,G62456,G62457,G62458,G62459,G62460,
       G62461,G62462,G62463,G62464,G62465,G62466,G62467,G62468,G62469,G62470,G62471,G62472,G62473,G62474,G62475,G62476,G62477,G62478,G62479,G62480,
       G62481,G62482,G62483,G62484,G62485,G62486,G62487,G62488,G62489,G62490,G62491,G62492,G62493,G62494,G62495,G62496,G62497,G62498,G62499,G62500,
       G62501,G62502,G62503,G62504,G62505,G62506,G62507,G62508,G62509,G62510,G62511,G62512,G62513,G62514,G62515,G62516,G62517,G62518,G62519,G62520,
       G62521,G62522,G62523,G62524,G62525,G62526,G62527,G62528,G62529,G62530,G62531,G62532,G62533,G62534,G62535,G62536,G62537,G62538,G62539,G62540,
       G62541,G62542,G62543,G62544,G62545,G62546,G62547,G62548,G62549,G62550,G62551,G62552,G62553,G62554,G62555,G62556,G62557,G62558,G62559,G62560,
       G62561,G62562,G62563,G62564,G62565,G62566,G62567,G62568,G62569,G62570,G62571,G62572,G62573,G62574,G62575,G62576,G62577,G62578,G62579,G62580,
       G62581,G62582,G62583,G62584,G62585,G62586,G62587,G62588,G62589,G62590,G62591,G62592,G62593,G62594,G62595,G62596,G62597,G62598,G62599,G62600,
       G62601,G62602,G62603,G62604,G62605,G62606,G62607,G62608,G62609,G62610,G62611,G62612,G62613,G62614,G62615,G62616,G62617,G62618,G62619,G62620,
       G62621,G62622,G62623,G62624,G62625,G62626,G62627,G62628,G62629,G62630,G62631,G62632,G62633,G62634,G62635,G62636,G62637,G62638,G62639,G62640,
       G62641,G62642,G62643,G62644,G62645,G62646,G62647,G62648,G62649,G62650,G62651,G62652,G62653,G62654,G62655,G62656,G62657,G62658,G62659,G62660,
       G62661,G62662,G62663,G62664,G62665,G62666,G62667,G62668,G62669,G62670,G62671,G62672,G62673,G62674,G62675,G62676,G62677,G62678,G62679,G62680,
       G62681,G62682,G62683,G62684,G62685,G62686,G62687,G62688,G62689,G62690,G62691,G62692,G62693,G62694,G62695,G62696,G62697,G62698,G62699,G62700,
       G62701,G62702,G62703,G62704,G62705,G62706,G62707,G62708,G62709,G62710,G62711,G62712,G62713,G62714,G62715,G62716,G62717,G62718,G62719,G62720,
       G62721,G62722,G62723,G62724,G62725,G62726,G62727,G62728,G62729,G62730,G62731,G62732,G62733,G62734,G62735,G62736,G62737,G62738,G62739,G62740,
       G62741,G62742,G62743,G62744,G62745,G62746,G62747,G62748,G62749,G62750,G62751,G62752,G62753,G62754,G62755,G62756,G62757,G62758,G62759,G62760,
       G62761,G62762,G62763,G62764,G62765,G62766,G62767,G62768,G62769,G62770,G62771,G62772,G62773,G62774,G62775,G62776,G62777,G62778,G62779,G62780,
       G62781,G62782,G62783,G62784,G62785,G62786,G62787,G62788,G62789,G62790,G62791,G62792,G62793,G62794,G62795,G62796,G62797,G62798,G62799,G62800,
       G62801,G62802,G62803,G62804,G62805,G62806,G62807,G62808,G62809,G62810,G62811,G62812,G62813,G62814,G62815,G62816,G62817,G62818,G62819,G62820,
       G62821,G62822,G62823,G62824,G62825,G62826,G62827,G62828,G62829,G62830,G62831,G62832,G62833,G62834,G62835,G62836,G62837,G62838,G62839,G62840,
       G62841,G62842,G62843,G62844,G62845,G62846,G62847,G62848,G62849,G62850,G62851,G62852,G62853,G62854,G62855,G62856,G62857,G62858,G62859,G62860,
       G62861,G62862,G62863,G62864,G62865,G62866,G62867,G62868,G62869,G62870,G62871,G62872,G62873,G62874,G62875,G62876,G62877,G62878,G62879,G62880,
       G62881,G62882,G62883,G62884,G62885,G62886,G62887,G62888,G62889,G62890,G62891,G62892,G62893,G62894,G62895,G62896,G62897,G62898,G62899,G62900,
       G62901,G62902,G62903,G62904,G62905,G62906,G62907,G62908,G62909,G62910,G62911,G62912,G62913,G62914,G62915,G62916,G62917,G62918,G62919,G62920,
       G62921,G62922,G62923,G62924,G62925,G62926,G62927,G62928,G62929,G62930,G62931,G62932,G62933,G62934,G62935,G62936,G62937,G62938,G62939,G62940,
       G62941,G62942,G62943,G62944,G62945,G62946,G62947,G62948,G62949,G62950,G62951,G62952,G62953,G62954,G62955,G62956,G62957,G62958,G62959,G62960,
       G62961,G62962,G62963,G62964,G62965,G62966,G62967,G62968,G62969,G62970,G62971,G62972,G62973,G62974,G62975,G62976,G62977,G62978,G62979,G62980,
       G62981,G62982,G62983,G62984,G62985,G62986,G62987,G62988,G62989,G62990,G62991,G62992,G62993,G62994,G62995,G62996,G62997,G62998,G62999,G63000,
       G63001,G63002,G63003,G63004,G63005,G63006,G63007,G63008,G63009,G63010,G63011,G63012,G63013,G63014,G63015,G63016,G63017,G63018,G63019,G63020,
       G63021,G63022,G63023,G63024,G63025,G63026,G63027,G63028,G63029,G63030,G63031,G63032,G63033,G63034,G63035,G63036,G63037,G63038,G63039,G63040,
       G63041,G63042,G63043,G63044,G63045,G63046,G63047,G63048,G63049,G63050,G63051,G63052,G63053,G63054,G63055,G63056,G63057,G63058,G63059,G63060,
       G63061,G63062,G63063,G63064,G63065,G63066,G63067,G63068,G63069,G63070,G63071,G63072,G63073,G63074,G63075,G63076,G63077,G63078,G63079,G63080,
       G63081,G63082,G63083,G63084,G63085,G63086,G63087,G63088,G63089,G63090,G63091,G63092,G63093,G63094,G63095,G63096,G63097,G63098,G63099,G63100,
       G63101,G63102,G63103,G63104,G63105,G63106,G63107,G63108,G63109,G63110,G63111,G63112,G63113,G63114,G63115,G63116,G63117,G63118,G63119,G63120,
       G63121,G63122,G63123,G63124,G63125,G63126,G63127,G63128,G63129,G63130,G63131,G63132,G63133,G63134,G63135,G63136,G63137,G63138,G63139,G63140,
       G63141,G63142,G63143,G63144,G63145,G63146,G63147,G63148,G63149,G63150,G63151,G63152,G63153,G63154,G63155,G63156,G63157,G63158,G63159,G63160,
       G63161,G63162,G63163,G63164,G63165,G63166,G63167,G63168,G63169,G63170,G63171,G63172,G63173,G63174,G63175,G63176,G63177,G63178,G63179,G63180,
       G63181,G63182,G63183,G63184,G63185,G63186,G63187,G63188,G63189,G63190,G63191,G63192,G63193,G63194,G63195,G63196,G63197,G63198,G63199,G63200,
       G63201,G63202,G63203,G63204,G63205,G63206,G63207,G63208,G63209,G63210,G63211,G63212,G63213,G63214,G63215,G63216,G63217,G63218,G63219,G63220,
       G63221,G63222,G63223,G63224,G63225,G63226,G63227,G63228,G63229,G63230,G63231,G63232,G63233,G63234,G63235,G63236,G63237,G63238,G63239,G63240,
       G63241,G63242,G63243,G63244,G63245,G63246,G63247,G63248,G63249,G63250,G63251,G63252,G63253,G63254,G63255,G63256,G63257,G63258,G63259,G63260,
       G63261,G63262,G63263,G63264,G63265,G63266,G63267,G63268,G63269,G63270,G63271,G63272,G63273,G63274,G63275,G63276,G63277,G63278,G63279,G63280,
       G63281,G63282,G63283,G63284,G63285,G63286,G63287,G63288,G63289,G63290,G63291,G63292,G63293,G63294,G63295,G63296,G63297,G63298,G63299,G63300,
       G63301,G63302,G63303,G63304,G63305,G63306,G63307,G63308,G63309,G63310,G63311,G63312,G63313,G63314,G63315,G63316,G63317,G63318,G63319,G63320,
       G63321,G63322,G63323,G63324,G63325,G63326,G63327,G63328,G63329,G63330,G63331,G63332,G63333,G63334,G63335,G63336,G63337,G63338,G63339,G63340,
       G63341,G63342,G63343,G63344,G63345,G63346,G63347,G63348,G63349,G63350,G63351,G63352,G63353,G63354,G63355,G63356,G63357,G63358,G63359,G63360,
       G63361,G63362,G63363,G63364,G63365,G63366,G63367,G63368,G63369,G63370,G63371,G63372,G63373,G63374,G63375,G63376,G63377,G63378,G63379,G63380,
       G63381,G63382,G63383,G63384,G63385,G63386,G63387,G63388,G63389,G63390,G63391,G63392,G63393,G63394,G63395,G63396,G63397,G63398,G63399,G63400,
       G63401,G63402,G63403,G63404,G63405,G63406,G63407,G63408,G63409,G63410,G63411,G63412,G63413,G63414,G63415,G63416,G63417,G63418,G63419,G63420,
       G63421,G63422,G63423,G63424,G63425,G63426,G63427,G63428,G63429,G63430,G63431,G63432,G63433,G63434,G63435,G63436,G63437,G63438,G63439,G63440,
       G63441,G63442,G63443,G63444,G63445,G63446,G63447,G63448,G63449,G63450,G63451,G63452,G63453,G63454,G63455,G63456,G63457,G63458,G63459,G63460,
       G63461,G63462,G63463,G63464,G63465,G63466,G63467,G63468,G63469,G63470,G63471,G63472,G63473,G63474,G63475,G63476,G63477,G63478,G63479,G63480,
       G63481,G63482,G63483,G63484,G63485,G63486,G63487,G63488,G63489,G63490,G63491,G63492,G63493,G63494,G63495,G63496,G63497,G63498,G63499,G63500,
       G63501,G63502,G63503,G63504,G63505,G63506,G63507,G63508,G63509,G63510,G63511,G63512,G63513,G63514,G63515,G63516,G63517,G63518,G63519,G63520,
       G63521,G63522,G63523,G63524,G63525,G63526,G63527,G63528,G63529,G63530,G63531,G63532,G63533,G63534,G63535,G63536,G63537,G63538,G63539,G63540,
       G63541,G63542,G63543,G63544,G63545,G63546,G63547,G63548,G63549,G63550,G63551,G63552,G63553,G63554,G63555,G63556,G63557,G63558,G63559,G63560,
       G63561,G63562,G63563,G63564,G63565,G63566,G63567,G63568,G63569,G63570,G63571,G63572,G63573,G63574,G63575,G63576,G63577,G63578,G63579,G63580,
       G63581,G63582,G63583,G63584,G63585,G63586,G63587,G63588,G63589,G63590,G63591,G63592,G63593,G63594,G63595,G63596,G63597,G63598,G63599,G63600,
       G63601,G63602,G63603,G63604,G63605,G63606,G63607,G63608,G63609,G63610,G63611,G63612,G63613,G63614,G63615,G63616,G63617,G63618,G63619,G63620,
       G63621,G63622,G63623,G63624,G63625,G63626,G63627,G63628,G63629,G63630,G63631,G63632,G63633,G63634,G63635,G63636,G63637,G63638,G63639,G63640,
       G63641,G63642,G63643,G63644,G63645,G63646,G63647,G63648,G63649,G63650,G63651,G63652,G63653,G63654,G63655,G63656,G63657,G63658,G63659,G63660,
       G63661,G63662,G63663,G63664,G63665,G63666,G63667,G63668,G63669,G63670,G63671,G63672,G63673,G63674,G63675,G63676,G63677,G63678,G63679,G63680,
       G63681,G63682,G63683,G63684,G63685,G63686,G63687,G63688,G63689,G63690,G63691,G63692,G63693,G63694,G63695,G63696,G63697,G63698,G63699,G63700,
       G63701,G63702,G63703,G63704,G63705,G63706,G63707,G63708,G63709,G63710,G63711,G63712,G63713,G63714,G63715,G63716,G63717,G63718,G63719,G63720,
       G63721,G63722,G63723,G63724,G63725,G63726,G63727,G63728,G63729,G63730,G63731,G63732,G63733,G63734,G63735,G63736,G63737,G63738,G63739,G63740,
       G63741,G63742,G63743,G63744,G63745,G63746,G63747,G63748,G63749,G63750,G63751,G63752,G63753,G63754,G63755,G63756,G63757,G63758,G63759,G63760,
       G63761,G63762,G63763,G63764,G63765,G63766,G63767,G63768,G63769,G63770,G63771,G63772,G63773,G63774,G63775,G63776,G63777,G63778,G63779,G63780,
       G63781,G63782,G63783,G63784,G63785,G63786,G63787,G63788,G63789,G63790,G63791,G63792,G63793,G63794,G63795,G63796,G63797,G63798,G63799,G63800,
       G63801,G63802,G63803,G63804,G63805,G63806,G63807,G63808,G63809,G63810,G63811,G63812,G63813,G63814,G63815,G63816,G63817,G63818,G63819,G63820,
       G63821,G63822,G63823,G63824,G63825,G63826,G63827,G63828,G63829,G63830,G63831,G63832,G63833,G63834,G63835,G63836,G63837,G63838,G63839,G63840,
       G63841,G63842,G63843,G63844,G63845,G63846,G63847,G63848,G63849,G63850,G63851,G63852,G63853,G63854,G63855,G63856,G63857,G63858,G63859,G63860,
       G63861,G63862,G63863,G63864,G63865,G63866,G63867,G63868,G63869,G63870,G63871,G63872,G63873,G63874,G63875,G63876,G63877,G63878,G63879,G63880,
       G63881,G63882,G63883,G63884,G63885,G63886,G63887,G63888,G63889,G63890,G63891,G63892,G63893,G63894,G63895,G63896,G63897,G63898,G63899,G63900,
       G63901,G63902,G63903,G63904,G63905,G63906,G63907,G63908,G63909,G63910,G63911,G63912,G63913,G63914,G63915,G63916,G63917,G63918,G63919,G63920,
       G63921,G63922,G63923,G63924,G63925,G63926,G63927,G63928,G63929,G63930,G63931,G63932,G63933,G63934,G63935,G63936,G63937,G63938,G63939,G63940,
       G63941,G63942,G63943,G63944,G63945,G63946,G63947,G63948,G63949,G63950,G63951,G63952,G63953,G63954,G63955,G63956,G63957,G63958,G63959,G63960,
       G63961,G63962,G63963,G63964,G63965,G63966,G63967,G63968,G63969,G63970,G63971,G63972,G63973,G63974,G63975,G63976,G63977,G63978,G63979,G63980,
       G63981,G63982,G63983,G63984,G63985,G63986,G63987,G63988,G63989,G63990,G63991,G63992,G63993,G63994,G63995,G63996,G63997,G63998,G63999,G64000,
       G64001,G64002,G64003,G64004,G64005,G64006,G64007,G64008,G64009,G64010,G64011,G64012,G64013,G64014,G64015,G64016,G64017,G64018,G64019,G64020,
       G64021,G64022,G64023,G64024,G64025,G64026,G64027,G64028,G64029,G64030,G64031,G64032,G64033,G64034,G64035,G64036,G64037,G64038,G64039,G64040,
       G64041,G64042,G64043,G64044,G64045,G64046,G64047,G64048,G64049,G64050,G64051,G64052,G64053,G64054,G64055,G64056,G64057,G64058,G64059,G64060,
       G64061,G64062,G64063,G64064,G64065,G64066,G64067,G64068,G64069,G64070,G64071,G64072,G64073,G64074,G64075,G64076,G64077,G64078,G64079,G64080,
       G64081,G64082,G64083,G64084,G64085,G64086,G64087,G64088,G64089,G64090,G64091,G64092,G64093,G64094,G64095,G64096,G64097,G64098,G64099,G64100,
       G64101,G64102,G64103,G64104,G64105,G64106,G64107,G64108,G64109,G64110,G64111,G64112,G64113,G64114,G64115,G64116,G64117,G64118,G64119,G64120,
       G64121,G64122,G64123,G64124,G64125,G64126,G64127,G64128,G64129,G64130,G64131,G64132,G64133,G64134,G64135,G64136,G64137,G64138,G64139,G64140,
       G64141,G64142,G64143,G64144,G64145,G64146,G64147,G64148,G64149,G64150,G64151,G64152,G64153,G64154,G64155,G64156,G64157,G64158,G64159,G64160,
       G64161,G64162,G64163,G64164,G64165,G64166,G64167,G64168,G64169,G64170,G64171,G64172,G64173,G64174,G64175,G64176,G64177,G64178,G64179,G64180,
       G64181,G64182,G64183,G64184,G64185,G64186,G64187,G64188,G64189,G64190,G64191,G64192,G64193,G64194,G64195,G64196,G64197,G64198,G64199,G64200,
       G64201,G64202,G64203,G64204,G64205,G64206,G64207,G64208,G64209,G64210,G64211,G64212,G64213,G64214,G64215,G64216,G64217,G64218,G64219,G64220,
       G64221,G64222,G64223,G64224,G64225,G64226,G64227,G64228,G64229,G64230,G64231,G64232,G64233,G64234,G64235,G64236,G64237,G64238,G64239,G64240,
       G64241,G64242,G64243,G64244,G64245,G64246,G64247,G64248,G64249,G64250,G64251,G64252,G64253,G64254,G64255,G64256,G64257,G64258,G64259,G64260,
       G64261,G64262,G64263,G64264,G64265,G64266,G64267,G64268,G64269,G64270,G64271,G64272,G64273,G64274,G64275,G64276,G64277,G64278,G64279,G64280,
       G64281,G64282,G64283,G64284,G64285,G64286,G64287,G64288,G64289,G64290,G64291,G64292,G64293,G64294,G64295,G64296,G64297,G64298,G64299,G64300,
       G64301,G64302,G64303,G64304,G64305,G64306,G64307,G64308,G64309,G64310,G64311,G64312,G64313,G64314,G64315,G64316,G64317,G64318,G64319,G64320,
       G64321,G64322,G64323,G64324,G64325,G64326,G64327,G64328,G64329,G64330,G64331,G64332,G64333,G64334,G64335,G64336,G64337,G64338,G64339,G64340,
       G64341,G64342,G64343,G64344,G64345,G64346,G64347,G64348,G64349,G64350,G64351,G64352,G64353,G64354,G64355,G64356,G64357,G64358,G64359,G64360,
       G64361,G64362,G64363,G64364,G64365,G64366,G64367,G64368,G64369,G64370,G64371,G64372,G64373,G64374,G64375,G64376,G64377,G64378,G64379,G64380,
       G64381,G64382,G64383,G64384,G64385,G64386,G64387,G64388,G64389,G64390,G64391,G64392,G64393,G64394,G64395,G64396,G64397,G64398,G64399,G64400,
       G64401,G64402,G64403,G64404,G64405,G64406,G64407,G64408,G64409,G64410,G64411,G64412,G64413,G64414,G64415,G64416,G64417,G64418,G64419,G64420,
       G64421,G64422,G64423,G64424,G64425,G64426,G64427,G64428,G64429,G64430,G64431,G64432,G64433,G64434,G64435,G64436,G64437,G64438,G64439,G64440,
       G64441,G64442,G64443,G64444,G64445,G64446,G64447,G64448,G64449,G64450,G64451,G64452,G64453,G64454,G64455,G64456,G64457,G64458,G64459,G64460,
       G64461,G64462,G64463,G64464,G64465,G64466,G64467,G64468,G64469,G64470,G64471,G64472,G64473,G64474,G64475,G64476,G64477,G64478,G64479,G64480,
       G64481,G64482,G64483,G64484,G64485,G64486,G64487,G64488,G64489,G64490,G64491,G64492,G64493,G64494,G64495,G64496,G64497,G64498,G64499,G64500,
       G64501,G64502,G64503,G64504,G64505,G64506,G64507,G64508,G64509,G64510,G64511,G64512,G64513,G64514,G64515,G64516,G64517,G64518,G64519,G64520,
       G64521,G64522,G64523,G64524,G64525,G64526,G64527,G64528,G64529,G64530,G64531,G64532,G64533,G64534,G64535,G64536,G64537,G64538,G64539,G64540,
       G64541,G64542,G64543,G64544,G64545,G64546,G64547,G64548,G64549,G64550,G64551,G64552,G64553,G64554,G64555,G64556,G64557,G64558,G64559,G64560,
       G64561,G64562,G64563,G64564,G64565,G64566,G64567,G64568,G64569,G64570,G64571,G64572,G64573,G64574,G64575,G64576,G64577,G64578,G64579,G64580,
       G64581,G64582,G64583,G64584,G64585,G64586,G64587,G64588,G64589,G64590,G64591,G64592,G64593,G64594,G64595,G64596,G64597,G64598,G64599,G64600,
       G64601,G64602,G64603,G64604,G64605,G64606,G64607,G64608,G64609,G64610,G64611,G64612,G64613,G64614,G64615,G64616,G64617,G64618,G64619,G64620,
       G64621,G64622,G64623,G64624,G64625,G64626,G64627,G64628,G64629,G64630,G64631,G64632,G64633,G64634,G64635,G64636,G64637,G64638,G64639,G64640,
       G64641,G64642,G64643,G64644,G64645,G64646,G64647,G64648,G64649,G64650,G64651,G64652,G64653,G64654,G64655,G64656,G64657,G64658,G64659,G64660,
       G64661,G64662,G64663,G64664,G64665,G64666,G64667,G64668,G64669,G64670,G64671,G64672,G64673,G64674,G64675,G64676,G64677,G64678,G64679,G64680,
       G64681,G64682,G64683,G64684,G64685,G64686,G64687,G64688,G64689,G64690,G64691,G64692,G64693,G64694,G64695,G64696,G64697,G64698,G64699,G64700,
       G64701,G64702,G64703,G64704,G64705,G64706,G64707,G64708,G64709,G64710,G64711,G64712,G64713,G64714,G64715,G64716,G64717,G64718,G64719,G64720,
       G64721,G64722,G64723,G64724,G64725,G64726,G64727,G64728,G64729,G64730,G64731,G64732,G64733,G64734,G64735,G64736,G64737,G64738,G64739,G64740,
       G64741,G64742,G64743,G64744,G64745,G64746,G64747,G64748,G64749,G64750,G64751,G64752,G64753,G64754,G64755,G64756,G64757,G64758,G64759,G64760,
       G64761,G64762,G64763,G64764,G64765,G64766,G64767,G64768,G64769,G64770,G64771,G64772,G64773,G64774,G64775,G64776,G64777,G64778,G64779,G64780,
       G64781,G64782,G64783,G64784,G64785,G64786,G64787,G64788,G64789,G64790,G64791,G64792,G64793,G64794,G64795,G64796,G64797,G64798,G64799,G64800,
       G64801,G64802,G64803,G64804,G64805,G64806,G64807,G64808,G64809,G64810,G64811,G64812,G64813,G64814,G64815,G64816,G64817,G64818,G64819,G64820,
       G64821,G64822,G64823,G64824,G64825,G64826,G64827,G64828,G64829,G64830,G64831,G64832,G64833,G64834,G64835,G64836,G64837,G64838,G64839,G64840,
       G64841,G64842,G64843,G64844,G64845,G64846,G64847,G64848,G64849,G64850,G64851,G64852,G64853,G64854,G64855,G64856,G64857,G64858,G64859,G64860,
       G64861,G64862,G64863,G64864,G64865,G64866,G64867,G64868,G64869,G64870,G64871,G64872,G64873,G64874,G64875,G64876,G64877,G64878,G64879,G64880,
       G64881,G64882,G64883,G64884,G64885,G64886,G64887,G64888,G64889,G64890,G64891,G64892,G64893,G64894,G64895,G64896,G64897,G64898,G64899,G64900,
       G64901,G64902,G64903,G64904,G64905,G64906,G64907,G64908,G64909,G64910,G64911,G64912,G64913,G64914,G64915,G64916,G64917,G64918,G64919,G64920,
       G64921,G64922,G64923,G64924,G64925,G64926,G64927,G64928,G64929,G64930,G64931,G64932,G64933,G64934,G64935,G64936,G64937,G64938,G64939,G64940,
       G64941,G64942,G64943,G64944,G64945,G64946,G64947,G64948,G64949,G64950,G64951,G64952,G64953,G64954,G64955,G64956,G64957,G64958,G64959,G64960,
       G64961,G64962,G64963,G64964,G64965,G64966,G64967,G64968,G64969,G64970,G64971,G64972,G64973,G64974,G64975,G64976,G64977,G64978,G64979,G64980,
       G64981,G64982,G64983,G64984,G64985,G64986,G64987,G64988,G64989,G64990,G64991,G64992,G64993,G64994,G64995,G64996,G64997,G64998,G64999,G65000,
       G65001,G65002,G65003,G65004,G65005,G65006,G65007,G65008,G65009,G65010,G65011,G65012,G65013,G65014,G65015,G65016,G65017,G65018,G65019,G65020,
       G65021,G65022,G65023,G65024,G65025,G65026,G65027,G65028,G65029,G65030,G65031,G65032,G65033,G65034,G65035,G65036,G65037,G65038,G65039,G65040,
       G65041,G65042,G65043,G65044,G65045,G65046,G65047,G65048,G65049,G65050,G65051,G65052,G65053,G65054,G65055,G65056,G65057,G65058,G65059,G65060,
       G65061,G65062,G65063,G65064,G65065,G65066,G65067,G65068,G65069,G65070,G65071,G65072,G65073,G65074,G65075,G65076,G65077,G65078,G65079,G65080,
       G65081,G65082,G65083,G65084,G65085,G65086,G65087,G65088,G65089,G65090,G65091,G65092,G65093,G65094,G65095,G65096,G65097,G65098,G65099,G65100,
       G65101,G65102,G65103,G65104,G65105,G65106,G65107,G65108,G65109,G65110,G65111,G65112,G65113,G65114,G65115,G65116,G65117,G65118,G65119,G65120,
       G65121,G65122,G65123,G65124,G65125,G65126,G65127,G65128,G65129,G65130,G65131,G65132,G65133,G65134,G65135,G65136,G65137,G65138,G65139,G65140,
       G65141,G65142,G65143,G65144,G65145,G65146,G65147,G65148,G65149,G65150,G65151,G65152,G65153,G65154,G65155,G65156,G65157,G65158,G65159,G65160,
       G65161,G65162,G65163,G65164,G65165,G65166,G65167,G65168,G65169,G65170,G65171,G65172,G65173,G65174,G65175,G65176,G65177,G65178,G65179,G65180,
       G65181,G65182,G65183,G65184,G65185,G65186,G65187,G65188,G65189,G65190,G65191,G65192,G65193,G65194,G65195,G65196,G65197,G65198,G65199,G65200,
       G65201,G65202,G65203,G65204,G65205,G65206,G65207,G65208,G65209,G65210,G65211,G65212,G65213,G65214,G65215,G65216,G65217,G65218,G65219,G65220,
       G65221,G65222,G65223,G65224,G65225,G65226,G65227,G65228,G65229,G65230,G65231,G65232,G65233,G65234,G65235,G65236,G65237,G65238,G65239,G65240,
       G65241,G65242,G65243,G65244,G65245,G65246,G65247,G65248,G65249,G65250,G65251,G65252,G65253,G65254,G65255,G65256,G65257,G65258,G65259,G65260,
       G65261,G65262,G65263,G65264,G65265,G65266,G65267,G65268,G65269,G65270,G65271,G65272,G65273,G65274,G65275,G65276,G65277,G65278,G65279,G65280,
       G65281,G65282,G65283,G65284,G65285,G65286,G65287,G65288,G65289,G65290,G65291,G65292,G65293,G65294,G65295,G65296,G65297,G65298,G65299,G65300,
       G65301,G65302,G65303,G65304,G65305,G65306,G65307,G65308,G65309,G65310,G65311,G65312,G65313,G65314,G65315,G65316,G65317,G65318,G65319,G65320,
       G65321,G65322,G65323,G65324,G65325,G65326,G65327,G65328,G65329,G65330,G65331,G65332,G65333,G65334,G65335,G65336,G65337,G65338,G65339,G65340,
       G65341,G65342,G65343,G65344,G65345,G65346,G65347,G65348,G65349,G65350,G65351,G65352,G65353,G65354,G65355,G65356,G65357,G65358,G65359,G65360,
       G65361,G65362,G65363,G65364,G65365,G65366,G65367,G65368,G65369,G65370,G65371,G65372,G65373,G65374,G65375,G65376,G65377,G65378,G65379,G65380,
       G65381,G65382,G65383,G65384,G65385,G65386,G65387,G65388,G65389,G65390,G65391,G65392,G65393,G65394,G65395,G65396,G65397,G65398,G65399,G65400,
       G65401,G65402,G65403,G65404,G65405,G65406,G65407,G65408,G65409,G65410,G65411,G65412,G65413,G65414,G65415,G65416,G65417,G65418,G65419,G65420,
       G65421,G65422,G65423,G65424,G65425,G65426,G65427,G65428,G65429,G65430,G65431,G65432,G65433,G65434,G65435,G65436,G65437,G65438,G65439,G65440,
       G65441,G65442,G65443,G65444,G65445,G65446,G65447,G65448,G65449,G65450,G65451,G65452,G65453,G65454,G65455,G65456,G65457,G65458,G65459,G65460,
       G65461,G65462,G65463,G65464,G65465,G65466,G65467,G65468,G65469,G65470,G65471,G65472,G65473,G65474,G65475,G65476,G65477,G65478,G65479,G65480,
       G65481,G65482,G65483,G65484,G65485,G65486,G65487,G65488,G65489,G65490,G65491,G65492,G65493,G65494,G65495,G65496,G65497,G65498,G65499,G65500,
       G65501,G65502,G65503,G65504,G65505,G65506,G65507,G65508,G65509,G65510,G65511,G65512,G65513,G65514,G65515,G65516,G65517,G65518,G65519,G65520,
       G65521,G65522,G65523,G65524,G65525,G65526,G65527,G65528,G65529,G65530,G65531,G65532,G65533,G65534,G65535,G65536,G65537,G65538,G65539,G65540,
       G65541,G65542,G65543,G65544,G65545,G65546,G65547,G65548,G65549,G65550,G65551,G65552,G65553,G65554,G65555,G65556,G65557,G65558,G65559,G65560,
       G65561,G65562,G65563,G65564,G65565,G65566,G65567,G65568,G65569,G65570,G65571,G65572,G65573,G65574,G65575,G65576,G65577,G65578,G65579,G65580,
       G65581,G65582,G65583,G65584,G65585,G65586,G65587,G65588,G65589,G65590,G65591,G65592,G65593,G65594,G65595,G65596,G65597,G65598,G65599,G65600,
       G65601,G65602,G65603,G65604,G65605,G65606,G65607,G65608,G65609,G65610,G65611,G65612,G65613,G65614,G65615,G65616,G65617,G65618,G65619,G65620,
       G65621,G65622,G65623,G65624,G65625,G65626,G65627,G65628,G65629,G65630,G65631,G65632,G65633,G65634,G65635,G65636,G65637,G65638,G65639,G65640,
       G65641,G65642,G65643,G65644,G65645,G65646,G65647,G65648,G65649,G65650,G65651,G65652,G65653,G65654,G65655,G65656,G65657,G65658,G65659,G65660,
       G65661,G65662,G65663,G65664,G65665,G65666,G65667,G65668,G65669,G65670,G65671,G65672,G65673,G65674,G65675,G65676,G65677,G65678,G65679,G65680,
       G65681,G65682,G65683,G65684,G65685,G65686,G65687,G65688,G65689,G65690,G65691,G65692,G65693,G65694,G65695,G65696,G65697,G65698,G65699,G65700,
       G65701,G65702,G65703,G65704,G65705,G65706,G65707,G65708,G65709,G65710,G65711,G65712,G65713,G65714,G65715,G65716,G65717,G65718,G65719,G65720,
       G65721,G65722,G65723,G65724,G65725,G65726,G65727,G65728,G65729,G65730,G65731,G65732,G65733,G65734,G65735,G65736,G65737,G65738,G65739,G65740,
       G65741,G65742,G65743,G65744,G65745,G65746,G65747,G65748,G65749,G65750,G65751,G65752,G65753,G65754,G65755,G65756,G65757,G65758,G65759,G65760,
       G65761,G65762,G65763,G65764,G65765,G65766,G65767,G65768,G65769,G65770,G65771,G65772,G65773,G65774,G65775,G65776,G65777,G65778,G65779,G65780,
       G65781,G65782,G65783,G65784,G65785,G65786,G65787,G65788,G65789,G65790,G65791,G65792,G65793,G65794,G65795,G65796,G65797,G65798,G65799,G65800,
       G65801,G65802,G65803,G65804,G65805,G65806,G65807,G65808,G65809,G65810,G65811,G65812,G65813,G65814,G65815,G65816,G65817,G65818,G65819,G65820,
       G65821,G65822,G65823,G65824,G65825,G65826,G65827,G65828,G65829,G65830,G65831,G65832,G65833,G65834,G65835,G65836,G65837,G65838,G65839,G65840,
       G65841,G65842,G65843,G65844,G65845,G65846,G65847,G65848,G65849,G65850,G65851,G65852,G65853,G65854,G65855,G65856,G65857,G65858,G65859,G65860,
       G65861,G65862,G65863,G65864,G65865,G65866,G65867,G65868,G65869,G65870,G65871,G65872,G65873,G65874,G65875,G65876,G65877,G65878,G65879,G65880,
       G65881,G65882,G65883,G65884,G65885,G65886,G65887,G65888,G65889,G65890,G65891,G65892,G65893,G65894,G65895,G65896,G65897,G65898,G65899,G65900,
       G65901,G65902,G65903,G65904,G65905,G65906,G65907,G65908,G65909,G65910,G65911,G65912,G65913,G65914,G65915,G65916,G65917,G65918,G65919,G65920,
       G65921,G65922,G65923,G65924,G65925,G65926,G65927,G65928,G65929,G65930,G65931,G65932,G65933,G65934,G65935,G65936,G65937,G65938,G65939,G65940,
       G65941,G65942,G65943,G65944,G65945,G65946,G65947,G65948,G65949,G65950,G65951,G65952,G65953,G65954,G65955,G65956,G65957,G65958,G65959,G65960,
       G65961,G65962,G65963,G65964,G65965,G65966,G65967,G65968,G65969,G65970,G65971,G65972,G65973,G65974,G65975,G65976,G65977,G65978,G65979,G65980,
       G65981,G65982,G65983,G65984,G65985,G65986,G65987,G65988,G65989,G65990,G65991,G65992,G65993,G65994,G65995,G65996,G65997,G65998,G65999,G66000,
       G66001,G66002,G66003,G66004,G66005,G66006,G66007,G66008,G66009,G66010,G66011,G66012,G66013,G66014,G66015,G66016,G66017,G66018,G66019,G66020,
       G66021,G66022,G66023,G66024,G66025,G66026,G66027,G66028,G66029,G66030,G66031,G66032,G66033,G66034,G66035,G66036,G66037,G66038,G66039,G66040,
       G66041,G66042,G66043,G66044,G66045,G66046,G66047,G66048,G66049,G66050,G66051,G66052,G66053,G66054,G66055,G66056,G66057,G66058,G66059,G66060,
       G66061,G66062,G66063,G66064,G66065,G66066,G66067,G66068,G66069,G66070,G66071,G66072,G66073,G66074,G66075,G66076,G66077,G66078,G66079,G66080,
       G66081,G66082,G66083,G66084,G66085,G66086,G66087,G66088,G66089,G66090,G66091,G66092,G66093,G66094,G66095,G66096,G66097,G66098,G66099,G66100,
       G66101,G66102,G66103,G66104,G66105,G66106,G66107,G66108,G66109,G66110,G66111,G66112,G66113,G66114,G66115,G66116,G66117,G66118,G66119,G66120,
       G66121,G66122,G66123,G66124,G66125,G66126,G66127,G66128,G66129,G66130,G66131,G66132,G66133,G66134,G66135,G66136,G66137,G66138,G66139,G66140,
       G66141,G66142,G66143,G66144,G66145,G66146,G66147,G66148,G66149,G66150,G66151,G66152,G66153,G66154,G66155,G66156,G66157,G66158,G66159,G66160,
       G66161,G66162,G66163,G66164,G66165,G66166,G66167,G66168,G66169,G66170,G66171,G66172,G66173,G66174,G66175,G66176,G66177,G66178,G66179,G66180,
       G66181,G66182,G66183,G66184,G66185,G66186,G66187,G66188,G66189,G66190,G66191,G66192,G66193,G66194,G66195,G66196,G66197,G66198,G66199,G66200,
       G66201,G66202,G66203,G66204,G66205,G66206,G66207,G66208,G66209,G66210,G66211,G66212,G66213,G66214,G66215,G66216,G66217,G66218,G66219,G66220,
       G66221,G66222,G66223,G66224,G66225,G66226,G66227,G66228,G66229,G66230,G66231,G66232,G66233,G66234,G66235,G66236,G66237,G66238,G66239,G66240,
       G66241,G66242,G66243,G66244,G66245,G66246,G66247,G66248,G66249,G66250,G66251,G66252,G66253,G66254,G66255,G66256,G66257,G66258,G66259,G66260,
       G66261,G66262,G66263,G66264,G66265,G66266,G66267,G66268,G66269,G66270,G66271,G66272,G66273,G66274,G66275,G66276,G66277,G66278,G66279,G66280,
       G66281,G66282,G66283,G66284,G66285,G66286,G66287,G66288,G66289,G66290,G66291,G66292,G66293,G66294,G66295,G66296,G66297,G66298,G66299,G66300,
       G66301,G66302,G66303,G66304,G66305,G66306,G66307,G66308,G66309,G66310,G66311,G66312,G66313,G66314,G66315,G66316,G66317,G66318,G66319,G66320,
       G66321,G66322,G66323,G66324,G66325,G66326,G66327,G66328,G66329,G66330,G66331,G66332,G66333,G66334,G66335,G66336,G66337,G66338,G66339,G66340,
       G66341,G66342,G66343,G66344,G66345,G66346,G66347,G66348,G66349,G66350,G66351,G66352,G66353,G66354,G66355,G66356,G66357,G66358,G66359,G66360,
       G66361,G66362,G66363,G66364,G66365,G66366,G66367,G66368,G66369,G66370,G66371,G66372,G66373,G66374,G66375,G66376,G66377,G66378,G66379,G66380,
       G66381,G66382,G66383,G66384,G66385,G66386,G66387,G66388,G66389,G66390,G66391,G66392,G66393,G66394,G66395,G66396,G66397,G66398,G66399,G66400,
       G66401,G66402,G66403,G66404,G66405,G66406,G66407,G66408,G66409,G66410,G66411,G66412,G66413,G66414,G66415,G66416,G66417,G66418,G66419,G66420,
       G66421,G66422,G66423,G66424,G66425,G66426,G66427,G66428,G66429,G66430,G66431,G66432,G66433,G66434,G66435,G66436,G66437,G66438,G66439,G66440,
       G66441,G66442,G66443,G66444,G66445,G66446,G66447,G66448,G66449,G66450,G66451,G66452,G66453,G66454,G66455,G66456,G66457,G66458,G66459,G66460,
       G66461,G66462,G66463,G66464,G66465,G66466,G66467,G66468,G66469,G66470,G66471,G66472,G66473,G66474,G66475,G66476,G66477,G66478,G66479,G66480,
       G66481,G66482,G66483,G66484,G66485,G66486,G66487,G66488,G66489,G66490,G66491,G66492,G66493,G66494,G66495,G66496,G66497,G66498,G66499,G66500,
       G66501,G66502,G66503,G66504,G66505,G66506,G66507,G66508,G66509,G66510,G66511,G66512,G66513,G66514,G66515,G66516,G66517,G66518,G66519,G66520,
       G66521,G66522,G66523,G66524,G66525,G66526,G66527,G66528,G66529,G66530,G66531,G66532,G66533,G66534,G66535,G66536,G66537,G66538,G66539,G66540,
       G66541,G66542,G66543,G66544,G66545,G66546,G66547,G66548,G66549,G66550,G66551,G66552,G66553,G66554,G66555,G66556,G66557,G66558,G66559,G66560,
       G66561,G66562,G66563,G66564,G66565,G66566,G66567,G66568,G66569,G66570,G66571,G66572,G66573,G66574,G66575,G66576,G66577,G66578,G66579,G66580,
       G66581,G66582,G66583,G66584,G66585,G66586,G66587,G66588,G66589,G66590,G66591,G66592,G66593,G66594,G66595,G66596,G66597,G66598,G66599,G66600,
       G66601,G66602,G66603,G66604,G66605,G66606,G66607,G66608,G66609,G66610,G66611,G66612,G66613,G66614,G66615,G66616,G66617,G66618,G66619,G66620,
       G66621,G66622,G66623,G66624,G66625,G66626,G66627,G66628,G66629,G66630,G66631,G66632,G66633,G66634,G66635,G66636,G66637,G66638,G66639,G66640,
       G66641,G66642,G66643,G66644,G66645,G66646,G66647,G66648,G66649,G66650,G66651,G66652,G66653,G66654,G66655,G66656,G66657,G66658,G66659,G66660,
       G66661,G66662,G66663,G66664,G66665,G66666,G66667,G66668,G66669,G66670,G66671,G66672,G66673,G66674,G66675,G66676,G66677,G66678,G66679,G66680,
       G66681,G66682,G66683,G66684,G66685,G66686,G66687,G66688,G66689,G66690,G66691,G66692,G66693,G66694,G66695,G66696,G66697,G66698,G66699,G66700,
       G66701,G66702,G66703,G66704,G66705,G66706,G66707,G66708,G66709,G66710,G66711,G66712,G66713,G66714,G66715,G66716,G66717,G66718,G66719,G66720,
       G66721,G66722,G66723,G66724,G66725,G66726,G66727,G66728,G66729,G66730,G66731,G66732,G66733,G66734,G66735,G66736,G66737,G66738,G66739,G66740,
       G66741,G66742,G66743,G66744,G66745,G66746,G66747,G66748,G66749,G66750,G66751,G66752,G66753,G66754,G66755,G66756,G66757,G66758,G66759,G66760,
       G66761,G66762,G66763,G66764,G66765,G66766,G66767,G66768,G66769,G66770,G66771,G66772,G66773,G66774,G66775,G66776,G66777,G66778,G66779,G66780,
       G66781,G66782,G66783,G66784,G66785,G66786,G66787,G66788,G66789,G66790,G66791,G66792,G66793,G66794,G66795,G66796,G66797,G66798,G66799,G66800,
       G66801,G66802,G66803,G66804,G66805,G66806,G66807,G66808,G66809,G66810,G66811,G66812,G66813,G66814,G66815,G66816,G66817,G66818,G66819,G66820,
       G66821,G66822,G66823,G66824,G66825,G66826,G66827,G66828,G66829,G66830,G66831,G66832,G66833,G66834,G66835,G66836,G66837,G66838,G66839,G66840,
       G66841,G66842,G66843,G66844,G66845,G66846,G66847,G66848,G66849,G66850,G66851,G66852,G66853,G66854,G66855,G66856,G66857,G66858,G66859,G66860,
       G66861,G66862,G66863,G66864,G66865,G66866,G66867,G66868,G66869,G66870,G66871,G66872,G66873,G66874,G66875,G66876,G66877,G66878,G66879,G66880,
       G66881,G66882,G66883,G66884,G66885,G66886,G66887,G66888,G66889,G66890,G66891,G66892,G66893,G66894,G66895,G66896,G66897,G66898,G66899,G66900,
       G66901,G66902,G66903,G66904,G66905,G66906,G66907,G66908,G66909,G66910,G66911,G66912,G66913,G66914,G66915,G66916,G66917,G66918,G66919,G66920,
       G66921,G66922,G66923,G66924,G66925,G66926,G66927,G66928,G66929,G66930,G66931,G66932,G66933,G66934,G66935,G66936,G66937,G66938,G66939,G66940,
       G66941,G66942,G66943,G66944,G66945,G66946,G66947,G66948,G66949,G66950,G66951,G66952,G66953,G66954,G66955,G66956,G66957,G66958,G66959,G66960,
       G66961,G66962,G66963,G66964,G66965,G66966,G66967,G66968,G66969,G66970,G66971,G66972,G66973,G66974,G66975,G66976,G66977,G66978,G66979,G66980,
       G66981,G66982,G66983,G66984,G66985,G66986,G66987,G66988,G66989,G66990,G66991,G66992,G66993,G66994,G66995,G66996,G66997,G66998,G66999,G67000,
       G67001,G67002,G67003,G67004,G67005,G67006,G67007,G67008,G67009,G67010,G67011,G67012,G67013,G67014,G67015,G67016,G67017,G67018,G67019,G67020,
       G67021,G67022,G67023,G67024,G67025,G67026,G67027,G67028,G67029,G67030,G67031,G67032,G67033,G67034,G67035,G67036,G67037,G67038,G67039,G67040,
       G67041,G67042,G67043,G67044,G67045,G67046,G67047,G67048,G67049,G67050,G67051,G67052,G67053,G67054,G67055,G67056,G67057,G67058,G67059,G67060,
       G67061,G67062,G67063,G67064,G67065,G67066,G67067,G67068,G67069,G67070,G67071,G67072,G67073,G67074,G67075,G67076,G67077,G67078,G67079,G67080,
       G67081,G67082,G67083,G67084,G67085,G67086,G67087,G67088,G67089,G67090,G67091,G67092,G67093,G67094,G67095,G67096,G67097,G67098,G67099,G67100,
       G67101,G67102,G67103,G67104,G67105,G67106,G67107,G67108,G67109,G67110,G67111,G67112,G67113,G67114,G67115,G67116,G67117,G67118,G67119,G67120,
       G67121,G67122,G67123,G67124,G67125,G67126,G67127,G67128,G67129,G67130,G67131,G67132,G67133,G67134,G67135,G67136,G67137,G67138,G67139,G67140,
       G67141,G67142,G67143,G67144,G67145,G67146,G67147,G67148,G67149,G67150,G67151,G67152,G67153,G67154,G67155,G67156,G67157,G67158,G67159,G67160,
       G67161,G67162,G67163,G67164,G67165,G67166,G67167,G67168,G67169,G67170,G67171,G67172,G67173,G67174,G67175,G67176,G67177,G67178,G67179,G67180,
       G67181,G67182,G67183,G67184,G67185,G67186,G67187,G67188,G67189,G67190,G67191,G67192,G67193,G67194,G67195,G67196,G67197,G67198,G67199,G67200,
       G67201,G67202,G67203,G67204,G67205,G67206,G67207,G67208,G67209,G67210,G67211,G67212,G67213,G67214,G67215,G67216,G67217,G67218,G67219,G67220,
       G67221,G67222,G67223,G67224,G67225,G67226,G67227,G67228,G67229,G67230,G67231,G67232,G67233,G67234,G67235,G67236,G67237,G67238,G67239,G67240,
       G67241,G67242,G67243,G67244,G67245,G67246,G67247,G67248,G67249,G67250,G67251,G67252,G67253,G67254,G67255,G67256,G67257,G67258,G67259,G67260,
       G67261,G67262,G67263,G67264,G67265,G67266,G67267,G67268,G67269,G67270,G67271,G67272,G67273,G67274,G67275,G67276,G67277,G67278,G67279,G67280,
       G67281,G67282,G67283,G67284,G67285,G67286,G67287,G67288,G67289,G67290,G67291,G67292,G67293,G67294,G67295,G67296,G67297,G67298,G67299,G67300,
       G67301,G67302,G67303,G67304,G67305,G67306,G67307,G67308,G67309,G67310,G67311,G67312,G67313,G67314,G67315,G67316,G67317,G67318,G67319,G67320,
       G67321,G67322,G67323,G67324,G67325,G67326,G67327,G67328,G67329,G67330,G67331,G67332,G67333,G67334,G67335,G67336,G67337,G67338,G67339,G67340,
       G67341,G67342,G67343,G67344,G67345,G67346,G67347,G67348,G67349,G67350,G67351,G67352,G67353,G67354,G67355,G67356,G67357,G67358,G67359,G67360,
       G67361,G67362,G67363,G67364,G67365,G67366,G67367,G67368,G67369,G67370,G67371,G67372,G67373,G67374,G67375,G67376,G67377,G67378,G67379,G67380,
       G67381,G67382,G67383,G67384,G67385,G67386,G67387,G67388,G67389,G67390,G67391,G67392,G67393,G67394,G67395,G67396,G67397,G67398,G67399,G67400,
       G67401,G67402,G67403,G67404,G67405,G67406,G67407,G67408,G67409,G67410,G67411,G67412,G67413,G67414,G67415,G67416,G67417,G67418,G67419,G67420,
       G67421,G67422,G67423,G67424,G67425,G67426,G67427,G67428,G67429,G67430,G67431,G67432,G67433,G67434,G67435,G67436,G67437,G67438,G67439,G67440,
       G67441,G67442,G67443,G67444,G67445,G67446,G67447,G67448,G67449,G67450,G67451,G67452,G67453,G67454,G67455,G67456,G67457,G67458,G67459,G67460,
       G67461,G67462,G67463,G67464,G67465,G67466,G67467,G67468,G67469,G67470,G67471,G67472,G67473,G67474,G67475,G67476,G67477,G67478,G67479,G67480,
       G67481,G67482,G67483,G67484,G67485,G67486,G67487,G67488,G67489,G67490,G67491,G67492,G67493,G67494,G67495,G67496,G67497,G67498,G67499,G67500,
       G67501,G67502,G67503,G67504,G67505,G67506,G67507,G67508,G67509,G67510,G67511,G67512,G67513,G67514,G67515,G67516,G67517,G67518,G67519,G67520,
       G67521,G67522,G67523,G67524,G67525,G67526,G67527,G67528,G67529,G67530,G67531,G67532,G67533,G67534,G67535,G67536,G67537,G67538,G67539,G67540,
       G67541,G67542,G67543,G67544,G67545,G67546,G67547,G67548,G67549,G67550,G67551,G67552,G67553,G67554,G67555,G67556,G67557,G67558,G67559,G67560,
       G67561,G67562,G67563,G67564,G67565,G67566,G67567,G67568,G67569,G67570,G67571,G67572,G67573,G67574,G67575,G67576,G67577,G67578,G67579,G67580,
       G67581,G67582,G67583,G67584,G67585,G67586,G67587,G67588,G67589,G67590,G67591,G67592,G67593,G67594,G67595,G67596,G67597,G67598,G67599,G67600,
       G67601,G67602,G67603,G67604,G67605,G67606,G67607,G67608,G67609,G67610,G67611,G67612,G67613,G67614,G67615,G67616,G67617,G67618,G67619,G67620,
       G67621,G67622,G67623,G67624,G67625,G67626,G67627,G67628,G67629,G67630,G67631,G67632,G67633,G67634,G67635,G67636,G67637,G67638,G67639,G67640,
       G67641,G67642,G67643,G67644,G67645,G67646,G67647,G67648,G67649,G67650,G67651,G67652,G67653,G67654,G67655,G67656,G67657,G67658,G67659,G67660,
       G67661,G67662,G67663,G67664,G67665,G67666,G67667,G67668,G67669,G67670,G67671,G67672,G67673,G67674,G67675,G67676,G67677,G67678,G67679,G67680,
       G67681,G67682,G67683,G67684,G67685,G67686,G67687,G67688,G67689,G67690,G67691,G67692,G67693,G67694,G67695,G67696,G67697,G67698,G67699,G67700,
       G67701,G67702,G67703,G67704,G67705,G67706,G67707,G67708,G67709,G67710,G67711,G67712,G67713,G67714,G67715,G67716,G67717,G67718,G67719,G67720,
       G67721,G67722,G67723,G67724,G67725,G67726,G67727,G67728,G67729,G67730,G67731,G67732,G67733,G67734,G67735,G67736,G67737,G67738,G67739,G67740,
       G67741,G67742,G67743,G67744,G67745,G67746,G67747,G67748,G67749,G67750,G67751,G67752,G67753,G67754,G67755,G67756,G67757,G67758,G67759,G67760,
       G67761,G67762,G67763,G67764,G67765,G67766,G67767,G67768,G67769,G67770,G67771,G67772,G67773,G67774,G67775,G67776,G67777,G67778,G67779,G67780,
       G67781,G67782,G67783,G67784,G67785,G67786,G67787,G67788,G67789,G67790,G67791,G67792,G67793,G67794,G67795,G67796,G67797,G67798,G67799,G67800,
       G67801,G67802,G67803,G67804,G67805,G67806,G67807,G67808,G67809,G67810,G67811,G67812,G67813,G67814,G67815,G67816,G67817,G67818,G67819,G67820,
       G67821,G67822,G67823,G67824,G67825,G67826,G67827,G67828,G67829,G67830,G67831,G67832,G67833,G67834,G67835,G67836,G67837,G67838,G67839,G67840,
       G67841,G67842,G67843,G67844,G67845,G67846,G67847,G67848,G67849,G67850,G67851,G67852,G67853,G67854,G67855,G67856,G67857,G67858,G67859,G67860,
       G67861,G67862,G67863,G67864,G67865,G67866,G67867,G67868,G67869,G67870,G67871,G67872,G67873,G67874,G67875,G67876,G67877,G67878,G67879,G67880,
       G67881,G67882,G67883,G67884,G67885,G67886,G67887,G67888,G67889,G67890,G67891,G67892,G67893,G67894,G67895,G67896,G67897,G67898,G67899,G67900,
       G67901,G67902,G67903,G67904,G67905,G67906,G67907,G67908,G67909,G67910,G67911,G67912,G67913,G67914,G67915,G67916,G67917,G67918,G67919,G67920,
       G67921,G67922,G67923,G67924,G67925,G67926,G67927,G67928,G67929,G67930,G67931,G67932,G67933,G67934,G67935,G67936,G67937,G67938,G67939,G67940,
       G67941,G67942,G67943,G67944,G67945,G67946,G67947,G67948,G67949,G67950,G67951,G67952,G67953,G67954,G67955,G67956,G67957,G67958,G67959,G67960,
       G67961,G67962,G67963,G67964,G67965,G67966,G67967,G67968,G67969,G67970,G67971,G67972,G67973,G67974,G67975,G67976,G67977,G67978,G67979,G67980,
       G67981,G67982,G67983,G67984,G67985,G67986,G67987,G67988,G67989,G67990,G67991,G67992,G67993,G67994,G67995,G67996,G67997,G67998,G67999,G68000,
       G68001,G68002,G68003,G68004,G68005,G68006,G68007,G68008,G68009,G68010,G68011,G68012,G68013,G68014,G68015,G68016,G68017,G68018,G68019,G68020,
       G68021,G68022,G68023,G68024,G68025,G68026,G68027,G68028,G68029,G68030,G68031,G68032,G68033,G68034,G68035,G68036,G68037,G68038,G68039,G68040,
       G68041,G68042,G68043,G68044,G68045,G68046,G68047,G68048,G68049,G68050,G68051,G68052,G68053,G68054,G68055,G68056,G68057,G68058,G68059,G68060,
       G68061,G68062,G68063,G68064,G68065,G68066,G68067,G68068,G68069,G68070,G68071,G68072,G68073,G68074,G68075,G68076,G68077,G68078,G68079,G68080,
       G68081,G68082,G68083,G68084,G68085,G68086,G68087,G68088,G68089,G68090,G68091,G68092,G68093,G68094,G68095,G68096,G68097,G68098,G68099,G68100,
       G68101,G68102,G68103,G68104,G68105,G68106,G68107,G68108,G68109,G68110,G68111,G68112,G68113,G68114,G68115,G68116,G68117,G68118,G68119,G68120,
       G68121,G68122,G68123,G68124,G68125,G68126,G68127,G68128,G68129,G68130,G68131,G68132,G68133,G68134,G68135,G68136,G68137,G68138,G68139,G68140,
       G68141,G68142,G68143,G68144,G68145,G68146,G68147,G68148,G68149,G68150,G68151,G68152,G68153,G68154,G68155,G68156,G68157,G68158,G68159,G68160,
       G68161,G68162,G68163,G68164,G68165,G68166,G68167,G68168,G68169,G68170,G68171,G68172,G68173,G68174,G68175,G68176,G68177,G68178,G68179,G68180,
       G68181,G68182,G68183,G68184,G68185,G68186,G68187,G68188,G68189,G68190,G68191,G68192,G68193,G68194,G68195,G68196,G68197,G68198,G68199,G68200,
       G68201,G68202,G68203,G68204,G68205,G68206,G68207,G68208,G68209,G68210,G68211,G68212,G68213,G68214,G68215,G68216,G68217,G68218,G68219,G68220,
       G68221,G68222,G68223,G68224,G68225,G68226,G68227,G68228,G68229,G68230,G68231,G68232,G68233,G68234,G68235,G68236,G68237,G68238,G68239,G68240,
       G68241,G68242,G68243,G68244,G68245,G68246,G68247,G68248,G68249,G68250,G68251,G68252,G68253,G68254,G68255,G68256,G68257,G68258,G68259,G68260,
       G68261,G68262,G68263,G68264,G68265,G68266,G68267,G68268,G68269,G68270,G68271,G68272,G68273,G68274,G68275,G68276,G68277,G68278,G68279,G68280,
       G68281,G68282,G68283,G68284,G68285,G68286,G68287,G68288,G68289,G68290,G68291,G68292,G68293,G68294,G68295,G68296,G68297,G68298,G68299,G68300,
       G68301,G68302,G68303,G68304,G68305,G68306,G68307,G68308,G68309,G68310,G68311,G68312,G68313,G68314,G68315,G68316,G68317,G68318,G68319,G68320,
       G68321,G68322,G68323,G68324,G68325,G68326,G68327,G68328,G68329,G68330,G68331,G68332,G68333,G68334,G68335,G68336,G68337,G68338,G68339,G68340,
       G68341,G68342,G68343,G68344,G68345,G68346,G68347,G68348,G68349,G68350,G68351,G68352,G68353,G68354,G68355,G68356,G68357,G68358,G68359,G68360,
       G68361,G68362,G68363,G68364,G68365,G68366,G68367,G68368,G68369,G68370,G68371,G68372,G68373,G68374,G68375,G68376,G68377,G68378,G68379,G68380,
       G68381,G68382,G68383,G68384,G68385,G68386,G68387,G68388,G68389,G68390,G68391,G68392,G68393,G68394,G68395,G68396,G68397,G68398,G68399,G68400,
       G68401,G68402,G68403,G68404,G68405,G68406,G68407,G68408,G68409,G68410,G68411,G68412,G68413,G68414,G68415,G68416,G68417,G68418,G68419,G68420,
       G68421,G68422,G68423,G68424,G68425,G68426,G68427,G68428,G68429,G68430,G68431,G68432,G68433,G68434,G68435,G68436,G68437,G68438,G68439,G68440,
       G68441,G68442,G68443,G68444,G68445,G68446,G68447,G68448,G68449,G68450,G68451,G68452,G68453,G68454,G68455,G68456,G68457,G68458,G68459,G68460,
       G68461,G68462,G68463,G68464,G68465,G68466,G68467,G68468,G68469,G68470,G68471,G68472,G68473,G68474,G68475,G68476,G68477,G68478,G68479,G68480,
       G68481,G68482,G68483,G68484,G68485,G68486,G68487,G68488,G68489,G68490,G68491,G68492,G68493,G68494,G68495,G68496,G68497,G68498,G68499,G68500,
       G68501,G68502,G68503,G68504,G68505,G68506,G68507,G68508,G68509,G68510,G68511,G68512,G68513,G68514,G68515,G68516,G68517,G68518,G68519,G68520,
       G68521,G68522,G68523,G68524,G68525,G68526,G68527,G68528,G68529,G68530,G68531,G68532,G68533,G68534,G68535,G68536,G68537,G68538,G68539,G68540,
       G68541,G68542,G68543,G68544,G68545,G68546,G68547,G68548,G68549,G68550,G68551,G68552,G68553,G68554,G68555,G68556,G68557,G68558,G68559,G68560,
       G68561,G68562,G68563,G68564,G68565,G68566,G68567,G68568,G68569,G68570,G68571,G68572,G68573,G68574,G68575,G68576,G68577,G68578,G68579,G68580,
       G68581,G68582,G68583,G68584,G68585,G68586,G68587,G68588,G68589,G68590,G68591,G68592,G68593,G68594,G68595,G68596,G68597,G68598,G68599,G68600,
       G68601,G68602,G68603,G68604,G68605,G68606,G68607,G68608,G68609,G68610,G68611,G68612,G68613,G68614,G68615,G68616,G68617,G68618,G68619,G68620,
       G68621,G68622,G68623,G68624,G68625,G68626,G68627,G68628,G68629,G68630,G68631,G68632,G68633,G68634,G68635,G68636,G68637,G68638,G68639,G68640,
       G68641,G68642,G68643,G68644,G68645,G68646,G68647,G68648,G68649,G68650,G68651,G68652,G68653,G68654,G68655,G68656,G68657,G68658,G68659,G68660,
       G68661,G68662,G68663,G68664,G68665,G68666,G68667,G68668,G68669,G68670,G68671,G68672,G68673,G68674,G68675,G68676,G68677,G68678,G68679,G68680,
       G68681,G68682,G68683,G68684,G68685,G68686,G68687,G68688,G68689,G68690,G68691,G68692,G68693,G68694,G68695,G68696,G68697,G68698,G68699,G68700,
       G68701,G68702,G68703,G68704,G68705,G68706,G68707,G68708,G68709,G68710,G68711,G68712,G68713,G68714,G68715,G68716,G68717,G68718,G68719,G68720,
       G68721,G68722,G68723,G68724,G68725,G68726,G68727,G68728,G68729,G68730,G68731,G68732,G68733,G68734,G68735,G68736,G68737,G68738,G68739,G68740,
       G68741,G68742,G68743,G68744,G68745,G68746,G68747,G68748,G68749,G68750,G68751,G68752,G68753,G68754,G68755,G68756,G68757,G68758,G68759,G68760,
       G68761,G68762,G68763,G68764,G68765,G68766,G68767,G68768,G68769,G68770,G68771,G68772,G68773,G68774,G68775,G68776,G68777,G68778,G68779,G68780,
       G68781,G68782,G68783,G68784,G68785,G68786,G68787,G68788,G68789,G68790,G68791,G68792,G68793,G68794,G68795,G68796,G68797,G68798,G68799,G68800,
       G68801,G68802,G68803,G68804,G68805,G68806,G68807,G68808,G68809,G68810,G68811,G68812,G68813,G68814,G68815,G68816,G68817,G68818,G68819,G68820,
       G68821,G68822,G68823,G68824,G68825,G68826,G68827,G68828,G68829,G68830,G68831,G68832,G68833,G68834,G68835,G68836,G68837,G68838,G68839,G68840,
       G68841,G68842,G68843,G68844,G68845,G68846,G68847,G68848,G68849,G68850,G68851,G68852,G68853,G68854,G68855,G68856,G68857,G68858,G68859,G68860,
       G68861,G68862,G68863,G68864,G68865,G68866,G68867,G68868,G68869,G68870,G68871,G68872,G68873,G68874,G68875,G68876,G68877,G68878,G68879,G68880,
       G68881,G68882,G68883,G68884,G68885,G68886,G68887,G68888,G68889,G68890,G68891,G68892,G68893,G68894,G68895,G68896,G68897,G68898,G68899,G68900,
       G68901,G68902,G68903,G68904,G68905,G68906,G68907,G68908,G68909,G68910,G68911,G68912,G68913,G68914,G68915,G68916,G68917,G68918,G68919,G68920,
       G68921,G68922,G68923,G68924,G68925,G68926,G68927,G68928,G68929,G68930,G68931,G68932,G68933,G68934,G68935,G68936,G68937,G68938,G68939,G68940,
       G68941,G68942,G68943,G68944,G68945,G68946,G68947,G68948,G68949,G68950,G68951,G68952,G68953,G68954,G68955,G68956,G68957,G68958,G68959,G68960,
       G68961,G68962,G68963,G68964,G68965,G68966,G68967,G68968,G68969,G68970,G68971,G68972,G68973,G68974,G68975,G68976,G68977,G68978,G68979,G68980,
       G68981,G68982,G68983,G68984,G68985,G68986,G68987,G68988,G68989,G68990,G68991,G68992,G68993,G68994,G68995,G68996,G68997,G68998,G68999,G69000,
       G69001,G69002,G69003,G69004,G69005,G69006,G69007,G69008,G69009,G69010,G69011,G69012,G69013,G69014,G69015,G69016,G69017,G69018,G69019,G69020,
       G69021,G69022,G69023,G69024,G69025,G69026,G69027,G69028,G69029,G69030,G69031,G69032,G69033,G69034,G69035,G69036,G69037,G69038,G69039,G69040,
       G69041,G69042,G69043,G69044,G69045,G69046,G69047,G69048,G69049,G69050,G69051,G69052,G69053,G69054,G69055,G69056,G69057,G69058,G69059,G69060,
       G69061,G69062,G69063,G69064,G69065,G69066,G69067,G69068,G69069,G69070,G69071,G69072,G69073,G69074,G69075,G69076,G69077,G69078,G69079,G69080,
       G69081,G69082,G69083,G69084,G69085,G69086,G69087,G69088,G69089,G69090,G69091,G69092,G69093,G69094,G69095,G69096,G69097,G69098,G69099,G69100,
       G69101,G69102,G69103,G69104,G69105,G69106,G69107,G69108,G69109,G69110,G69111,G69112,G69113,G69114,G69115,G69116,G69117,G69118,G69119,G69120,
       G69121,G69122,G69123,G69124,G69125,G69126,G69127,G69128,G69129,G69130,G69131,G69132,G69133,G69134,G69135,G69136,G69137,G69138,G69139,G69140,
       G69141,G69142,G69143,G69144,G69145,G69146,G69147,G69148,G69149,G69150,G69151,G69152,G69153,G69154,G69155,G69156,G69157,G69158,G69159,G69160,
       G69161,G69162,G69163,G69164,G69165,G69166,G69167,G69168,G69169,G69170,G69171,G69172,G69173,G69174,G69175,G69176,G69177,G69178,G69179,G69180,
       G69181,G69182,G69183,G69184,G69185,G69186,G69187,G69188,G69189,G69190,G69191,G69192,G69193,G69194,G69195,G69196,G69197,G69198,G69199,G69200,
       G69201,G69202,G69203,G69204,G69205,G69206,G69207,G69208,G69209,G69210,G69211,G69212,G69213,G69214,G69215,G69216,G69217,G69218,G69219,G69220,
       G69221,G69222,G69223,G69224,G69225,G69226,G69227,G69228,G69229,G69230,G69231,G69232,G69233,G69234,G69235,G69236,G69237,G69238,G69239,G69240,
       G69241,G69242,G69243,G69244,G69245,G69246,G69247,G69248,G69249,G69250,G69251,G69252,G69253,G69254,G69255,G69256,G69257,G69258,G69259,G69260,
       G69261,G69262,G69263,G69264,G69265,G69266,G69267,G69268,G69269,G69270,G69271,G69272,G69273,G69274,G69275,G69276,G69277,G69278,G69279,G69280,
       G69281,G69282,G69283,G69284,G69285,G69286,G69287,G69288,G69289,G69290,G69291,G69292,G69293,G69294,G69295,G69296,G69297,G69298,G69299,G69300,
       G69301,G69302,G69303,G69304,G69305,G69306,G69307,G69308,G69309,G69310,G69311,G69312,G69313,G69314,G69315,G69316,G69317,G69318,G69319,G69320,
       G69321,G69322,G69323,G69324,G69325,G69326,G69327,G69328,G69329,G69330,G69331,G69332,G69333,G69334,G69335,G69336,G69337,G69338,G69339,G69340,
       G69341,G69342,G69343,G69344,G69345,G69346,G69347,G69348,G69349,G69350,G69351,G69352,G69353,G69354,G69355,G69356,G69357,G69358,G69359,G69360,
       G69361,G69362,G69363,G69364,G69365,G69366,G69367,G69368,G69369,G69370,G69371,G69372,G69373,G69374,G69375,G69376,G69377,G69378,G69379,G69380,
       G69381,G69382,G69383,G69384,G69385,G69386,G69387,G69388,G69389,G69390,G69391,G69392,G69393,G69394,G69395,G69396,G69397,G69398,G69399,G69400,
       G69401,G69402,G69403,G69404,G69405,G69406,G69407,G69408,G69409,G69410,G69411,G69412,G69413,G69414,G69415,G69416,G69417,G69418,G69419,G69420,
       G69421,G69422,G69423,G69424,G69425,G69426,G69427,G69428,G69429,G69430,G69431,G69432,G69433,G69434,G69435,G69436,G69437,G69438,G69439,G69440,
       G69441,G69442,G69443,G69444,G69445,G69446,G69447,G69448,G69449,G69450,G69451,G69452,G69453,G69454,G69455,G69456,G69457,G69458,G69459,G69460,
       G69461,G69462,G69463,G69464,G69465,G69466,G69467,G69468,G69469,G69470,G69471,G69472,G69473,G69474,G69475,G69476,G69477,G69478,G69479,G69480,
       G69481,G69482,G69483,G69484,G69485,G69486,G69487,G69488,G69489,G69490,G69491,G69492,G69493,G69494,G69495,G69496,G69497,G69498,G69499,G69500,
       G69501,G69502,G69503,G69504,G69505,G69506,G69507,G69508,G69509,G69510,G69511,G69512,G69513,G69514,G69515,G69516,G69517,G69518,G69519,G69520,
       G69521,G69522,G69523,G69524,G69525,G69526,G69527,G69528,G69529,G69530,G69531,G69532,G69533,G69534,G69535,G69536,G69537,G69538,G69539,G69540,
       G69541,G69542,G69543,G69544,G69545,G69546,G69547,G69548,G69549,G69550,G69551,G69552,G69553,G69554,G69555,G69556,G69557,G69558,G69559,G69560,
       G69561,G69562,G69563,G69564,G69565,G69566,G69567,G69568,G69569,G69570,G69571,G69572,G69573,G69574,G69575,G69576,G69577,G69578,G69579,G69580,
       G69581,G69582,G69583,G69584,G69585,G69586,G69587,G69588,G69589,G69590,G69591,G69592,G69593,G69594,G69595,G69596,G69597,G69598,G69599,G69600,
       G69601,G69602,G69603,G69604,G69605,G69606,G69607,G69608,G69609,G69610,G69611,G69612,G69613,G69614,G69615,G69616,G69617,G69618,G69619,G69620,
       G69621,G69622,G69623,G69624,G69625,G69626,G69627,G69628,G69629,G69630,G69631,G69632,G69633,G69634,G69635,G69636,G69637,G69638,G69639,G69640,
       G69641,G69642,G69643,G69644,G69645,G69646,G69647,G69648,G69649,G69650,G69651,G69652,G69653,G69654,G69655,G69656,G69657,G69658,G69659,G69660,
       G69661,G69662,G69663,G69664,G69665,G69666,G69667,G69668,G69669,G69670,G69671,G69672,G69673,G69674,G69675,G69676,G69677,G69678,G69679,G69680,
       G69681,G69682,G69683,G69684,G69685,G69686,G69687,G69688,G69689,G69690,G69691,G69692,G69693,G69694,G69695,G69696,G69697,G69698,G69699,G69700,
       G69701,G69702,G69703,G69704,G69705,G69706,G69707,G69708,G69709,G69710,G69711,G69712,G69713,G69714,G69715,G69716,G69717,G69718,G69719,G69720,
       G69721,G69722,G69723,G69724,G69725,G69726,G69727,G69728,G69729,G69730,G69731,G69732,G69733,G69734,G69735,G69736,G69737,G69738,G69739,G69740,
       G69741,G69742,G69743,G69744,G69745,G69746,G69747,G69748,G69749,G69750,G69751,G69752,G69753,G69754,G69755,G69756,G69757,G69758,G69759,G69760,
       G69761,G69762,G69763,G69764,G69765,G69766,G69767,G69768,G69769,G69770,G69771,G69772,G69773,G69774,G69775,G69776,G69777,G69778,G69779,G69780,
       G69781,G69782,G69783,G69784,G69785,G69786,G69787,G69788,G69789,G69790,G69791,G69792,G69793,G69794,G69795,G69796,G69797,G69798,G69799,G69800,
       G69801,G69802,G69803,G69804,G69805,G69806,G69807,G69808,G69809,G69810,G69811,G69812,G69813,G69814,G69815,G69816,G69817,G69818,G69819,G69820,
       G69821,G69822,G69823,G69824,G69825,G69826,G69827,G69828,G69829,G69830,G69831,G69832,G69833,G69834,G69835,G69836,G69837,G69838,G69839,G69840,
       G69841,G69842,G69843,G69844,G69845,G69846,G69847,G69848,G69849,G69850,G69851,G69852,G69853,G69854,G69855,G69856,G69857,G69858,G69859,G69860,
       G69861,G69862,G69863,G69864,G69865,G69866,G69867,G69868,G69869,G69870,G69871,G69872,G69873,G69874,G69875,G69876,G69877,G69878,G69879,G69880,
       G69881,G69882,G69883,G69884,G69885,G69886,G69887,G69888,G69889,G69890,G69891,G69892,G69893,G69894,G69895,G69896,G69897,G69898,G69899,G69900,
       G69901,G69902,G69903,G69904,G69905,G69906,G69907,G69908,G69909,G69910,G69911,G69912,G69913,G69914,G69915,G69916,G69917,G69918,G69919,G69920,
       G69921,G69922,G69923,G69924,G69925,G69926,G69927,G69928,G69929,G69930,G69931,G69932,G69933,G69934,G69935,G69936,G69937,G69938,G69939,G69940,
       G69941,G69942,G69943,G69944,G69945,G69946,G69947,G69948,G69949,G69950,G69951,G69952,G69953,G69954,G69955,G69956,G69957,G69958,G69959,G69960,
       G69961,G69962,G69963,G69964,G69965,G69966,G69967,G69968,G69969,G69970,G69971,G69972,G69973,G69974,G69975,G69976,G69977,G69978,G69979,G69980,
       G69981,G69982,G69983,G69984,G69985,G69986,G69987,G69988,G69989,G69990,G69991,G69992,G69993,G69994,G69995,G69996,G69997,G69998,G69999,G70000,
       G70001,G70002,G70003,G70004,G70005,G70006,G70007,G70008,G70009,G70010,G70011,G70012,G70013,G70014,G70015,G70016,G70017,G70018,G70019,G70020,
       G70021,G70022,G70023,G70024,G70025,G70026,G70027,G70028,G70029,G70030,G70031,G70032,G70033,G70034,G70035,G70036,G70037,G70038,G70039,G70040,
       G70041,G70042,G70043,G70044,G70045,G70046,G70047,G70048,G70049,G70050,G70051,G70052,G70053,G70054,G70055,G70056,G70057,G70058,G70059,G70060,
       G70061,G70062,G70063,G70064,G70065,G70066,G70067,G70068,G70069,G70070,G70071,G70072,G70073,G70074,G70075,G70076,G70077,G70078,G70079,G70080,
       G70081,G70082,G70083,G70084,G70085,G70086,G70087,G70088,G70089,G70090,G70091,G70092,G70093,G70094,G70095,G70096,G70097,G70098,G70099,G70100,
       G70101,G70102,G70103,G70104,G70105,G70106,G70107,G70108,G70109,G70110,G70111,G70112,G70113,G70114,G70115,G70116,G70117,G70118,G70119,G70120,
       G70121,G70122,G70123,G70124,G70125,G70126,G70127,G70128,G70129,G70130,G70131,G70132,G70133,G70134,G70135,G70136,G70137,G70138,G70139,G70140,
       G70141,G70142,G70143,G70144,G70145,G70146,G70147,G70148,G70149,G70150,G70151,G70152,G70153,G70154,G70155,G70156,G70157,G70158,G70159,G70160,
       G70161,G70162,G70163,G70164,G70165,G70166,G70167,G70168,G70169,G70170,G70171,G70172,G70173,G70174,G70175,G70176,G70177,G70178,G70179,G70180,
       G70181,G70182,G70183,G70184,G70185,G70186,G70187,G70188,G70189,G70190,G70191,G70192,G70193,G70194,G70195,G70196,G70197,G70198,G70199,G70200,
       G70201,G70202,G70203,G70204,G70205,G70206,G70207,G70208,G70209,G70210,G70211,G70212,G70213,G70214,G70215,G70216,G70217,G70218,G70219,G70220,
       G70221,G70222,G70223,G70224,G70225,G70226,G70227,G70228,G70229,G70230,G70231,G70232,G70233,G70234,G70235,G70236,G70237,G70238,G70239,G70240,
       G70241,G70242,G70243,G70244,G70245,G70246,G70247,G70248,G70249,G70250,G70251,G70252,G70253,G70254,G70255,G70256,G70257,G70258,G70259,G70260,
       G70261,G70262,G70263,G70264,G70265,G70266,G70267,G70268,G70269,G70270,G70271,G70272,G70273,G70274,G70275,G70276,G70277,G70278,G70279,G70280,
       G70281,G70282,G70283,G70284,G70285,G70286,G70287,G70288,G70289,G70290,G70291,G70292,G70293,G70294,G70295,G70296,G70297,G70298,G70299,G70300,
       G70301,G70302,G70303,G70304,G70305,G70306,G70307,G70308,G70309,G70310,G70311,G70312,G70313,G70314,G70315,G70316,G70317,G70318,G70319,G70320,
       G70321,G70322,G70323,G70324,G70325,G70326,G70327,G70328,G70329,G70330,G70331,G70332,G70333,G70334,G70335,G70336,G70337,G70338,G70339,G70340,
       G70341,G70342,G70343,G70344,G70345,G70346,G70347,G70348,G70349,G70350,G70351,G70352,G70353,G70354,G70355,G70356,G70357,G70358,G70359,G70360,
       G70361,G70362,G70363,G70364,G70365,G70366,G70367,G70368,G70369,G70370,G70371,G70372,G70373,G70374,G70375,G70376,G70377,G70378,G70379,G70380,
       G70381,G70382,G70383,G70384,G70385,G70386,G70387,G70388,G70389,G70390,G70391,G70392,G70393,G70394,G70395,G70396,G70397,G70398,G70399,G70400,
       G70401,G70402,G70403,G70404,G70405,G70406,G70407,G70408,G70409,G70410,G70411,G70412,G70413,G70414,G70415,G70416,G70417,G70418,G70419,G70420,
       G70421,G70422,G70423,G70424,G70425,G70426,G70427,G70428,G70429,G70430,G70431,G70432,G70433,G70434,G70435,G70436,G70437,G70438,G70439,G70440,
       G70441,G70442,G70443,G70444,G70445,G70446,G70447,G70448,G70449,G70450,G70451,G70452,G70453,G70454,G70455,G70456,G70457,G70458,G70459,G70460,
       G70461,G70462,G70463,G70464,G70465,G70466,G70467,G70468,G70469,G70470,G70471,G70472,G70473,G70474,G70475,G70476,G70477,G70478,G70479,G70480,
       G70481,G70482,G70483,G70484,G70485,G70486,G70487,G70488,G70489,G70490,G70491,G70492,G70493,G70494,G70495,G70496,G70497,G70498,G70499,G70500,
       G70501,G70502,G70503,G70504,G70505,G70506,G70507,G70508,G70509,G70510,G70511,G70512,G70513,G70514,G70515,G70516,G70517,G70518,G70519,G70520,
       G70521,G70522,G70523,G70524,G70525,G70526,G70527,G70528,G70529,G70530,G70531,G70532,G70533,G70534,G70535,G70536,G70537,G70538,G70539,G70540,
       G70541,G70542,G70543,G70544,G70545,G70546,G70547,G70548,G70549,G70550,G70551,G70552,G70553,G70554,G70555,G70556,G70557,G70558,G70559,G70560,
       G70561,G70562,G70563,G70564,G70565,G70566,G70567,G70568,G70569,G70570,G70571,G70572,G70573,G70574,G70575,G70576,G70577,G70578,G70579,G70580,
       G70581,G70582,G70583,G70584,G70585,G70586,G70587,G70588,G70589,G70590,G70591,G70592,G70593,G70594,G70595,G70596,G70597,G70598,G70599,G70600,
       G70601,G70602,G70603,G70604,G70605,G70606,G70607,G70608,G70609,G70610,G70611,G70612,G70613,G70614,G70615,G70616,G70617,G70618,G70619,G70620,
       G70621,G70622,G70623,G70624,G70625,G70626,G70627,G70628,G70629,G70630,G70631,G70632,G70633,G70634,G70635,G70636,G70637,G70638,G70639,G70640,
       G70641,G70642,G70643,G70644,G70645,G70646,G70647,G70648,G70649,G70650,G70651,G70652,G70653,G70654,G70655,G70656,G70657,G70658,G70659,G70660,
       G70661,G70662,G70663,G70664,G70665,G70666,G70667,G70668,G70669,G70670,G70671,G70672,G70673,G70674,G70675,G70676,G70677,G70678,G70679,G70680,
       G70681,G70682,G70683,G70684,G70685,G70686,G70687,G70688,G70689,G70690,G70691,G70692,G70693,G70694,G70695,G70696,G70697,G70698,G70699,G70700,
       G70701,G70702,G70703,G70704,G70705,G70706,G70707,G70708,G70709,G70710,G70711,G70712,G70713,G70714,G70715,G70716,G70717,G70718,G70719,G70720,
       G70721,G70722,G70723,G70724,G70725,G70726,G70727,G70728,G70729,G70730,G70731,G70732,G70733,G70734,G70735,G70736,G70737,G70738,G70739,G70740,
       G70741,G70742,G70743,G70744,G70745,G70746,G70747,G70748,G70749,G70750,G70751,G70752,G70753,G70754,G70755,G70756,G70757,G70758,G70759,G70760,
       G70761,G70762,G70763,G70764,G70765,G70766,G70767,G70768,G70769,G70770,G70771,G70772,G70773,G70774,G70775,G70776,G70777,G70778,G70779,G70780,
       G70781,G70782,G70783,G70784,G70785,G70786,G70787,G70788,G70789,G70790,G70791,G70792,G70793,G70794,G70795,G70796,G70797,G70798,G70799,G70800,
       G70801,G70802,G70803,G70804,G70805,G70806,G70807,G70808,G70809,G70810,G70811,G70812,G70813,G70814,G70815,G70816,G70817,G70818,G70819,G70820,
       G70821,G70822,G70823,G70824,G70825,G70826,G70827,G70828,G70829,G70830,G70831,G70832,G70833,G70834,G70835,G70836,G70837,G70838,G70839,G70840,
       G70841,G70842,G70843,G70844,G70845,G70846,G70847,G70848,G70849,G70850,G70851,G70852,G70853,G70854,G70855,G70856,G70857,G70858,G70859,G70860,
       G70861,G70862,G70863,G70864,G70865,G70866,G70867,G70868,G70869,G70870,G70871,G70872,G70873,G70874,G70875,G70876,G70877,G70878,G70879,G70880,
       G70881,G70882,G70883,G70884,G70885,G70886,G70887,G70888,G70889,G70890,G70891,G70892,G70893,G70894,G70895,G70896,G70897,G70898,G70899,G70900,
       G70901,G70902,G70903,G70904,G70905,G70906,G70907,G70908,G70909,G70910,G70911,G70912,G70913,G70914,G70915,G70916,G70917,G70918,G70919,G70920,
       G70921,G70922,G70923,G70924,G70925,G70926,G70927,G70928,G70929,G70930,G70931,G70932,G70933,G70934,G70935,G70936,G70937,G70938,G70939,G70940,
       G70941,G70942,G70943,G70944,G70945,G70946,G70947,G70948,G70949,G70950,G70951,G70952,G70953,G70954,G70955,G70956,G70957,G70958,G70959,G70960,
       G70961,G70962,G70963,G70964,G70965,G70966,G70967,G70968,G70969,G70970,G70971,G70972,G70973,G70974,G70975,G70976,G70977,G70978,G70979,G70980,
       G70981,G70982,G70983,G70984,G70985,G70986,G70987,G70988,G70989,G70990,G70991,G70992,G70993,G70994,G70995,G70996,G70997,G70998,G70999,G71000,
       G71001,G71002,G71003,G71004,G71005,G71006,G71007,G71008,G71009,G71010,G71011,G71012,G71013,G71014,G71015,G71016,G71017,G71018,G71019,G71020,
       G71021,G71022,G71023,G71024,G71025,G71026,G71027,G71028,G71029,G71030,G71031,G71032,G71033,G71034,G71035,G71036,G71037,G71038,G71039,G71040,
       G71041,G71042,G71043,G71044,G71045,G71046,G71047,G71048,G71049,G71050,G71051,G71052,G71053,G71054,G71055,G71056,G71057,G71058,G71059,G71060,
       G71061,G71062,G71063,G71064,G71065,G71066,G71067,G71068,G71069,G71070,G71071,G71072,G71073,G71074,G71075,G71076,G71077,G71078,G71079,G71080,
       G71081,G71082,G71083,G71084,G71085,G71086,G71087,G71088,G71089,G71090,G71091,G71092,G71093,G71094,G71095,G71096,G71097,G71098,G71099,G71100,
       G71101,G71102,G71103,G71104,G71105,G71106,G71107,G71108,G71109,G71110,G71111,G71112,G71113,G71114,G71115,G71116,G71117,G71118,G71119,G71120,
       G71121,G71122,G71123,G71124,G71125,G71126,G71127,G71128,G71129,G71130,G71131,G71132,G71133,G71134,G71135,G71136,G71137,G71138,G71139,G71140,
       G71141,G71142,G71143,G71144,G71145,G71146,G71147,G71148,G71149,G71150,G71151,G71152,G71153,G71154,G71155,G71156,G71157,G71158,G71159,G71160,
       G71161,G71162,G71163,G71164,G71165,G71166,G71167,G71168,G71169,G71170,G71171,G71172,G71173,G71174,G71175,G71176,G71177,G71178,G71179,G71180,
       G71181,G71182,G71183,G71184,G71185,G71186,G71187,G71188,G71189,G71190,G71191,G71192,G71193,G71194,G71195,G71196,G71197,G71198,G71199,G71200,
       G71201,G71202,G71203,G71204,G71205,G71206,G71207,G71208,G71209,G71210,G71211,G71212,G71213,G71214,G71215,G71216,G71217,G71218,G71219,G71220,
       G71221,G71222,G71223,G71224,G71225,G71226,G71227,G71228,G71229,G71230,G71231,G71232,G71233,G71234,G71235,G71236,G71237,G71238,G71239,G71240,
       G71241,G71242,G71243,G71244,G71245,G71246,G71247,G71248,G71249,G71250,G71251,G71252,G71253,G71254,G71255,G71256,G71257,G71258,G71259,G71260,
       G71261,G71262,G71263,G71264,G71265,G71266,G71267,G71268,G71269,G71270,G71271,G71272,G71273,G71274,G71275,G71276,G71277,G71278,G71279,G71280,
       G71281,G71282,G71283,G71284,G71285,G71286,G71287,G71288,G71289,G71290,G71291,G71292,G71293,G71294,G71295,G71296,G71297,G71298,G71299,G71300,
       G71301,G71302,G71303,G71304,G71305,G71306,G71307,G71308,G71309,G71310,G71311,G71312,G71313,G71314,G71315,G71316,G71317,G71318,G71319,G71320,
       G71321,G71322,G71323,G71324,G71325,G71326,G71327,G71328,G71329,G71330,G71331,G71332,G71333,G71334,G71335,G71336,G71337,G71338,G71339,G71340,
       G71341,G71342,G71343,G71344,G71345,G71346,G71347,G71348,G71349,G71350,G71351,G71352,G71353,G71354,G71355,G71356,G71357,G71358,G71359,G71360,
       G71361,G71362,G71363,G71364,G71365,G71366,G71367,G71368,G71369,G71370,G71371,G71372,G71373,G71374,G71375,G71376,G71377,G71378,G71379,G71380,
       G71381,G71382,G71383,G71384,G71385,G71386,G71387,G71388,G71389,G71390,G71391,G71392,G71393,G71394,G71395,G71396,G71397,G71398,G71399,G71400,
       G71401,G71402,G71403,G71404,G71405,G71406,G71407,G71408,G71409,G71410,G71411,G71412,G71413,G71414,G71415,G71416,G71417,G71418,G71419,G71420,
       G71421,G71422,G71423,G71424,G71425,G71426,G71427,G71428,G71429,G71430,G71431,G71432,G71433,G71434,G71435,G71436,G71437,G71438,G71439,G71440,
       G71441,G71442,G71443,G71444,G71445,G71446,G71447,G71448,G71449,G71450,G71451,G71452,G71453,G71454,G71455,G71456,G71457,G71458,G71459,G71460,
       G71461,G71462,G71463,G71464,G71465,G71466,G71467,G71468,G71469,G71470,G71471,G71472,G71473,G71474,G71475,G71476,G71477,G71478,G71479,G71480,
       G71481,G71482,G71483,G71484,G71485,G71486,G71487,G71488,G71489,G71490,G71491,G71492,G71493,G71494,G71495,G71496,G71497,G71498,G71499,G71500,
       G71501,G71502,G71503,G71504,G71505,G71506,G71507,G71508,G71509,G71510,G71511,G71512,G71513,G71514,G71515,G71516,G71517,G71518,G71519,G71520,
       G71521,G71522,G71523,G71524,G71525,G71526,G71527,G71528,G71529,G71530,G71531,G71532,G71533,G71534,G71535,G71536,G71537,G71538,G71539,G71540,
       G71541,G71542,G71543,G71544,G71545,G71546,G71547,G71548,G71549,G71550,G71551,G71552,G71553,G71554,G71555,G71556,G71557,G71558,G71559,G71560,
       G71561,G71562,G71563,G71564,G71565,G71566,G71567,G71568,G71569,G71570,G71571,G71572,G71573,G71574,G71575,G71576,G71577,G71578,G71579,G71580,
       G71581,G71582,G71583,G71584,G71585,G71586,G71587,G71588,G71589,G71590,G71591,G71592,G71593,G71594,G71595,G71596,G71597,G71598,G71599,G71600,
       G71601,G71602,G71603,G71604,G71605,G71606,G71607,G71608,G71609,G71610,G71611,G71612,G71613,G71614,G71615,G71616,G71617,G71618,G71619,G71620,
       G71621,G71622,G71623,G71624,G71625,G71626,G71627,G71628,G71629,G71630,G71631,G71632,G71633,G71634,G71635,G71636,G71637,G71638,G71639,G71640,
       G71641,G71642,G71643,G71644,G71645,G71646,G71647,G71648,G71649,G71650,G71651,G71652,G71653,G71654,G71655,G71656,G71657,G71658,G71659,G71660,
       G71661,G71662,G71663,G71664,G71665,G71666,G71667,G71668,G71669,G71670,G71671,G71672,G71673,G71674,G71675,G71676,G71677,G71678,G71679,G71680,
       G71681,G71682,G71683,G71684,G71685,G71686,G71687,G71688,G71689,G71690,G71691,G71692,G71693,G71694,G71695,G71696,G71697,G71698,G71699,G71700,
       G71701,G71702,G71703,G71704,G71705,G71706,G71707,G71708,G71709,G71710,G71711,G71712,G71713,G71714,G71715,G71716,G71717,G71718,G71719,G71720,
       G71721,G71722,G71723,G71724,G71725,G71726,G71727,G71728,G71729,G71730,G71731,G71732,G71733,G71734,G71735,G71736,G71737,G71738,G71739,G71740,
       G71741,G71742,G71743,G71744,G71745,G71746,G71747,G71748,G71749,G71750,G71751,G71752,G71753,G71754,G71755,G71756,G71757,G71758,G71759,G71760,
       G71761,G71762,G71763,G71764,G71765,G71766,G71767,G71768,G71769,G71770,G71771,G71772,G71773,G71774,G71775,G71776,G71777,G71778,G71779,G71780,
       G71781,G71782,G71783,G71784,G71785,G71786,G71787,G71788,G71789,G71790,G71791,G71792,G71793,G71794,G71795,G71796,G71797,G71798,G71799,G71800,
       G71801,G71802,G71803,G71804,G71805,G71806,G71807,G71808,G71809,G71810,G71811,G71812,G71813,G71814,G71815,G71816,G71817,G71818,G71819,G71820,
       G71821,G71822,G71823,G71824,G71825,G71826,G71827,G71828,G71829,G71830,G71831,G71832,G71833,G71834,G71835,G71836,G71837,G71838,G71839,G71840,
       G71841,G71842,G71843,G71844,G71845,G71846,G71847,G71848,G71849,G71850,G71851,G71852,G71853,G71854,G71855,G71856,G71857,G71858,G71859,G71860,
       G71861,G71862,G71863,G71864,G71865,G71866,G71867,G71868,G71869,G71870,G71871,G71872,G71873,G71874,G71875,G71876,G71877,G71878,G71879,G71880,
       G71881,G71882,G71883,G71884,G71885,G71886,G71887,G71888,G71889,G71890,G71891,G71892,G71893,G71894,G71895,G71896,G71897,G71898,G71899,G71900,
       G71901,G71902,G71903,G71904,G71905,G71906,G71907,G71908,G71909,G71910,G71911,G71912,G71913,G71914,G71915,G71916,G71917,G71918,G71919,G71920,
       G71921,G71922,G71923,G71924,G71925,G71926,G71927,G71928,G71929,G71930,G71931,G71932,G71933,G71934,G71935,G71936,G71937,G71938,G71939,G71940,
       G71941,G71942,G71943,G71944,G71945,G71946,G71947,G71948,G71949,G71950,G71951,G71952,G71953,G71954,G71955,G71956,G71957,G71958,G71959,G71960,
       G71961,G71962,G71963,G71964,G71965,G71966,G71967,G71968,G71969,G71970,G71971,G71972,G71973,G71974,G71975,G71976,G71977,G71978,G71979,G71980,
       G71981,G71982,G71983,G71984,G71985,G71986,G71987,G71988,G71989,G71990,G71991,G71992,G71993,G71994,G71995,G71996,G71997,G71998,G71999,G72000,
       G72001,G72002,G72003,G72004,G72005,G72006,G72007,G72008,G72009,G72010,G72011,G72012,G72013,G72014,G72015,G72016,G72017,G72018,G72019,G72020,
       G72021,G72022,G72023,G72024,G72025,G72026,G72027,G72028,G72029,G72030,G72031,G72032,G72033,G72034,G72035,G72036,G72037,G72038,G72039,G72040,
       G72041,G72042,G72043,G72044,G72045,G72046,G72047,G72048,G72049,G72050,G72051,G72052,G72053,G72054,G72055,G72056,G72057,G72058,G72059,G72060,
       G72061,G72062,G72063,G72064,G72065,G72066,G72067,G72068,G72069,G72070,G72071,G72072,G72073,G72074,G72075,G72076,G72077,G72078,G72079,G72080,
       G72081,G72082,G72083,G72084,G72085,G72086,G72087,G72088,G72089,G72090,G72091,G72092,G72093,G72094,G72095,G72096,G72097,G72098,G72099,G72100,
       G72101,G72102,G72103,G72104,G72105,G72106,G72107,G72108,G72109,G72110,G72111,G72112,G72113,G72114,G72115,G72116,G72117,G72118,G72119,G72120,
       G72121,G72122,G72123,G72124,G72125,G72126,G72127,G72128,G72129,G72130,G72131,G72132,G72133,G72134,G72135,G72136,G72137,G72138,G72139,G72140,
       G72141,G72142,G72143,G72144,G72145,G72146,G72147,G72148,G72149,G72150,G72151,G72152,G72153,G72154,G72155,G72156,G72157,G72158,G72159,G72160,
       G72161,G72162,G72163,G72164,G72165,G72166,G72167,G72168,G72169,G72170,G72171,G72172,G72173,G72174,G72175,G72176,G72177,G72178,G72179,G72180,
       G72181,G72182,G72183,G72184,G72185,G72186,G72187,G72188,G72189,G72190,G72191,G72192,G72193,G72194,G72195,G72196,G72197,G72198,G72199,G72200,
       G72201,G72202,G72203,G72204,G72205,G72206,G72207,G72208,G72209,G72210,G72211,G72212,G72213,G72214,G72215,G72216,G72217,G72218,G72219,G72220,
       G72221,G72222,G72223,G72224,G72225,G72226,G72227,G72228,G72229,G72230,G72231,G72232,G72233,G72234,G72235,G72236,G72237,G72238,G72239,G72240,
       G72241,G72242,G72243,G72244,G72245,G72246,G72247,G72248,G72249,G72250,G72251,G72252,G72253,G72254,G72255,G72256,G72257,G72258,G72259,G72260,
       G72261,G72262,G72263,G72264,G72265,G72266,G72267,G72268,G72269,G72270,G72271,G72272,G72273,G72274,G72275,G72276,G72277,G72278,G72279,G72280,
       G72281,G72282,G72283,G72284,G72285,G72286,G72287,G72288,G72289,G72290,G72291,G72292,G72293,G72294,G72295,G72296,G72297,G72298,G72299,G72300,
       G72301,G72302,G72303,G72304,G72305,G72306,G72307,G72308,G72309,G72310,G72311,G72312,G72313,G72314,G72315,G72316,G72317,G72318,G72319,G72320,
       G72321,G72322,G72323,G72324,G72325,G72326,G72327,G72328,G72329,G72330,G72331,G72332,G72333,G72334,G72335,G72336,G72337,G72338,G72339,G72340,
       G72341,G72342,G72343,G72344,G72345,G72346,G72347,G72348,G72349,G72350,G72351,G72352,G72353,G72354,G72355,G72356,G72357,G72358,G72359,G72360,
       G72361,G72362,G72363,G72364,G72365,G72366,G72367,G72368,G72369,G72370,G72371,G72372,G72373,G72374,G72375,G72376,G72377,G72378,G72379,G72380,
       G72381,G72382,G72383,G72384,G72385,G72386,G72387,G72388,G72389,G72390,G72391,G72392,G72393,G72394,G72395,G72396,G72397,G72398,G72399,G72400,
       G72401,G72402,G72403,G72404,G72405,G72406,G72407,G72408,G72409,G72410,G72411,G72412,G72413,G72414,G72415,G72416,G72417,G72418,G72419,G72420,
       G72421,G72422,G72423,G72424,G72425,G72426,G72427,G72428,G72429,G72430,G72431,G72432,G72433,G72434,G72435,G72436,G72437,G72438,G72439,G72440,
       G72441,G72442,G72443,G72444,G72445,G72446,G72447,G72448,G72449,G72450,G72451,G72452,G72453,G72454,G72455,G72456,G72457,G72458,G72459,G72460,
       G72461,G72462,G72463,G72464,G72465,G72466,G72467,G72468,G72469,G72470,G72471,G72472,G72473,G72474,G72475,G72476,G72477,G72478,G72479,G72480,
       G72481,G72482,G72483,G72484,G72485,G72486,G72487,G72488,G72489,G72490,G72491,G72492,G72493,G72494,G72495,G72496,G72497,G72498,G72499,G72500,
       G72501,G72502,G72503,G72504,G72505,G72506,G72507,G72508,G72509,G72510,G72511,G72512,G72513,G72514,G72515,G72516,G72517,G72518,G72519,G72520,
       G72521,G72522,G72523,G72524,G72525,G72526,G72527,G72528,G72529,G72530,G72531,G72532,G72533,G72534,G72535,G72536,G72537,G72538,G72539,G72540,
       G72541,G72542,G72543,G72544,G72545,G72546,G72547,G72548,G72549,G72550,G72551,G72552,G72553,G72554,G72555,G72556,G72557,G72558,G72559,G72560,
       G72561,G72562,G72563,G72564,G72565,G72566,G72567,G72568,G72569,G72570,G72571,G72572,G72573,G72574,G72575,G72576,G72577,G72578,G72579,G72580,
       G72581,G72582,G72583,G72584,G72585,G72586,G72587,G72588,G72589,G72590,G72591,G72592,G72593,G72594,G72595,G72596,G72597,G72598,G72599,G72600,
       G72601,G72602,G72603,G72604,G72605,G72606,G72607,G72608,G72609,G72610,G72611,G72612,G72613,G72614,G72615,G72616,G72617,G72618,G72619,G72620,
       G72621,G72622,G72623,G72624,G72625,G72626,G72627,G72628,G72629,G72630,G72631,G72632,G72633,G72634,G72635,G72636,G72637,G72638,G72639,G72640,
       G72641,G72642,G72643,G72644,G72645,G72646,G72647,G72648,G72649,G72650,G72651,G72652,G72653,G72654,G72655,G72656,G72657,G72658,G72659,G72660,
       G72661,G72662,G72663,G72664,G72665,G72666,G72667,G72668,G72669,G72670,G72671,G72672,G72673,G72674,G72675,G72676,G72677,G72678,G72679,G72680,
       G72681,G72682,G72683,G72684,G72685,G72686,G72687,G72688,G72689,G72690,G72691,G72692,G72693,G72694,G72695,G72696,G72697,G72698,G72699,G72700,
       G72701,G72702,G72703,G72704,G72705,G72706,G72707,G72708,G72709,G72710,G72711,G72712,G72713,G72714,G72715,G72716,G72717,G72718,G72719,G72720,
       G72721,G72722,G72723,G72724,G72725,G72726,G72727,G72728,G72729,G72730,G72731,G72732,G72733,G72734,G72735,G72736,G72737,G72738,G72739,G72740,
       G72741,G72742,G72743,G72744,G72745,G72746,G72747,G72748,G72749,G72750,G72751,G72752,G72753,G72754,G72755,G72756,G72757,G72758,G72759,G72760,
       G72761,G72762,G72763,G72764,G72765,G72766,G72767,G72768,G72769,G72770,G72771,G72772,G72773,G72774,G72775,G72776,G72777,G72778,G72779,G72780,
       G72781,G72782,G72783,G72784,G72785,G72786,G72787,G72788,G72789,G72790,G72791,G72792,G72793,G72794,G72795,G72796,G72797,G72798,G72799,G72800,
       G72801,G72802,G72803,G72804,G72805,G72806,G72807,G72808,G72809,G72810,G72811,G72812,G72813,G72814,G72815,G72816,G72817,G72818,G72819,G72820,
       G72821,G72822,G72823,G72824,G72825,G72826,G72827,G72828,G72829,G72830,G72831,G72832,G72833,G72834,G72835,G72836,G72837,G72838,G72839,G72840,
       G72841,G72842,G72843,G72844,G72845,G72846,G72847,G72848,G72849,G72850,G72851,G72852,G72853,G72854,G72855,G72856,G72857,G72858,G72859,G72860,
       G72861,G72862,G72863,G72864,G72865,G72866,G72867,G72868,G72869,G72870,G72871,G72872,G72873,G72874,G72875,G72876,G72877,G72878,G72879,G72880,
       G72881,G72882,G72883,G72884,G72885,G72886,G72887,G72888,G72889,G72890,G72891,G72892,G72893,G72894,G72895,G72896,G72897,G72898,G72899,G72900,
       G72901,G72902,G72903,G72904,G72905,G72906,G72907,G72908,G72909,G72910,G72911,G72912,G72913,G72914,G72915,G72916,G72917,G72918,G72919,G72920,
       G72921,G72922,G72923,G72924,G72925,G72926,G72927,G72928,G72929,G72930,G72931,G72932,G72933,G72934,G72935,G72936,G72937,G72938,G72939,G72940,
       G72941,G72942,G72943,G72944,G72945,G72946,G72947,G72948,G72949,G72950,G72951,G72952,G72953,G72954,G72955,G72956,G72957,G72958,G72959,G72960,
       G72961,G72962,G72963,G72964,G72965,G72966,G72967,G72968,G72969,G72970,G72971,G72972,G72973,G72974,G72975,G72976,G72977,G72978,G72979,G72980,
       G72981,G72982,G72983,G72984,G72985,G72986,G72987,G72988,G72989,G72990,G72991,G72992,G72993,G72994,G72995,G72996,G72997,G72998,G72999,G73000,
       G73001,G73002,G73003,G73004,G73005,G73006,G73007,G73008,G73009,G73010,G73011,G73012,G73013,G73014,G73015,G73016,G73017,G73018,G73019,G73020,
       G73021,G73022,G73023,G73024,G73025,G73026,G73027,G73028,G73029,G73030,G73031,G73032,G73033,G73034,G73035,G73036,G73037,G73038,G73039,G73040,
       G73041,G73042,G73043,G73044,G73045,G73046,G73047,G73048,G73049,G73050,G73051,G73052,G73053,G73054,G73055,G73056,G73057,G73058,G73059,G73060,
       G73061,G73062,G73063,G73064,G73065,G73066,G73067,G73068,G73069,G73070,G73071,G73072,G73073,G73074,G73075,G73076,G73077,G73078,G73079,G73080,
       G73081,G73082,G73083,G73084,G73085,G73086,G73087,G73088,G73089,G73090,G73091,G73092,G73093,G73094,G73095,G73096,G73097,G73098,G73099,G73100,
       G73101,G73102,G73103,G73104,G73105,G73106,G73107,G73108,G73109,G73110,G73111,G73112,G73113,G73114,G73115,G73116,G73117,G73118,G73119,G73120,
       G73121,G73122,G73123,G73124,G73125,G73126,G73127,G73128,G73129,G73130,G73131,G73132,G73133,G73134,G73135,G73136,G73137,G73138,G73139,G73140,
       G73141,G73142,G73143,G73144,G73145,G73146,G73147,G73148,G73149,G73150,G73151,G73152,G73153,G73154,G73155,G73156,G73157,G73158,G73159,G73160,
       G73161,G73162,G73163,G73164,G73165,G73166,G73167,G73168,G73169,G73170,G73171,G73172,G73173,G73174,G73175,G73176,G73177,G73178,G73179,G73180,
       G73181,G73182,G73183,G73184,G73185,G73186,G73187,G73188,G73189,G73190,G73191,G73192,G73193,G73194,G73195,G73196,G73197,G73198,G73199,G73200,
       G73201,G73202,G73203,G73204,G73205,G73206,G73207,G73208,G73209,G73210,G73211,G73212,G73213,G73214,G73215,G73216,G73217,G73218,G73219,G73220,
       G73221,G73222,G73223,G73224,G73225,G73226,G73227,G73228,G73229,G73230,G73231,G73232,G73233,G73234,G73235,G73236,G73237,G73238,G73239,G73240,
       G73241,G73242,G73243,G73244,G73245,G73246,G73247,G73248,G73249,G73250,G73251,G73252,G73253,G73254,G73255,G73256,G73257,G73258,G73259,G73260,
       G73261,G73262,G73263,G73264,G73265,G73266,G73267,G73268,G73269,G73270,G73271,G73272,G73273,G73274,G73275,G73276,G73277,G73278,G73279,G73280,
       G73281,G73282,G73283,G73284,G73285,G73286,G73287,G73288,G73289,G73290,G73291,G73292,G73293,G73294,G73295,G73296,G73297,G73298,G73299,G73300,
       G73301,G73302,G73303,G73304,G73305,G73306,G73307,G73308,G73309,G73310,G73311,G73312,G73313,G73314,G73315,G73316,G73317,G73318,G73319,G73320,
       G73321,G73322,G73323,G73324,G73325,G73326,G73327,G73328,G73329,G73330,G73331,G73332,G73333,G73334,G73335,G73336,G73337,G73338,G73339,G73340,
       G73341,G73342,G73343,G73344,G73345,G73346,G73347,G73348,G73349,G73350,G73351,G73352,G73353,G73354,G73355,G73356,G73357,G73358,G73359,G73360,
       G73361,G73362,G73363,G73364,G73365,G73366,G73367,G73368,G73369,G73370,G73371,G73372,G73373,G73374,G73375,G73376,G73377,G73378,G73379,G73380,
       G73381,G73382,G73383,G73384,G73385,G73386,G73387,G73388,G73389,G73390,G73391,G73392,G73393,G73394,G73395,G73396,G73397,G73398,G73399,G73400,
       G73401,G73402,G73403,G73404,G73405,G73406,G73407,G73408,G73409,G73410,G73411,G73412,G73413,G73414,G73415,G73416,G73417,G73418,G73419,G73420,
       G73421,G73422,G73423,G73424,G73425,G73426,G73427,G73428,G73429,G73430,G73431,G73432,G73433,G73434,G73435,G73436,G73437,G73438,G73439,G73440,
       G73441,G73442,G73443,G73444,G73445,G73446,G73447,G73448,G73449,G73450,G73451,G73452,G73453,G73454,G73455,G73456,G73457,G73458,G73459,G73460,
       G73461,G73462,G73463,G73464,G73465,G73466,G73467,G73468,G73469,G73470,G73471,G73472,G73473,G73474,G73475,G73476,G73477,G73478,G73479,G73480,
       G73481,G73482,G73483,G73484,G73485,G73486,G73487,G73488,G73489,G73490,G73491,G73492,G73493,G73494,G73495,G73496,G73497,G73498,G73499,G73500,
       G73501,G73502,G73503,G73504,G73505,G73506,G73507,G73508,G73509,G73510,G73511,G73512,G73513,G73514,G73515,G73516,G73517,G73518,G73519,G73520,
       G73521,G73522,G73523,G73524,G73525,G73526,G73527,G73528,G73529,G73530,G73531,G73532,G73533,G73534,G73535,G73536,G73537,G73538,G73539,G73540,
       G73541,G73542,G73543,G73544,G73545,G73546,G73547,G73548,G73549,G73550,G73551,G73552,G73553,G73554,G73555,G73556,G73557,G73558,G73559,G73560,
       G73561,G73562,G73563,G73564,G73565,G73566,G73567,G73568,G73569,G73570,G73571,G73572,G73573,G73574,G73575,G73576,G73577,G73578,G73579,G73580,
       G73581,G73582,G73583,G73584,G73585,G73586,G73587,G73588,G73589,G73590,G73591,G73592,G73593,G73594,G73595,G73596,G73597,G73598,G73599,G73600,
       G73601,G73602,G73603,G73604,G73605,G73606,G73607,G73608,G73609,G73610,G73611,G73612,G73613,G73614,G73615,G73616,G73617,G73618,G73619,G73620,
       G73621,G73622,G73623,G73624,G73625,G73626,G73627,G73628,G73629,G73630,G73631,G73632,G73633,G73634,G73635,G73636,G73637,G73638,G73639,G73640,
       G73641,G73642,G73643,G73644,G73645,G73646,G73647,G73648,G73649,G73650,G73651,G73652,G73653,G73654,G73655,G73656,G73657,G73658,G73659,G73660,
       G73661,G73662,G73663,G73664,G73665,G73666,G73667,G73668,G73669,G73670,G73671,G73672,G73673,G73674,G73675,G73676,G73677,G73678,G73679,G73680,
       G73681,G73682,G73683,G73684,G73685,G73686,G73687,G73688,G73689,G73690,G73691,G73692,G73693,G73694,G73695,G73696,G73697,G73698,G73699,G73700,
       G73701,G73702,G73703,G73704,G73705,G73706,G73707,G73708,G73709,G73710,G73711,G73712,G73713,G73714,G73715,G73716,G73717,G73718,G73719,G73720,
       G73721,G73722,G73723,G73724,G73725,G73726,G73727,G73728,G73729,G73730,G73731,G73732,G73733,G73734,G73735,G73736,G73737,G73738,G73739,G73740,
       G73741,G73742,G73743,G73744,G73745,G73746,G73747,G73748,G73749,G73750,G73751,G73752,G73753,G73754,G73755,G73756,G73757,G73758,G73759,G73760,
       G73761,G73762,G73763,G73764,G73765,G73766,G73767,G73768,G73769,G73770,G73771,G73772,G73773,G73774,G73775,G73776,G73777,G73778,G73779,G73780,
       G73781,G73782,G73783,G73784,G73785,G73786,G73787,G73788,G73789,G73790,G73791,G73792,G73793,G73794,G73795,G73796,G73797,G73798,G73799,G73800,
       G73801,G73802,G73803,G73804,G73805,G73806,G73807,G73808,G73809,G73810,G73811,G73812,G73813,G73814,G73815,G73816,G73817,G73818,G73819,G73820,
       G73821,G73822,G73823,G73824,G73825,G73826,G73827,G73828,G73829,G73830,G73831,G73832,G73833,G73834,G73835,G73836,G73837,G73838,G73839,G73840,
       G73841,G73842,G73843,G73844,G73845,G73846,G73847,G73848,G73849,G73850,G73851,G73852,G73853,G73854,G73855,G73856,G73857,G73858,G73859,G73860,
       G73861,G73862,G73863,G73864,G73865,G73866,G73867,G73868,G73869,G73870,G73871,G73872,G73873,G73874,G73875,G73876,G73877,G73878,G73879,G73880,
       G73881,G73882,G73883,G73884,G73885,G73886,G73887,G73888,G73889,G73890,G73891,G73892,G73893,G73894,G73895,G73896,G73897,G73898,G73899,G73900,
       G73901,G73902,G73903,G73904,G73905,G73906,G73907,G73908,G73909,G73910,G73911,G73912,G73913,G73914,G73915,G73916,G73917,G73918,G73919,G73920,
       G73921,G73922,G73923,G73924,G73925,G73926,G73927,G73928,G73929,G73930,G73931,G73932,G73933,G73934,G73935,G73936,G73937,G73938,G73939,G73940,
       G73941,G73942,G73943,G73944,G73945,G73946,G73947,G73948,G73949,G73950,G73951,G73952,G73953,G73954,G73955,G73956,G73957,G73958,G73959,G73960,
       G73961,G73962,G73963,G73964,G73965,G73966,G73967,G73968,G73969,G73970,G73971,G73972,G73973,G73974,G73975,G73976,G73977,G73978,G73979,G73980,
       G73981,G73982,G73983,G73984,G73985,G73986,G73987,G73988,G73989,G73990,G73991,G73992,G73993,G73994,G73995,G73996,G73997,G73998,G73999,G74000,
       G74001,G74002,G74003,G74004,G74005,G74006,G74007,G74008,G74009,G74010,G74011,G74012,G74013,G74014,G74015,G74016,G74017,G74018,G74019,G74020,
       G74021,G74022,G74023,G74024,G74025,G74026,G74027,G74028,G74029,G74030,G74031,G74032,G74033,G74034,G74035,G74036,G74037,G74038,G74039,G74040,
       G74041,G74042,G74043,G74044,G74045,G74046,G74047,G74048,G74049,G74050,G74051,G74052,G74053,G74054,G74055,G74056,G74057,G74058,G74059,G74060,
       G74061,G74062,G74063,G74064,G74065,G74066,G74067,G74068,G74069,G74070,G74071,G74072,G74073,G74074,G74075,G74076,G74077,G74078,G74079,G74080,
       G74081,G74082,G74083,G74084,G74085,G74086,G74087,G74088,G74089,G74090,G74091,G74092,G74093,G74094,G74095,G74096,G74097,G74098,G74099,G74100,
       G74101,G74102,G74103,G74104,G74105,G74106,G74107,G74108,G74109,G74110,G74111,G74112,G74113,G74114,G74115,G74116,G74117,G74118,G74119,G74120,
       G74121,G74122,G74123,G74124,G74125,G74126,G74127,G74128,G74129,G74130,G74131,G74132,G74133,G74134,G74135,G74136,G74137,G74138,G74139,G74140,
       G74141,G74142,G74143,G74144,G74145,G74146,G74147,G74148,G74149,G74150,G74151,G74152,G74153,G74154,G74155,G74156,G74157,G74158,G74159,G74160,
       G74161,G74162,G74163,G74164,G74165,G74166,G74167,G74168,G74169,G74170,G74171,G74172,G74173,G74174,G74175,G74176,G74177,G74178,G74179,G74180,
       G74181,G74182,G74183,G74184,G74185,G74186,G74187,G74188,G74189,G74190,G74191,G74192,G74193,G74194,G74195,G74196,G74197,G74198,G74199,G74200,
       G74201,G74202,G74203,G74204,G74205,G74206,G74207,G74208,G74209,G74210,G74211,G74212,G74213,G74214,G74215,G74216,G74217,G74218,G74219,G74220,
       G74221,G74222,G74223,G74224,G74225,G74226,G74227,G74228,G74229,G74230,G74231,G74232,G74233,G74234,G74235,G74236,G74237,G74238,G74239,G74240,
       G74241,G74242,G74243,G74244,G74245,G74246,G74247,G74248,G74249,G74250,G74251,G74252,G74253,G74254,G74255,G74256,G74257,G74258,G74259,G74260,
       G74261,G74262,G74263,G74264,G74265,G74266,G74267,G74268,G74269,G74270,G74271,G74272,G74273,G74274,G74275,G74276,G74277,G74278,G74279,G74280,
       G74281,G74282,G74283,G74284,G74285,G74286,G74287,G74288,G74289,G74290,G74291,G74292,G74293,G74294,G74295,G74296,G74297,G74298,G74299,G74300,
       G74301,G74302,G74303,G74304,G74305,G74306,G74307,G74308,G74309,G74310,G74311,G74312,G74313,G74314,G74315,G74316,G74317,G74318,G74319,G74320,
       G74321,G74322,G74323,G74324,G74325,G74326,G74327,G74328,G74329,G74330,G74331,G74332,G74333,G74334,G74335,G74336,G74337,G74338,G74339,G74340,
       G74341,G74342,G74343,G74344,G74345,G74346,G74347,G74348,G74349,G74350,G74351,G74352,G74353,G74354,G74355,G74356,G74357,G74358,G74359,G74360,
       G74361,G74362,G74363,G74364,G74365,G74366,G74367,G74368,G74369,G74370,G74371,G74372,G74373,G74374,G74375,G74376,G74377,G74378,G74379,G74380,
       G74381,G74382,G74383,G74384,G74385,G74386,G74387,G74388,G74389,G74390,G74391,G74392,G74393,G74394,G74395,G74396,G74397,G74398,G74399,G74400,
       G74401,G74402,G74403,G74404,G74405,G74406,G74407,G74408,G74409,G74410,G74411,G74412,G74413,G74414,G74415,G74416,G74417,G74418,G74419,G74420,
       G74421,G74422,G74423,G74424,G74425,G74426,G74427,G74428,G74429,G74430,G74431,G74432,G74433,G74434,G74435,G74436,G74437,G74438,G74439,G74440,
       G74441,G74442,G74443,G74444,G74445,G74446,G74447,G74448,G74449,G74450,G74451,G74452,G74453,G74454,G74455,G74456,G74457,G74458,G74459,G74460,
       G74461,G74462,G74463,G74464,G74465,G74466,G74467,G74468,G74469,G74470,G74471,G74472,G74473,G74474,G74475,G74476,G74477,G74478,G74479,G74480,
       G74481,G74482,G74483,G74484,G74485,G74486,G74487,G74488,G74489,G74490,G74491,G74492,G74493,G74494,G74495,G74496,G74497,G74498,G74499,G74500,
       G74501,G74502,G74503,G74504,G74505,G74506,G74507,G74508,G74509,G74510,G74511,G74512,G74513,G74514,G74515,G74516,G74517,G74518,G74519,G74520,
       G74521,G74522,G74523,G74524,G74525,G74526,G74527,G74528,G74529,G74530,G74531,G74532,G74533,G74534,G74535,G74536,G74537,G74538,G74539,G74540,
       G74541,G74542,G74543,G74544,G74545,G74546,G74547,G74548,G74549,G74550,G74551,G74552,G74553,G74554,G74555,G74556,G74557,G74558,G74559,G74560,
       G74561,G74562,G74563,G74564,G74565,G74566,G74567,G74568,G74569,G74570,G74571,G74572,G74573,G74574,G74575,G74576,G74577,G74578,G74579,G74580,
       G74581,G74582,G74583,G74584,G74585,G74586,G74587,G74588,G74589,G74590,G74591,G74592,G74593,G74594,G74595,G74596,G74597,G74598,G74599,G74600,
       G74601,G74602,G74603,G74604,G74605,G74606,G74607,G74608,G74609,G74610,G74611,G74612,G74613,G74614,G74615,G74616,G74617,G74618,G74619,G74620,
       G74621,G74622,G74623,G74624,G74625,G74626,G74627,G74628,G74629,G74630,G74631,G74632,G74633,G74634,G74635,G74636,G74637,G74638,G74639,G74640,
       G74641,G74642,G74643,G74644,G74645,G74646,G74647,G74648,G74649,G74650,G74651,G74652,G74653,G74654,G74655,G74656,G74657,G74658,G74659,G74660,
       G74661,G74662,G74663,G74664,G74665,G74666,G74667,G74668,G74669,G74670,G74671,G74672,G74673,G74674,G74675,G74676,G74677,G74678,G74679,G74680,
       G74681,G74682,G74683,G74684,G74685,G74686,G74687,G74688,G74689,G74690,G74691,G74692,G74693,G74694,G74695,G74696,G74697,G74698,G74699,G74700,
       G74701,G74702,G74703,G74704,G74705,G74706,G74707,G74708,G74709,G74710,G74711,G74712,G74713,G74714,G74715,G74716,G74717,G74718,G74719,G74720,
       G74721,G74722,G74723,G74724,G74725,G74726,G74727,G74728,G74729,G74730,G74731,G74732,G74733,G74734,G74735,G74736,G74737,G74738,G74739,G74740,
       G74741,G74742,G74743,G74744,G74745,G74746,G74747,G74748,G74749,G74750,G74751,G74752,G74753,G74754,G74755,G74756,G74757,G74758,G74759,G74760,
       G74761,G74762,G74763,G74764,G74765,G74766,G74767,G74768,G74769,G74770,G74771,G74772,G74773,G74774,G74775,G74776,G74777,G74778,G74779,G74780,
       G74781,G74782,G74783,G74784,G74785,G74786,G74787,G74788,G74789,G74790,G74791,G74792,G74793,G74794,G74795,G74796,G74797,G74798,G74799,G74800,
       G74801,G74802,G74803,G74804,G74805,G74806,G74807,G74808,G74809,G74810,G74811,G74812,G74813,G74814,G74815,G74816,G74817,G74818,G74819,G74820,
       G74821,G74822,G74823,G74824,G74825,G74826,G74827,G74828,G74829,G74830,G74831,G74832,G74833,G74834,G74835,G74836,G74837,G74838,G74839,G74840,
       G74841,G74842,G74843,G74844,G74845,G74846,G74847,G74848,G74849,G74850,G74851,G74852,G74853,G74854,G74855,G74856,G74857,G74858,G74859,G74860,
       G74861,G74862,G74863,G74864,G74865,G74866,G74867,G74868,G74869,G74870,G74871,G74872,G74873,G74874,G74875,G74876,G74877,G74878,G74879,G74880,
       G74881,G74882,G74883,G74884,G74885,G74886,G74887,G74888,G74889,G74890,G74891,G74892,G74893,G74894,G74895,G74896,G74897,G74898,G74899,G74900,
       G74901,G74902,G74903,G74904,G74905,G74906,G74907,G74908,G74909,G74910,G74911,G74912,G74913,G74914,G74915,G74916,G74917,G74918,G74919,G74920,
       G74921,G74922,G74923,G74924,G74925,G74926,G74927,G74928,G74929,G74930,G74931,G74932,G74933,G74934,G74935,G74936,G74937,G74938,G74939,G74940,
       G74941,G74942,G74943,G74944,G74945,G74946,G74947,G74948,G74949,G74950,G74951,G74952,G74953,G74954,G74955,G74956,G74957,G74958,G74959,G74960,
       G74961,G74962,G74963,G74964,G74965,G74966,G74967,G74968,G74969,G74970,G74971,G74972,G74973,G74974,G74975,G74976,G74977,G74978,G74979,G74980,
       G74981,G74982,G74983,G74984,G74985,G74986,G74987,G74988,G74989,G74990,G74991,G74992,G74993,G74994,G74995,G74996,G74997,G74998,G74999,G75000,
       G75001,G75002,G75003,G75004,G75005,G75006,G75007,G75008,G75009,G75010,G75011,G75012,G75013,G75014,G75015,G75016,G75017,G75018,G75019,G75020,
       G75021,G75022,G75023,G75024,G75025,G75026,G75027,G75028,G75029,G75030,G75031,G75032,G75033,G75034,G75035,G75036,G75037,G75038,G75039,G75040,
       G75041,G75042,G75043,G75044,G75045,G75046,G75047,G75048,G75049,G75050,G75051,G75052,G75053,G75054,G75055,G75056,G75057,G75058,G75059,G75060,
       G75061,G75062,G75063,G75064,G75065,G75066,G75067,G75068,G75069,G75070,G75071,G75072,G75073,G75074,G75075,G75076,G75077,G75078,G75079,G75080,
       G75081,G75082,G75083,G75084,G75085,G75086,G75087,G75088,G75089,G75090,G75091,G75092,G75093,G75094,G75095,G75096,G75097,G75098,G75099,G75100,
       G75101,G75102,G75103,G75104,G75105,G75106,G75107,G75108,G75109,G75110,G75111,G75112,G75113,G75114,G75115,G75116,G75117,G75118,G75119,G75120,
       G75121,G75122,G75123,G75124,G75125,G75126,G75127,G75128,G75129,G75130,G75131,G75132,G75133,G75134,G75135,G75136,G75137,G75138,G75139,G75140,
       G75141,G75142,G75143,G75144,G75145,G75146,G75147,G75148,G75149,G75150,G75151,G75152,G75153,G75154,G75155,G75156,G75157,G75158,G75159,G75160,
       G75161,G75162,G75163,G75164,G75165,G75166,G75167,G75168,G75169,G75170,G75171,G75172,G75173,G75174,G75175,G75176,G75177,G75178,G75179,G75180,
       G75181,G75182,G75183,G75184,G75185,G75186,G75187,G75188,G75189,G75190,G75191,G75192,G75193,G75194,G75195,G75196,G75197,G75198,G75199,G75200,
       G75201,G75202,G75203,G75204,G75205,G75206,G75207,G75208,G75209,G75210,G75211,G75212,G75213,G75214,G75215,G75216,G75217,G75218,G75219,G75220,
       G75221,G75222,G75223,G75224,G75225,G75226,G75227,G75228,G75229,G75230,G75231,G75232,G75233,G75234,G75235,G75236,G75237,G75238,G75239,G75240,
       G75241,G75242,G75243,G75244,G75245,G75246,G75247,G75248,G75249,G75250,G75251,G75252,G75253,G75254,G75255,G75256,G75257,G75258,G75259,G75260,
       G75261,G75262,G75263,G75264,G75265,G75266,G75267,G75268,G75269,G75270,G75271,G75272,G75273,G75274,G75275,G75276,G75277,G75278,G75279,G75280,
       G75281,G75282,G75283,G75284,G75285,G75286,G75287,G75288,G75289,G75290,G75291,G75292,G75293,G75294,G75295,G75296,G75297,G75298,G75299,G75300,
       G75301,G75302,G75303,G75304,G75305,G75306,G75307,G75308,G75309,G75310,G75311,G75312,G75313,G75314,G75315,G75316,G75317,G75318,G75319,G75320,
       G75321,G75322,G75323,G75324,G75325,G75326,G75327,G75328,G75329,G75330,G75331,G75332,G75333,G75334,G75335,G75336,G75337,G75338,G75339,G75340,
       G75341,G75342,G75343,G75344,G75345,G75346,G75347,G75348,G75349,G75350,G75351,G75352,G75353,G75354,G75355,G75356,G75357,G75358,G75359,G75360,
       G75361,G75362,G75363,G75364,G75365,G75366,G75367,G75368,G75369,G75370,G75371,G75372,G75373,G75374,G75375,G75376,G75377,G75378,G75379,G75380,
       G75381,G75382,G75383,G75384,G75385,G75386,G75387,G75388,G75389,G75390,G75391,G75392,G75393,G75394,G75395,G75396,G75397,G75398,G75399,G75400,
       G75401,G75402,G75403,G75404,G75405,G75406,G75407,G75408,G75409,G75410,G75411,G75412,G75413,G75414,G75415,G75416,G75417,G75418,G75419,G75420,
       G75421,G75422,G75423,G75424,G75425,G75426,G75427,G75428,G75429,G75430,G75431,G75432,G75433,G75434,G75435,G75436,G75437,G75438,G75439,G75440,
       G75441,G75442,G75443,G75444,G75445,G75446,G75447,G75448,G75449,G75450,G75451,G75452,G75453,G75454,G75455,G75456,G75457,G75458,G75459,G75460,
       G75461,G75462,G75463,G75464,G75465,G75466,G75467,G75468,G75469,G75470,G75471,G75472,G75473,G75474,G75475,G75476,G75477,G75478,G75479,G75480,
       G75481,G75482,G75483,G75484,G75485,G75486,G75487,G75488,G75489,G75490,G75491,G75492,G75493,G75494,G75495,G75496,G75497,G75498,G75499,G75500,
       G75501,G75502,G75503,G75504,G75505,G75506,G75507,G75508,G75509,G75510,G75511,G75512,G75513,G75514,G75515,G75516,G75517,G75518,G75519,G75520,
       G75521,G75522,G75523,G75524,G75525,G75526,G75527,G75528,G75529,G75530,G75531,G75532,G75533,G75534,G75535,G75536,G75537,G75538,G75539,G75540,
       G75541,G75542,G75543,G75544,G75545,G75546,G75547,G75548,G75549,G75550,G75551,G75552,G75553,G75554,G75555,G75556,G75557,G75558,G75559,G75560,
       G75561,G75562,G75563,G75564,G75565,G75566,G75567,G75568,G75569,G75570,G75571,G75572,G75573,G75574,G75575,G75576,G75577,G75578,G75579,G75580,
       G75581,G75582,G75583,G75584,G75585,G75586,G75587,G75588,G75589,G75590,G75591,G75592,G75593,G75594,G75595,G75596,G75597,G75598,G75599,G75600,
       G75601,G75602,G75603,G75604,G75605,G75606,G75607,G75608,G75609,G75610,G75611,G75612,G75613,G75614,G75615,G75616,G75617,G75618,G75619,G75620,
       G75621,G75622,G75623,G75624,G75625,G75626,G75627,G75628,G75629,G75630,G75631,G75632,G75633,G75634,G75635,G75636,G75637,G75638,G75639,G75640,
       G75641,G75642,G75643,G75644,G75645,G75646,G75647,G75648,G75649,G75650,G75651,G75652,G75653,G75654,G75655,G75656,G75657,G75658,G75659,G75660,
       G75661,G75662,G75663,G75664,G75665,G75666,G75667,G75668,G75669,G75670,G75671,G75672,G75673,G75674,G75675,G75676,G75677,G75678,G75679,G75680,
       G75681,G75682,G75683,G75684,G75685,G75686,G75687,G75688,G75689,G75690,G75691,G75692,G75693,G75694,G75695,G75696,G75697,G75698,G75699,G75700,
       G75701,G75702,G75703,G75704,G75705,G75706,G75707,G75708,G75709,G75710,G75711,G75712,G75713,G75714,G75715,G75716,G75717,G75718,G75719,G75720,
       G75721,G75722,G75723,G75724,G75725,G75726,G75727,G75728,G75729,G75730,G75731,G75732,G75733,G75734,G75735,G75736,G75737,G75738,G75739,G75740,
       G75741,G75742,G75743,G75744,G75745,G75746,G75747,G75748,G75749,G75750,G75751,G75752,G75753,G75754,G75755,G75756,G75757,G75758,G75759,G75760,
       G75761,G75762,G75763,G75764,G75765,G75766,G75767,G75768,G75769,G75770,G75771,G75772,G75773,G75774,G75775,G75776,G75777,G75778,G75779,G75780,
       G75781,G75782,G75783,G75784,G75785,G75786,G75787,G75788,G75789,G75790,G75791,G75792,G75793,G75794,G75795,G75796,G75797,G75798,G75799,G75800,
       G75801,G75802,G75803,G75804,G75805,G75806,G75807,G75808,G75809,G75810,G75811,G75812,G75813,G75814,G75815,G75816,G75817,G75818,G75819,G75820,
       G75821,G75822,G75823,G75824,G75825,G75826,G75827,G75828,G75829,G75830,G75831,G75832,G75833,G75834,G75835,G75836,G75837,G75838,G75839,G75840,
       G75841,G75842,G75843,G75844,G75845,G75846,G75847,G75848,G75849,G75850,G75851,G75852,G75853,G75854,G75855,G75856,G75857,G75858,G75859,G75860,
       G75861,G75862,G75863,G75864,G75865,G75866,G75867,G75868,G75869,G75870,G75871,G75872,G75873,G75874,G75875,G75876,G75877,G75878,G75879,G75880,
       G75881,G75882,G75883,G75884,G75885,G75886,G75887,G75888,G75889,G75890,G75891,G75892,G75893,G75894,G75895,G75896,G75897,G75898,G75899,G75900,
       G75901,G75902,G75903,G75904,G75905,G75906,G75907,G75908,G75909,G75910,G75911,G75912,G75913,G75914,G75915,G75916,G75917,G75918,G75919,G75920,
       G75921,G75922,G75923,G75924,G75925,G75926,G75927,G75928,G75929,G75930,G75931,G75932,G75933,G75934,G75935,G75936,G75937,G75938,G75939,G75940,
       G75941,G75942,G75943,G75944,G75945,G75946,G75947,G75948,G75949,G75950,G75951,G75952,G75953,G75954,G75955,G75956,G75957,G75958,G75959,G75960,
       G75961,G75962,G75963,G75964,G75965,G75966,G75967,G75968,G75969,G75970,G75971,G75972,G75973,G75974,G75975,G75976,G75977,G75978,G75979,G75980,
       G75981,G75982,G75983,G75984,G75985,G75986,G75987,G75988,G75989,G75990,G75991,G75992,G75993,G75994,G75995,G75996,G75997,G75998,G75999,G76000,
       G76001,G76002,G76003,G76004,G76005,G76006,G76007,G76008,G76009,G76010,G76011,G76012,G76013,G76014,G76015,G76016,G76017,G76018,G76019,G76020,
       G76021,G76022,G76023,G76024,G76025,G76026,G76027,G76028,G76029,G76030,G76031,G76032,G76033,G76034,G76035,G76036,G76037,G76038,G76039,G76040,
       G76041,G76042,G76043,G76044,G76045,G76046,G76047,G76048,G76049,G76050,G76051,G76052,G76053,G76054,G76055,G76056,G76057,G76058,G76059,G76060,
       G76061,G76062,G76063,G76064,G76065,G76066,G76067,G76068,G76069,G76070,G76071,G76072,G76073,G76074,G76075,G76076,G76077,G76078,G76079,G76080,
       G76081,G76082,G76083,G76084,G76085,G76086,G76087,G76088,G76089,G76090,G76091,G76092,G76093,G76094,G76095,G76096,G76097,G76098,G76099,G76100,
       G76101,G76102,G76103,G76104,G76105,G76106,G76107,G76108,G76109,G76110,G76111,G76112,G76113,G76114,G76115,G76116,G76117,G76118,G76119,G76120,
       G76121,G76122,G76123,G76124,G76125,G76126,G76127,G76128,G76129,G76130,G76131,G76132,G76133,G76134,G76135,G76136,G76137,G76138,G76139,G76140,
       G76141,G76142,G76143,G76144,G76145,G76146,G76147,G76148,G76149,G76150,G76151,G76152,G76153,G76154,G76155,G76156,G76157,G76158,G76159,G76160,
       G76161,G76162,G76163,G76164,G76165,G76166,G76167,G76168,G76169,G76170,G76171,G76172,G76173,G76174,G76175,G76176,G76177,G76178,G76179,G76180,
       G76181,G76182,G76183,G76184,G76185,G76186,G76187,G76188,G76189,G76190,G76191,G76192,G76193,G76194,G76195,G76196,G76197,G76198,G76199,G76200,
       G76201,G76202,G76203,G76204,G76205,G76206,G76207,G76208,G76209,G76210,G76211,G76212,G76213,G76214,G76215,G76216,G76217,G76218,G76219,G76220,
       G76221,G76222,G76223,G76224,G76225,G76226,G76227,G76228,G76229,G76230,G76231,G76232,G76233,G76234,G76235,G76236,G76237,G76238,G76239,G76240,
       G76241,G76242,G76243,G76244,G76245,G76246,G76247,G76248,G76249,G76250,G76251,G76252,G76253,G76254,G76255,G76256,G76257,G76258,G76259,G76260,
       G76261,G76262,G76263,G76264,G76265,G76266,G76267,G76268,G76269,G76270,G76271,G76272,G76273,G76274,G76275,G76276,G76277,G76278,G76279,G76280,
       G76281,G76282,G76283,G76284,G76285,G76286,G76287,G76288,G76289,G76290,G76291,G76292,G76293,G76294,G76295,G76296,G76297,G76298,G76299,G76300,
       G76301,G76302,G76303,G76304,G76305,G76306,G76307,G76308,G76309,G76310,G76311,G76312,G76313,G76314,G76315,G76316,G76317,G76318,G76319,G76320,
       G76321,G76322,G76323,G76324,G76325,G76326,G76327,G76328,G76329,G76330,G76331,G76332,G76333,G76334,G76335,G76336,G76337,G76338,G76339,G76340,
       G76341,G76342,G76343,G76344,G76345,G76346,G76347,G76348,G76349,G76350,G76351,G76352,G76353,G76354,G76355,G76356,G76357,G76358,G76359,G76360,
       G76361,G76362,G76363,G76364,G76365,G76366,G76367,G76368,G76369,G76370,G76371,G76372,G76373,G76374,G76375,G76376,G76377,G76378,G76379,G76380,
       G76381,G76382,G76383,G76384,G76385,G76386,G76387,G76388,G76389,G76390,G76391,G76392,G76393,G76394,G76395,G76396,G76397,G76398,G76399,G76400,
       G76401,G76402,G76403,G76404,G76405,G76406,G76407,G76408,G76409,G76410,G76411,G76412,G76413,G76414,G76415,G76416,G76417,G76418,G76419,G76420,
       G76421,G76422,G76423,G76424,G76425,G76426,G76427,G76428,G76429,G76430,G76431,G76432,G76433,G76434,G76435,G76436,G76437,G76438,G76439,G76440,
       G76441,G76442,G76443,G76444,G76445,G76446,G76447,G76448,G76449,G76450,G76451,G76452,G76453,G76454,G76455,G76456,G76457,G76458,G76459,G76460,
       G76461,G76462,G76463,G76464,G76465,G76466,G76467,G76468,G76469,G76470,G76471,G76472,G76473,G76474,G76475,G76476,G76477,G76478,G76479,G76480,
       G76481,G76482,G76483,G76484,G76485,G76486,G76487,G76488,G76489,G76490,G76491,G76492,G76493,G76494,G76495,G76496,G76497,G76498,G76499,G76500,
       G76501,G76502,G76503,G76504,G76505,G76506,G76507,G76508,G76509,G76510,G76511,G76512,G76513,G76514,G76515,G76516,G76517,G76518,G76519,G76520,
       G76521,G76522,G76523,G76524,G76525,G76526,G76527,G76528,G76529,G76530,G76531,G76532,G76533,G76534,G76535,G76536,G76537,G76538,G76539,G76540,
       G76541,G76542,G76543,G76544,G76545,G76546,G76547,G76548,G76549,G76550,G76551,G76552,G76553,G76554,G76555,G76556,G76557,G76558,G76559,G76560,
       G76561,G76562,G76563,G76564,G76565,G76566,G76567,G76568,G76569,G76570,G76571,G76572,G76573,G76574,G76575,G76576,G76577,G76578,G76579,G76580,
       G76581,G76582,G76583,G76584,G76585,G76586,G76587,G76588,G76589,G76590,G76591,G76592,G76593,G76594,G76595,G76596,G76597,G76598,G76599,G76600,
       G76601,G76602,G76603,G76604,G76605,G76606,G76607,G76608,G76609,G76610,G76611,G76612,G76613,G76614,G76615,G76616,G76617,G76618,G76619,G76620,
       G76621,G76622,G76623,G76624,G76625,G76626,G76627,G76628,G76629,G76630,G76631,G76632,G76633,G76634,G76635,G76636,G76637,G76638,G76639,G76640,
       G76641,G76642,G76643,G76644,G76645,G76646,G76647,G76648,G76649,G76650,G76651,G76652,G76653,G76654,G76655,G76656,G76657,G76658,G76659,G76660,
       G76661,G76662,G76663,G76664,G76665,G76666,G76667,G76668,G76669,G76670,G76671,G76672,G76673,G76674,G76675,G76676,G76677,G76678,G76679,G76680,
       G76681,G76682,G76683,G76684,G76685,G76686,G76687,G76688,G76689,G76690,G76691,G76692,G76693,G76694,G76695,G76696,G76697,G76698,G76699,G76700,
       G76701,G76702,G76703,G76704,G76705,G76706,G76707,G76708,G76709,G76710,G76711,G76712,G76713,G76714,G76715,G76716,G76717,G76718,G76719,G76720,
       G76721,G76722,G76723,G76724,G76725,G76726,G76727,G76728,G76729,G76730,G76731,G76732,G76733,G76734,G76735,G76736,G76737,G76738,G76739,G76740,
       G76741,G76742,G76743,G76744,G76745,G76746,G76747,G76748,G76749,G76750,G76751,G76752,G76753,G76754,G76755,G76756,G76757,G76758,G76759,G76760,
       G76761,G76762,G76763,G76764,G76765,G76766,G76767,G76768,G76769,G76770,G76771,G76772,G76773,G76774,G76775,G76776,G76777,G76778,G76779,G76780,
       G76781,G76782,G76783,G76784,G76785,G76786,G76787,G76788,G76789,G76790,G76791,G76792,G76793,G76794,G76795,G76796,G76797,G76798,G76799,G76800,
       G76801,G76802,G76803,G76804,G76805,G76806,G76807,G76808,G76809,G76810,G76811,G76812,G76813,G76814,G76815,G76816,G76817,G76818,G76819,G76820,
       G76821,G76822,G76823,G76824,G76825,G76826,G76827,G76828,G76829,G76830,G76831,G76832,G76833,G76834,G76835,G76836,G76837,G76838,G76839,G76840,
       G76841,G76842,G76843,G76844,G76845,G76846,G76847,G76848,G76849,G76850,G76851,G76852,G76853,G76854,G76855,G76856,G76857,G76858,G76859,G76860,
       G76861,G76862,G76863,G76864,G76865,G76866,G76867,G76868,G76869,G76870,G76871,G76872,G76873,G76874,G76875,G76876,G76877,G76878,G76879,G76880,
       G76881,G76882,G76883,G76884,G76885,G76886,G76887,G76888,G76889,G76890,G76891,G76892,G76893,G76894,G76895,G76896,G76897,G76898,G76899,G76900,
       G76901,G76902,G76903,G76904,G76905,G76906,G76907,G76908,G76909,G76910,G76911,G76912,G76913,G76914,G76915,G76916,G76917,G76918,G76919,G76920,
       G76921,G76922,G76923,G76924,G76925,G76926,G76927,G76928,G76929,G76930,G76931,G76932,G76933,G76934,G76935,G76936,G76937,G76938,G76939,G76940,
       G76941,G76942,G76943,G76944,G76945,G76946,G76947,G76948,G76949,G76950,G76951,G76952,G76953,G76954,G76955,G76956,G76957,G76958,G76959,G76960,
       G76961,G76962,G76963,G76964,G76965,G76966,G76967,G76968,G76969,G76970,G76971,G76972,G76973,G76974,G76975,G76976,G76977,G76978,G76979,G76980,
       G76981,G76982,G76983,G76984,G76985,G76986,G76987,G76988,G76989,G76990,G76991,G76992,G76993,G76994,G76995,G76996,G76997,G76998,G76999,G77000,
       G77001,G77002,G77003,G77004,G77005,G77006,G77007,G77008,G77009,G77010,G77011,G77012,G77013,G77014,G77015,G77016,G77017,G77018,G77019,G77020,
       G77021,G77022,G77023,G77024,G77025,G77026,G77027,G77028,G77029,G77030,G77031,G77032,G77033,G77034,G77035,G77036,G77037,G77038,G77039,G77040,
       G77041,G77042,G77043,G77044,G77045,G77046,G77047,G77048,G77049,G77050,G77051,G77052,G77053,G77054,G77055,G77056,G77057,G77058,G77059,G77060,
       G77061,G77062,G77063,G77064,G77065,G77066,G77067,G77068,G77069,G77070,G77071,G77072,G77073,G77074,G77075,G77076,G77077,G77078,G77079,G77080,
       G77081,G77082,G77083,G77084,G77085,G77086,G77087,G77088,G77089,G77090,G77091,G77092,G77093,G77094,G77095,G77096,G77097,G77098,G77099,G77100,
       G77101,G77102,G77103,G77104,G77105,G77106,G77107,G77108,G77109,G77110,G77111,G77112,G77113,G77114,G77115,G77116,G77117,G77118,G77119,G77120,
       G77121,G77122,G77123,G77124,G77125,G77126,G77127,G77128,G77129,G77130,G77131,G77132,G77133,G77134,G77135,G77136,G77137,G77138,G77139,G77140,
       G77141,G77142,G77143,G77144,G77145,G77146,G77147,G77148,G77149,G77150,G77151,G77152,G77153,G77154,G77155,G77156,G77157,G77158,G77159,G77160,
       G77161,G77162,G77163,G77164,G77165,G77166,G77167,G77168,G77169,G77170,G77171,G77172,G77173,G77174,G77175,G77176,G77177,G77178,G77179,G77180,
       G77181,G77182,G77183,G77184,G77185,G77186,G77187,G77188,G77189,G77190,G77191,G77192,G77193,G77194,G77195,G77196,G77197,G77198,G77199,G77200,
       G77201,G77202,G77203,G77204,G77205,G77206,G77207,G77208,G77209,G77210,G77211,G77212,G77213,G77214,G77215,G77216,G77217,G77218,G77219,G77220,
       G77221,G77222,G77223,G77224,G77225,G77226,G77227,G77228,G77229,G77230,G77231,G77232,G77233,G77234,G77235,G77236,G77237,G77238,G77239,G77240,
       G77241,G77242,G77243,G77244,G77245,G77246,G77247,G77248,G77249,G77250,G77251,G77252,G77253,G77254,G77255,G77256,G77257,G77258,G77259,G77260,
       G77261,G77262,G77263,G77264,G77265,G77266,G77267,G77268,G77269,G77270,G77271,G77272,G77273,G77274,G77275,G77276,G77277,G77278,G77279,G77280,
       G77281,G77282,G77283,G77284,G77285,G77286,G77287,G77288,G77289,G77290,G77291,G77292,G77293,G77294,G77295,G77296,G77297,G77298,G77299,G77300,
       G77301,G77302,G77303,G77304,G77305,G77306,G77307,G77308,G77309,G77310,G77311,G77312,G77313,G77314,G77315,G77316,G77317,G77318,G77319,G77320,
       G77321,G77322,G77323,G77324,G77325,G77326,G77327,G77328,G77329,G77330,G77331,G77332,G77333,G77334,G77335,G77336,G77337,G77338,G77339,G77340,
       G77341,G77342,G77343,G77344,G77345,G77346,G77347,G77348,G77349,G77350,G77351,G77352,G77353,G77354,G77355,G77356,G77357,G77358,G77359,G77360,
       G77361,G77362,G77363,G77364,G77365,G77366,G77367,G77368,G77369,G77370,G77371,G77372,G77373,G77374,G77375,G77376,G77377,G77378,G77379,G77380,
       G77381,G77382,G77383,G77384,G77385,G77386,G77387,G77388,G77389,G77390,G77391,G77392,G77393,G77394,G77395,G77396,G77397,G77398,G77399,G77400,
       G77401,G77402,G77403,G77404,G77405,G77406,G77407,G77408,G77409,G77410,G77411,G77412,G77413,G77414,G77415,G77416,G77417,G77418,G77419,G77420,
       G77421,G77422,G77423,G77424,G77425,G77426,G77427,G77428,G77429,G77430,G77431,G77432,G77433,G77434,G77435,G77436,G77437,G77438,G77439,G77440,
       G77441,G77442,G77443,G77444,G77445,G77446,G77447,G77448,G77449,G77450,G77451,G77452,G77453,G77454,G77455,G77456,G77457,G77458,G77459,G77460,
       G77461,G77462,G77463,G77464,G77465,G77466,G77467,G77468,G77469,G77470,G77471,G77472,G77473,G77474,G77475,G77476,G77477,G77478,G77479,G77480,
       G77481,G77482,G77483,G77484,G77485,G77486,G77487,G77488,G77489,G77490,G77491,G77492,G77493,G77494,G77495,G77496,G77497,G77498,G77499,G77500,
       G77501,G77502,G77503,G77504,G77505,G77506,G77507,G77508,G77509,G77510,G77511,G77512,G77513,G77514,G77515,G77516,G77517,G77518,G77519,G77520,
       G77521,G77522,G77523,G77524,G77525,G77526,G77527,G77528,G77529,G77530,G77531,G77532,G77533,G77534,G77535,G77536,G77537,G77538,G77539,G77540,
       G77541,G77542,G77543,G77544,G77545,G77546,G77547,G77548,G77549,G77550,G77551,G77552,G77553,G77554,G77555,G77556,G77557,G77558,G77559,G77560,
       G77561,G77562,G77563,G77564,G77565,G77566,G77567,G77568,G77569,G77570,G77571,G77572,G77573,G77574,G77575,G77576,G77577,G77578,G77579,G77580,
       G77581,G77582,G77583,G77584,G77585,G77586,G77587,G77588,G77589,G77590,G77591,G77592,G77593,G77594,G77595,G77596,G77597,G77598,G77599,G77600,
       G77601,G77602,G77603,G77604,G77605,G77606,G77607,G77608,G77609,G77610,G77611,G77612,G77613,G77614,G77615,G77616,G77617,G77618,G77619,G77620,
       G77621,G77622,G77623,G77624,G77625,G77626,G77627,G77628,G77629,G77630,G77631,G77632,G77633,G77634,G77635,G77636,G77637,G77638,G77639,G77640,
       G77641,G77642,G77643,G77644,G77645,G77646,G77647,G77648,G77649,G77650,G77651,G77652,G77653,G77654,G77655,G77656,G77657,G77658,G77659,G77660,
       G77661,G77662,G77663,G77664,G77665,G77666,G77667,G77668,G77669,G77670,G77671,G77672,G77673,G77674,G77675,G77676,G77677,G77678,G77679,G77680,
       G77681,G77682,G77683,G77684,G77685,G77686,G77687,G77688,G77689,G77690,G77691,G77692,G77693,G77694,G77695,G77696,G77697,G77698,G77699,G77700,
       G77701,G77702,G77703,G77704,G77705,G77706,G77707,G77708,G77709,G77710,G77711,G77712,G77713,G77714,G77715,G77716,G77717,G77718,G77719,G77720,
       G77721,G77722,G77723,G77724,G77725,G77726,G77727,G77728,G77729,G77730,G77731,G77732,G77733,G77734,G77735,G77736,G77737,G77738,G77739,G77740,
       G77741,G77742,G77743,G77744,G77745,G77746,G77747,G77748,G77749,G77750,G77751,G77752,G77753,G77754,G77755,G77756,G77757,G77758,G77759,G77760,
       G77761,G77762,G77763,G77764,G77765,G77766,G77767,G77768,G77769,G77770,G77771,G77772,G77773,G77774,G77775,G77776,G77777,G77778,G77779,G77780,
       G77781,G77782,G77783,G77784,G77785,G77786,G77787,G77788,G77789,G77790,G77791,G77792,G77793,G77794,G77795,G77796,G77797,G77798,G77799,G77800,
       G77801,G77802,G77803,G77804,G77805,G77806,G77807,G77808,G77809,G77810,G77811,G77812,G77813,G77814,G77815,G77816,G77817,G77818,G77819,G77820,
       G77821,G77822,G77823,G77824,G77825,G77826,G77827,G77828,G77829,G77830,G77831,G77832,G77833,G77834,G77835,G77836,G77837,G77838,G77839,G77840,
       G77841,G77842,G77843,G77844,G77845,G77846,G77847,G77848,G77849,G77850,G77851,G77852,G77853,G77854,G77855,G77856,G77857,G77858,G77859,G77860,
       G77861,G77862,G77863,G77864,G77865,G77866,G77867,G77868,G77869,G77870,G77871,G77872,G77873,G77874,G77875,G77876,G77877,G77878,G77879,G77880,
       G77881,G77882,G77883,G77884,G77885,G77886,G77887,G77888,G77889,G77890,G77891,G77892,G77893,G77894,G77895,G77896,G77897,G77898,G77899,G77900,
       G77901,G77902,G77903,G77904,G77905,G77906,G77907,G77908,G77909,G77910,G77911,G77912,G77913,G77914,G77915,G77916,G77917,G77918,G77919,G77920,
       G77921,G77922,G77923,G77924,G77925,G77926,G77927,G77928,G77929,G77930,G77931,G77932,G77933,G77934,G77935,G77936,G77937,G77938,G77939,G77940,
       G77941,G77942,G77943,G77944,G77945,G77946,G77947,G77948,G77949,G77950,G77951,G77952,G77953,G77954,G77955,G77956,G77957,G77958,G77959,G77960,
       G77961,G77962,G77963,G77964,G77965,G77966,G77967,G77968,G77969,G77970,G77971,G77972,G77973,G77974,G77975,G77976,G77977,G77978,G77979,G77980,
       G77981,G77982,G77983,G77984,G77985,G77986,G77987,G77988,G77989,G77990,G77991,G77992,G77993,G77994,G77995,G77996,G77997,G77998,G77999,G78000,
       G78001,G78002,G78003,G78004,G78005,G78006,G78007,G78008,G78009,G78010,G78011,G78012,G78013,G78014,G78015,G78016,G78017,G78018,G78019,G78020,
       G78021,G78022,G78023,G78024,G78025,G78026,G78027,G78028,G78029,G78030,G78031,G78032,G78033,G78034,G78035,G78036,G78037,G78038,G78039,G78040,
       G78041,G78042,G78043,G78044,G78045,G78046,G78047,G78048,G78049,G78050,G78051,G78052,G78053,G78054,G78055,G78056,G78057,G78058,G78059,G78060,
       G78061,G78062,G78063,G78064,G78065,G78066,G78067,G78068,G78069,G78070,G78071,G78072,G78073,G78074,G78075,G78076,G78077,G78078,G78079,G78080,
       G78081,G78082,G78083,G78084,G78085,G78086,G78087,G78088,G78089,G78090,G78091,G78092,G78093,G78094,G78095,G78096,G78097,G78098,G78099,G78100,
       G78101,G78102,G78103,G78104,G78105,G78106,G78107,G78108,G78109,G78110,G78111,G78112,G78113,G78114,G78115,G78116,G78117,G78118,G78119,G78120,
       G78121,G78122,G78123,G78124,G78125,G78126,G78127,G78128,G78129,G78130,G78131,G78132,G78133,G78134,G78135,G78136,G78137,G78138,G78139,G78140,
       G78141,G78142,G78143,G78144,G78145,G78146,G78147,G78148,G78149,G78150,G78151,G78152,G78153,G78154,G78155,G78156,G78157,G78158,G78159,G78160,
       G78161,G78162,G78163,G78164,G78165,G78166,G78167,G78168,G78169,G78170,G78171,G78172,G78173,G78174,G78175,G78176,G78177,G78178,G78179,G78180,
       G78181,G78182,G78183,G78184,G78185,G78186,G78187,G78188,G78189,G78190,G78191,G78192,G78193,G78194,G78195,G78196,G78197,G78198,G78199,G78200,
       G78201,G78202,G78203,G78204,G78205,G78206,G78207,G78208,G78209,G78210,G78211,G78212,G78213,G78214,G78215,G78216,G78217,G78218,G78219,G78220,
       G78221,G78222,G78223,G78224,G78225,G78226,G78227,G78228,G78229,G78230,G78231,G78232,G78233,G78234,G78235,G78236,G78237,G78238,G78239,G78240,
       G78241,G78242,G78243,G78244,G78245,G78246,G78247,G78248,G78249,G78250,G78251,G78252,G78253,G78254,G78255,G78256,G78257,G78258,G78259,G78260,
       G78261,G78262,G78263,G78264,G78265,G78266,G78267,G78268,G78269,G78270,G78271,G78272,G78273,G78274,G78275,G78276,G78277,G78278,G78279,G78280,
       G78281,G78282,G78283,G78284,G78285,G78286,G78287,G78288,G78289,G78290,G78291,G78292,G78293,G78294,G78295,G78296,G78297,G78298,G78299,G78300,
       G78301,G78302,G78303,G78304,G78305,G78306,G78307,G78308,G78309,G78310,G78311,G78312,G78313,G78314,G78315,G78316,G78317,G78318,G78319,G78320,
       G78321,G78322,G78323,G78324,G78325,G78326,G78327,G78328,G78329,G78330,G78331,G78332,G78333,G78334,G78335,G78336,G78337,G78338,G78339,G78340,
       G78341,G78342,G78343,G78344,G78345,G78346,G78347,G78348,G78349,G78350,G78351,G78352,G78353,G78354,G78355,G78356,G78357,G78358,G78359,G78360,
       G78361,G78362,G78363,G78364,G78365,G78366,G78367,G78368,G78369,G78370,G78371,G78372,G78373,G78374,G78375,G78376,G78377,G78378,G78379,G78380,
       G78381,G78382,G78383,G78384,G78385,G78386,G78387,G78388,G78389,G78390,G78391,G78392,G78393,G78394,G78395,G78396,G78397,G78398,G78399,G78400,
       G78401,G78402,G78403,G78404,G78405,G78406,G78407,G78408,G78409,G78410,G78411,G78412,G78413,G78414,G78415,G78416,G78417,G78418,G78419,G78420,
       G78421,G78422,G78423,G78424,G78425,G78426,G78427,G78428,G78429,G78430,G78431,G78432,G78433,G78434,G78435,G78436,G78437,G78438,G78439,G78440,
       G78441,G78442,G78443,G78444,G78445,G78446,G78447,G78448,G78449,G78450,G78451,G78452,G78453,G78454,G78455,G78456,G78457,G78458,G78459,G78460,
       G78461,G78462,G78463,G78464,G78465,G78466,G78467,G78468,G78469,G78470,G78471,G78472,G78473,G78474,G78475,G78476,G78477,G78478,G78479,G78480,
       G78481,G78482,G78483,G78484,G78485,G78486,G78487,G78488,G78489,G78490,G78491,G78492,G78493,G78494,G78495,G78496,G78497,G78498,G78499,G78500,
       G78501,G78502,G78503,G78504,G78505,G78506,G78507,G78508,G78509,G78510,G78511,G78512,G78513,G78514,G78515,G78516,G78517,G78518,G78519,G78520,
       G78521,G78522,G78523,G78524,G78525,G78526,G78527,G78528,G78529,G78530,G78531,G78532,G78533,G78534,G78535,G78536,G78537,G78538,G78539,G78540,
       G78541,G78542,G78543,G78544,G78545,G78546,G78547,G78548,G78549,G78550,G78551,G78552,G78553,G78554,G78555,G78556,G78557,G78558,G78559,G78560,
       G78561,G78562,G78563,G78564,G78565,G78566,G78567,G78568,G78569,G78570,G78571,G78572,G78573,G78574,G78575,G78576,G78577,G78578,G78579,G78580,
       G78581,G78582,G78583,G78584,G78585,G78586,G78587,G78588,G78589,G78590,G78591,G78592,G78593,G78594,G78595,G78596,G78597,G78598,G78599,G78600,
       G78601,G78602,G78603,G78604,G78605,G78606,G78607,G78608,G78609,G78610,G78611,G78612,G78613,G78614,G78615,G78616,G78617,G78618,G78619,G78620,
       G78621,G78622,G78623,G78624,G78625,G78626,G78627,G78628,G78629,G78630,G78631,G78632,G78633,G78634,G78635,G78636,G78637,G78638,G78639,G78640,
       G78641,G78642,G78643,G78644,G78645,G78646,G78647,G78648,G78649,G78650,G78651,G78652,G78653,G78654,G78655,G78656,G78657,G78658,G78659,G78660,
       G78661,G78662,G78663,G78664,G78665,G78666,G78667,G78668,G78669,G78670,G78671,G78672,G78673,G78674,G78675,G78676,G78677,G78678,G78679,G78680,
       G78681,G78682,G78683,G78684,G78685,G78686,G78687,G78688,G78689,G78690,G78691,G78692,G78693,G78694,G78695,G78696,G78697,G78698,G78699,G78700,
       G78701,G78702,G78703,G78704,G78705,G78706,G78707,G78708,G78709,G78710,G78711,G78712,G78713,G78714,G78715,G78716,G78717,G78718,G78719,G78720,
       G78721,G78722,G78723,G78724,G78725,G78726,G78727,G78728,G78729,G78730,G78731,G78732,G78733,G78734,G78735,G78736,G78737,G78738,G78739,G78740,
       G78741,G78742,G78743,G78744,G78745,G78746,G78747,G78748,G78749,G78750,G78751,G78752,G78753,G78754,G78755,G78756,G78757,G78758,G78759,G78760,
       G78761,G78762,G78763,G78764,G78765,G78766,G78767,G78768,G78769,G78770,G78771,G78772,G78773,G78774,G78775,G78776,G78777,G78778,G78779,G78780,
       G78781,G78782,G78783,G78784,G78785,G78786,G78787,G78788,G78789,G78790,G78791,G78792,G78793,G78794,G78795,G78796,G78797,G78798,G78799,G78800,
       G78801,G78802,G78803,G78804,G78805,G78806,G78807,G78808,G78809,G78810,G78811,G78812,G78813,G78814,G78815,G78816,G78817,G78818,G78819,G78820,
       G78821,G78822,G78823,G78824,G78825,G78826,G78827,G78828,G78829,G78830,G78831,G78832,G78833,G78834,G78835,G78836,G78837,G78838,G78839,G78840,
       G78841,G78842,G78843,G78844,G78845,G78846,G78847,G78848,G78849,G78850,G78851,G78852,G78853,G78854,G78855,G78856,G78857,G78858,G78859,G78860,
       G78861,G78862,G78863,G78864,G78865,G78866,G78867,G78868,G78869,G78870,G78871,G78872,G78873,G78874,G78875,G78876,G78877,G78878,G78879,G78880,
       G78881,G78882,G78883,G78884,G78885,G78886,G78887,G78888,G78889,G78890,G78891,G78892,G78893,G78894,G78895,G78896,G78897,G78898,G78899,G78900,
       G78901,G78902,G78903,G78904,G78905,G78906,G78907,G78908,G78909,G78910,G78911,G78912,G78913,G78914,G78915,G78916,G78917,G78918,G78919,G78920,
       G78921,G78922,G78923,G78924,G78925,G78926,G78927,G78928,G78929,G78930,G78931,G78932,G78933,G78934,G78935,G78936,G78937,G78938,G78939,G78940,
       G78941,G78942,G78943,G78944,G78945,G78946,G78947,G78948,G78949,G78950,G78951,G78952,G78953,G78954,G78955,G78956,G78957,G78958,G78959,G78960,
       G78961,G78962,G78963,G78964,G78965,G78966,G78967,G78968,G78969,G78970,G78971,G78972,G78973,G78974,G78975,G78976,G78977,G78978,G78979,G78980,
       G78981,G78982,G78983,G78984,G78985,G78986,G78987,G78988,G78989,G78990,G78991,G78992,G78993,G78994,G78995,G78996,G78997,G78998,G78999,G79000,
       G79001,G79002,G79003,G79004,G79005,G79006,G79007,G79008,G79009,G79010,G79011,G79012,G79013,G79014,G79015,G79016,G79017,G79018,G79019,G79020,
       G79021,G79022,G79023,G79024,G79025,G79026,G79027,G79028,G79029,G79030,G79031,G79032,G79033,G79034,G79035,G79036,G79037,G79038,G79039,G79040,
       G79041,G79042,G79043,G79044,G79045,G79046,G79047,G79048,G79049,G79050,G79051,G79052,G79053,G79054,G79055,G79056,G79057,G79058,G79059,G79060,
       G79061,G79062,G79063,G79064,G79065,G79066,G79067,G79068,G79069,G79070,G79071,G79072,G79073,G79074,G79075,G79076,G79077,G79078,G79079,G79080,
       G79081,G79082,G79083,G79084,G79085,G79086,G79087,G79088,G79089,G79090,G79091,G79092,G79093,G79094,G79095,G79096,G79097,G79098,G79099,G79100,
       G79101,G79102,G79103,G79104,G79105,G79106,G79107,G79108,G79109,G79110,G79111,G79112,G79113,G79114,G79115,G79116,G79117,G79118,G79119,G79120,
       G79121,G79122,G79123,G79124,G79125,G79126,G79127,G79128,G79129,G79130,G79131,G79132,G79133,G79134,G79135,G79136,G79137,G79138,G79139,G79140,
       G79141,G79142,G79143,G79144,G79145,G79146,G79147,G79148,G79149,G79150,G79151,G79152,G79153,G79154,G79155,G79156,G79157,G79158,G79159,G79160,
       G79161,G79162,G79163,G79164,G79165,G79166,G79167,G79168,G79169,G79170,G79171,G79172,G79173,G79174,G79175,G79176,G79177,G79178,G79179,G79180,
       G79181,G79182,G79183,G79184,G79185,G79186,G79187,G79188,G79189,G79190,G79191,G79192,G79193,G79194,G79195,G79196,G79197,G79198,G79199,G79200,
       G79201,G79202,G79203,G79204,G79205,G79206,G79207,G79208,G79209,G79210,G79211,G79212,G79213,G79214,G79215,G79216,G79217,G79218,G79219,G79220,
       G79221,G79222,G79223,G79224,G79225,G79226,G79227,G79228,G79229,G79230,G79231,G79232,G79233,G79234,G79235,G79236,G79237,G79238,G79239,G79240,
       G79241,G79242,G79243,G79244,G79245,G79246,G79247,G79248,G79249,G79250,G79251,G79252,G79253,G79254,G79255,G79256,G79257,G79258,G79259,G79260,
       G79261,G79262,G79263,G79264,G79265,G79266,G79267,G79268,G79269,G79270,G79271,G79272,G79273,G79274,G79275,G79276,G79277,G79278,G79279,G79280,
       G79281,G79282,G79283,G79284,G79285,G79286,G79287,G79288,G79289,G79290,G79291,G79292,G79293,G79294,G79295,G79296,G79297,G79298,G79299,G79300,
       G79301,G79302,G79303,G79304,G79305,G79306,G79307,G79308,G79309,G79310,G79311,G79312,G79313,G79314,G79315,G79316,G79317,G79318,G79319,G79320,
       G79321,G79322,G79323,G79324,G79325,G79326,G79327,G79328,G79329,G79330,G79331,G79332,G79333,G79334,G79335,G79336,G79337,G79338,G79339,G79340,
       G79341,G79342,G79343,G79344,G79345,G79346,G79347,G79348,G79349,G79350,G79351,G79352,G79353,G79354,G79355,G79356,G79357,G79358,G79359,G79360,
       G79361,G79362,G79363,G79364,G79365,G79366,G79367,G79368,G79369,G79370,G79371,G79372,G79373,G79374,G79375,G79376,G79377,G79378,G79379,G79380,
       G79381,G79382,G79383,G79384,G79385,G79386,G79387,G79388,G79389,G79390,G79391,G79392,G79393,G79394,G79395,G79396,G79397,G79398,G79399,G79400,
       G79401,G79402,G79403,G79404,G79405,G79406,G79407,G79408,G79409,G79410,G79411,G79412,G79413,G79414,G79415,G79416,G79417,G79418,G79419,G79420,
       G79421,G79422,G79423,G79424,G79425,G79426,G79427,G79428,G79429,G79430,G79431,G79432,G79433,G79434,G79435,G79436,G79437,G79438,G79439,G79440,
       G79441,G79442,G79443,G79444,G79445,G79446,G79447,G79448,G79449,G79450,G79451,G79452,G79453,G79454,G79455,G79456,G79457,G79458,G79459,G79460,
       G79461,G79462,G79463,G79464,G79465,G79466,G79467,G79468,G79469,G79470,G79471,G79472,G79473,G79474,G79475,G79476,G79477,G79478,G79479,G79480,
       G79481,G79482,G79483,G79484,G79485,G79486,G79487,G79488,G79489,G79490,G79491,G79492,G79493,G79494,G79495,G79496,G79497,G79498,G79499,G79500,
       G79501,G79502,G79503,G79504,G79505,G79506,G79507,G79508,G79509,G79510,G79511,G79512,G79513,G79514,G79515,G79516,G79517,G79518,G79519,G79520,
       G79521,G79522,G79523,G79524,G79525,G79526,G79527,G79528,G79529,G79530,G79531,G79532,G79533,G79534,G79535,G79536,G79537,G79538,G79539,G79540,
       G79541,G79542,G79543,G79544,G79545,G79546,G79547,G79548,G79549,G79550,G79551,G79552,G79553,G79554,G79555,G79556,G79557,G79558,G79559,G79560,
       G79561,G79562,G79563,G79564,G79565,G79566,G79567,G79568,G79569,G79570,G79571,G79572,G79573,G79574,G79575,G79576,G79577,G79578,G79579,G79580,
       G79581,G79582,G79583,G79584,G79585,G79586,G79587,G79588,G79589,G79590,G79591,G79592,G79593,G79594,G79595,G79596,G79597,G79598,G79599,G79600,
       G79601,G79602,G79603,G79604,G79605,G79606,G79607,G79608,G79609,G79610,G79611,G79612,G79613,G79614,G79615,G79616,G79617,G79618,G79619,G79620,
       G79621,G79622,G79623,G79624,G79625,G79626,G79627,G79628,G79629,G79630,G79631,G79632,G79633,G79634,G79635,G79636,G79637,G79638,G79639,G79640,
       G79641,G79642,G79643,G79644,G79645,G79646,G79647,G79648,G79649,G79650,G79651,G79652,G79653,G79654,G79655,G79656,G79657,G79658,G79659,G79660,
       G79661,G79662,G79663,G79664,G79665,G79666,G79667,G79668,G79669,G79670,G79671,G79672,G79673,G79674,G79675,G79676,G79677,G79678,G79679,G79680,
       G79681,G79682,G79683,G79684,G79685,G79686,G79687,G79688,G79689,G79690,G79691,G79692,G79693,G79694,G79695,G79696,G79697,G79698,G79699,G79700,
       G79701,G79702,G79703,G79704,G79705,G79706,G79707,G79708,G79709,G79710,G79711,G79712,G79713,G79714,G79715,G79716,G79717,G79718,G79719,G79720,
       G79721,G79722,G79723,G79724,G79725,G79726,G79727,G79728,G79729,G79730,G79731,G79732,G79733,G79734,G79735,G79736,G79737,G79738,G79739,G79740,
       G79741,G79742,G79743,G79744,G79745,G79746,G79747,G79748,G79749,G79750,G79751,G79752,G79753,G79754,G79755,G79756,G79757,G79758,G79759,G79760,
       G79761,G79762,G79763,G79764,G79765,G79766,G79767,G79768,G79769,G79770,G79771,G79772,G79773,G79774,G79775,G79776,G79777,G79778,G79779,G79780,
       G79781,G79782,G79783,G79784,G79785,G79786,G79787,G79788,G79789,G79790,G79791,G79792,G79793,G79794,G79795,G79796,G79797,G79798,G79799,G79800,
       G79801,G79802,G79803,G79804,G79805,G79806,G79807,G79808,G79809,G79810,G79811,G79812,G79813,G79814,G79815,G79816,G79817,G79818,G79819,G79820,
       G79821,G79822,G79823,G79824,G79825,G79826,G79827,G79828,G79829,G79830,G79831,G79832,G79833,G79834,G79835,G79836,G79837,G79838,G79839,G79840,
       G79841,G79842,G79843,G79844,G79845,G79846,G79847,G79848,G79849,G79850,G79851,G79852,G79853,G79854,G79855,G79856,G79857,G79858,G79859,G79860,
       G79861,G79862,G79863,G79864,G79865,G79866,G79867,G79868,G79869,G79870,G79871,G79872,G79873,G79874,G79875,G79876,G79877,G79878,G79879,G79880,
       G79881,G79882,G79883,G79884,G79885,G79886,G79887,G79888,G79889,G79890,G79891,G79892,G79893,G79894,G79895,G79896,G79897,G79898,G79899,G79900,
       G79901,G79902,G79903,G79904,G79905,G79906,G79907,G79908,G79909,G79910,G79911,G79912,G79913,G79914,G79915,G79916,G79917,G79918,G79919,G79920,
       G79921,G79922,G79923,G79924,G79925,G79926,G79927,G79928,G79929,G79930,G79931,G79932,G79933,G79934,G79935,G79936,G79937,G79938,G79939,G79940,
       G79941,G79942,G79943,G79944,G79945,G79946,G79947,G79948,G79949,G79950,G79951,G79952,G79953,G79954,G79955,G79956,G79957,G79958,G79959,G79960,
       G79961,G79962,G79963,G79964,G79965,G79966,G79967,G79968,G79969,G79970,G79971,G79972,G79973,G79974,G79975,G79976,G79977,G79978,G79979,G79980,
       G79981,G79982,G79983,G79984,G79985,G79986,G79987,G79988,G79989,G79990,G79991,G79992,G79993,G79994,G79995,G79996,G79997,G79998,G79999,G80000,
       G80001,G80002,G80003,G80004,G80005,G80006,G80007,G80008,G80009,G80010,G80011,G80012,G80013,G80014,G80015,G80016,G80017,G80018,G80019,G80020,
       G80021,G80022,G80023,G80024,G80025,G80026,G80027,G80028,G80029,G80030,G80031,G80032,G80033,G80034,G80035,G80036,G80037,G80038,G80039,G80040,
       G80041,G80042,G80043,G80044,G80045,G80046,G80047,G80048,G80049,G80050,G80051,G80052,G80053,G80054,G80055,G80056,G80057,G80058,G80059,G80060,
       G80061,G80062,G80063,G80064,G80065,G80066,G80067,G80068,G80069,G80070,G80071,G80072,G80073,G80074,G80075,G80076,G80077,G80078,G80079,G80080,
       G80081,G80082,G80083,G80084,G80085,G80086,G80087,G80088,G80089,G80090,G80091,G80092,G80093,G80094,G80095,G80096,G80097,G80098,G80099,G80100,
       G80101,G80102,G80103,G80104,G80105,G80106,G80107,G80108,G80109,G80110,G80111,G80112,G80113,G80114,G80115,G80116,G80117,G80118,G80119,G80120,
       G80121,G80122,G80123,G80124,G80125,G80126,G80127,G80128,G80129,G80130,G80131,G80132,G80133,G80134,G80135,G80136,G80137,G80138,G80139,G80140,
       G80141,G80142,G80143,G80144,G80145,G80146,G80147,G80148,G80149,G80150,G80151,G80152,G80153,G80154,G80155,G80156,G80157,G80158,G80159,G80160,
       G80161,G80162,G80163,G80164,G80165,G80166,G80167,G80168,G80169,G80170,G80171,G80172,G80173,G80174,G80175,G80176,G80177,G80178,G80179,G80180,
       G80181,G80182,G80183,G80184,G80185,G80186,G80187,G80188,G80189,G80190,G80191,G80192,G80193,G80194,G80195,G80196,G80197,G80198,G80199,G80200,
       G80201,G80202,G80203,G80204,G80205,G80206,G80207,G80208,G80209,G80210,G80211,G80212,G80213,G80214,G80215,G80216,G80217,G80218,G80219,G80220,
       G80221,G80222,G80223,G80224,G80225,G80226,G80227,G80228,G80229,G80230,G80231,G80232,G80233,G80234,G80235,G80236,G80237,G80238,G80239,G80240,
       G80241,G80242,G80243,G80244,G80245,G80246,G80247,G80248,G80249,G80250,G80251,G80252,G80253,G80254,G80255,G80256,G80257,G80258,G80259,G80260,
       G80261,G80262,G80263,G80264,G80265,G80266,G80267,G80268,G80269,G80270,G80271,G80272,G80273,G80274,G80275,G80276,G80277,G80278,G80279,G80280,
       G80281,G80282,G80283,G80284,G80285,G80286,G80287,G80288,G80289,G80290,G80291,G80292,G80293,G80294,G80295,G80296,G80297,G80298,G80299,G80300,
       G80301,G80302,G80303,G80304,G80305,G80306,G80307,G80308,G80309,G80310,G80311,G80312,G80313,G80314,G80315,G80316,G80317,G80318,G80319,G80320,
       G80321,G80322,G80323,G80324,G80325,G80326,G80327,G80328,G80329,G80330,G80331,G80332,G80333,G80334,G80335,G80336,G80337,G80338,G80339,G80340,
       G80341,G80342,G80343,G80344,G80345,G80346,G80347,G80348,G80349,G80350,G80351,G80352,G80353,G80354,G80355,G80356,G80357,G80358,G80359,G80360,
       G80361,G80362,G80363,G80364,G80365,G80366,G80367,G80368,G80369,G80370,G80371,G80372,G80373,G80374,G80375,G80376,G80377,G80378,G80379,G80380,
       G80381,G80382,G80383,G80384,G80385,G80386,G80387,G80388,G80389,G80390,G80391,G80392,G80393,G80394,G80395,G80396,G80397,G80398,G80399,G80400,
       G80401,G80402,G80403,G80404,G80405,G80406,G80407,G80408,G80409,G80410,G80411,G80412,G80413,G80414,G80415,G80416,G80417,G80418,G80419,G80420,
       G80421,G80422,G80423,G80424,G80425,G80426,G80427,G80428,G80429,G80430,G80431,G80432,G80433,G80434,G80435,G80436,G80437,G80438,G80439,G80440,
       G80441,G80442,G80443,G80444,G80445,G80446,G80447,G80448,G80449,G80450,G80451,G80452,G80453,G80454,G80455,G80456,G80457,G80458,G80459,G80460,
       G80461,G80462,G80463,G80464,G80465,G80466,G80467,G80468,G80469,G80470,G80471,G80472,G80473,G80474,G80475,G80476,G80477,G80478,G80479,G80480,
       G80481,G80482,G80483,G80484,G80485,G80486,G80487,G80488,G80489,G80490,G80491,G80492,G80493,G80494,G80495,G80496,G80497,G80498,G80499,G80500,
       G80501,G80502,G80503,G80504,G80505,G80506,G80507,G80508,G80509,G80510,G80511,G80512,G80513,G80514,G80515,G80516,G80517,G80518,G80519,G80520,
       G80521,G80522,G80523,G80524,G80525,G80526,G80527,G80528,G80529,G80530,G80531,G80532,G80533,G80534,G80535,G80536,G80537,G80538,G80539,G80540,
       G80541,G80542,G80543,G80544,G80545,G80546,G80547,G80548,G80549,G80550,G80551,G80552,G80553,G80554,G80555,G80556,G80557,G80558,G80559,G80560,
       G80561,G80562,G80563,G80564,G80565,G80566,G80567,G80568,G80569,G80570,G80571,G80572,G80573,G80574,G80575,G80576,G80577,G80578,G80579,G80580,
       G80581,G80582,G80583,G80584,G80585,G80586,G80587,G80588,G80589,G80590,G80591,G80592,G80593,G80594,G80595,G80596,G80597,G80598,G80599,G80600,
       G80601,G80602,G80603,G80604,G80605,G80606,G80607,G80608,G80609,G80610,G80611,G80612,G80613,G80614,G80615,G80616,G80617,G80618,G80619,G80620,
       G80621,G80622,G80623,G80624,G80625,G80626,G80627,G80628,G80629,G80630,G80631,G80632,G80633,G80634,G80635,G80636,G80637,G80638,G80639,G80640,
       G80641,G80642,G80643,G80644,G80645,G80646,G80647,G80648,G80649,G80650,G80651,G80652,G80653,G80654,G80655,G80656,G80657,G80658,G80659,G80660,
       G80661,G80662,G80663,G80664,G80665,G80666,G80667,G80668,G80669,G80670,G80671,G80672,G80673,G80674,G80675,G80676,G80677,G80678,G80679,G80680,
       G80681,G80682,G80683,G80684,G80685,G80686,G80687,G80688,G80689,G80690,G80691,G80692,G80693,G80694,G80695,G80696,G80697,G80698,G80699,G80700,
       G80701,G80702,G80703,G80704,G80705,G80706,G80707,G80708,G80709,G80710,G80711,G80712,G80713,G80714,G80715,G80716,G80717,G80718,G80719,G80720,
       G80721,G80722,G80723,G80724,G80725,G80726,G80727,G80728,G80729,G80730,G80731,G80732,G80733,G80734,G80735,G80736,G80737,G80738,G80739,G80740,
       G80741,G80742,G80743,G80744,G80745,G80746,G80747,G80748,G80749,G80750,G80751,G80752,G80753,G80754,G80755,G80756,G80757,G80758,G80759,G80760,
       G80761,G80762,G80763,G80764,G80765,G80766,G80767,G80768,G80769,G80770,G80771,G80772,G80773,G80774,G80775,G80776,G80777,G80778,G80779,G80780,
       G80781,G80782,G80783,G80784,G80785,G80786,G80787,G80788,G80789,G80790,G80791,G80792,G80793,G80794,G80795,G80796,G80797,G80798,G80799,G80800,
       G80801,G80802,G80803,G80804,G80805,G80806,G80807,G80808,G80809,G80810,G80811,G80812,G80813,G80814,G80815,G80816,G80817,G80818,G80819,G80820,
       G80821,G80822,G80823,G80824,G80825,G80826,G80827,G80828,G80829,G80830,G80831,G80832,G80833,G80834,G80835,G80836,G80837,G80838,G80839,G80840,
       G80841,G80842,G80843,G80844,G80845,G80846,G80847,G80848,G80849,G80850,G80851,G80852,G80853,G80854,G80855,G80856,G80857,G80858,G80859,G80860,
       G80861,G80862,G80863,G80864,G80865,G80866,G80867,G80868,G80869,G80870,G80871,G80872,G80873,G80874,G80875,G80876,G80877,G80878,G80879,G80880,
       G80881,G80882,G80883,G80884,G80885,G80886,G80887,G80888,G80889,G80890,G80891,G80892,G80893,G80894,G80895,G80896,G80897,G80898,G80899,G80900,
       G80901,G80902,G80903,G80904,G80905,G80906,G80907,G80908,G80909,G80910,G80911,G80912,G80913,G80914,G80915,G80916,G80917,G80918,G80919,G80920,
       G80921,G80922,G80923,G80924,G80925,G80926,G80927,G80928,G80929,G80930,G80931,G80932,G80933,G80934,G80935,G80936,G80937,G80938,G80939,G80940,
       G80941,G80942,G80943,G80944,G80945,G80946,G80947,G80948,G80949,G80950,G80951,G80952,G80953,G80954,G80955,G80956,G80957,G80958,G80959,G80960,
       G80961,G80962,G80963,G80964,G80965,G80966,G80967,G80968,G80969,G80970,G80971,G80972,G80973,G80974,G80975,G80976,G80977,G80978,G80979,G80980,
       G80981,G80982,G80983,G80984,G80985,G80986,G80987,G80988,G80989,G80990,G80991,G80992,G80993,G80994,G80995,G80996,G80997,G80998,G80999,G81000,
       G81001,G81002,G81003,G81004,G81005,G81006,G81007,G81008,G81009,G81010,G81011,G81012,G81013,G81014,G81015,G81016,G81017,G81018,G81019,G81020,
       G81021,G81022,G81023,G81024,G81025,G81026,G81027,G81028,G81029,G81030,G81031,G81032,G81033,G81034,G81035,G81036,G81037,G81038,G81039,G81040,
       G81041,G81042,G81043,G81044,G81045,G81046,G81047,G81048,G81049,G81050,G81051,G81052,G81053,G81054,G81055,G81056,G81057,G81058,G81059,G81060,
       G81061,G81062,G81063,G81064,G81065,G81066,G81067,G81068,G81069,G81070,G81071,G81072,G81073,G81074,G81075,G81076,G81077,G81078,G81079,G81080,
       G81081,G81082,G81083;

  buf GNAME80(G80,G39);
  buf GNAME81(G81,G38);
  buf GNAME82(G82,G37);
  buf GNAME83(G83,G36);
  buf GNAME84(G84,G35);
  buf GNAME85(G85,G34);
  buf GNAME86(G86,G33);
  buf GNAME87(G87,G32);
  buf GNAME88(G88,G31);
  buf GNAME89(G89,G30);
  buf GNAME90(G90,G29);
  buf GNAME91(G91,G28);
  buf GNAME92(G92,G27);
  buf GNAME93(G93,G7);
  buf GNAME94(G94,G8);
  buf GNAME95(G95,G9);
  buf GNAME96(G96,G10);
  buf GNAME97(G97,G11);
  buf GNAME98(G98,G12);
  buf GNAME99(G99,G13);
  buf GNAME100(G100,G14);
  buf GNAME101(G101,G26);
  buf GNAME102(G102,G1);
  buf GNAME103(G103,G2);
  buf GNAME104(G104,G3);
  buf GNAME105(G105,G4);
  buf GNAME106(G106,G5);
  buf GNAME107(G107,G6);
  buf GNAME108(G108,G25);
  buf GNAME109(G109,G24);
  buf GNAME110(G110,G23);
  buf GNAME112(G112,G626);
  buf GNAME114(G114,G8670);
  buf GNAME116(G116,G5218);
  buf GNAME118(G118,G80198);
  buf GNAME120(G120,G80666);
  buf GNAME122(G122,G80718);
  buf GNAME124(G124,G57344);
  buf GNAME126(G126,G57565);
  buf GNAME128(G128,G34594);
  buf GNAME130(G130,G34360);
  buf GNAME132(G132,G11490);
  buf GNAME134(G134,G11468);
  buf GNAME136(G136,G11447);
  buf GNAME138(G138,G11426);
  buf GNAME140(G140,G11405);
  buf GNAME142(G142,G11384);
  buf GNAME144(G144,G11363);
  buf GNAME146(G146,G11342);
  not GNAME387(G387,G389);
  not GNAME388(G388,G108);
  or GNAME389(G389,G494,G388);
  not GNAME390(G390,G392);
  not GNAME391(G391,G611);
  or GNAME392(G392,G624,G391);
  nor GNAME393(G393,G459,G507);
  nor GNAME394(G394,G507,G520);
  nor GNAME395(G395,G633,G467);
  nor GNAME396(G396,G634,G468);
  nor GNAME397(G397,G629,G475);
  nor GNAME398(G398,G633,G468);
  nor GNAME399(G399,G635,G468);
  nor GNAME400(G400,G629,G468);
  nor GNAME401(G401,G634,G467);
  nor GNAME402(G402,G632,G467);
  nor GNAME403(G403,G628,G467);
  nor GNAME404(G404,G631,G469);
  nor GNAME405(G405,G630,G469);
  nor GNAME406(G406,G635,G469);
  nor GNAME407(G407,G628,G469);
  nor GNAME408(G408,G631,G470);
  nor GNAME409(G409,G630,G470);
  nor GNAME410(G410,G632,G470);
  nor GNAME411(G411,G629,G470);
  nor GNAME412(G412,G631,G471);
  nor GNAME413(G413,G630,G471);
  nor GNAME414(G414,G632,G471);
  nor GNAME415(G415,G628,G471);
  nor GNAME416(G416,G631,G472);
  nor GNAME417(G417,G630,G472);
  nor GNAME418(G418,G635,G472);
  nor GNAME419(G419,G628,G472);
  nor GNAME420(G420,G631,G473);
  nor GNAME421(G421,G630,G473);
  nor GNAME422(G422,G635,G473);
  nor GNAME423(G423,G629,G473);
  nor GNAME424(G424,G631,G474);
  nor GNAME425(G425,G630,G474);
  nor GNAME426(G426,G632,G474);
  nor GNAME427(G427,G629,G474);
  nor GNAME428(G428,G631,G475);
  nor GNAME429(G429,G630,G475);
  nor GNAME430(G430,G632,G475);
  nor GNAME431(G431,G634,G476);
  nor GNAME432(G432,G633,G476);
  nor GNAME433(G433,G632,G476);
  nor GNAME434(G434,G628,G476);
  nor GNAME435(G435,G629,G477);
  nor GNAME436(G436,G635,G477);
  nor GNAME437(G437,G635,G482);
  nor GNAME438(G438,G477,G634);
  nor GNAME439(G439,G477,G633);
  nor GNAME440(G440,G482,G634);
  nor GNAME441(G441,G482,G633);
  nor GNAME442(G442,G482,G629);
  nor GNAME443(G443,G633,G478);
  nor GNAME444(G444,G628,G478);
  nor GNAME445(G445,G633,G480);
  nor GNAME446(G446,G635,G478);
  nor GNAME447(G447,G634,G480);
  nor GNAME448(G448,G632,G480);
  nor GNAME449(G449,G634,G481);
  nor GNAME450(G450,G628,G481);
  nor GNAME451(G451,G629,G480);
  nor GNAME452(G452,G633,G481);
  nor GNAME453(G453,G634,G478);
  nor GNAME454(G454,G635,G481);
  not GNAME455(G455,G572);
  not GNAME456(G456,G559);
  not GNAME457(G457,G546);
  not GNAME458(G458,G533);
  not GNAME459(G459,G520);
  and GNAME460(G460,G455,G598,G456);
  and GNAME461(G461,G598,G456,G572);
  and GNAME462(G462,G598,G455,G559);
  and GNAME463(G463,G572,G585,G559);
  nand GNAME464(G464,G546,G458);
  nand GNAME465(G465,G533,G457);
  nand GNAME466(G466,G533,G546);
  nand GNAME467(G467,G484,G460);
  nand GNAME468(G468,G483,G460);
  nand GNAME469(G469,G484,G462);
  nand GNAME470(G470,G484,G461);
  nand GNAME471(G471,G462,G483);
  nand GNAME472(G472,G462,G393);
  nand GNAME473(G473,G462,G394);
  nand GNAME474(G474,G461,G483);
  nand GNAME475(G475,G461,G393);
  nand GNAME476(G476,G461,G394);
  nand GNAME477(G477,G394,G460);
  nand GNAME478(G478,G463,G484);
  nand GNAME479(G479,G458,G457);
  nand GNAME480(G480,G463,G393);
  nand GNAME481(G481,G463,G394);
  nand GNAME482(G482,G460,G393);
  and GNAME483(G483,G507,G520);
  and GNAME484(G484,G507,G459);
  dff DFF_493(CK,G492,G108);
  and GNAME494(G494,G492,G495);
  nand GNAME495(G495,G80,G497);
  buf GNAME496(G496,G492);
  buf GNAME497(G497,G487);
  dff DFF_506(CK,G505,G104);
  and GNAME507(G507,G505,G508);
  nand GNAME508(G508,G80,G510);
  buf GNAME509(G509,G505);
  buf GNAME510(G510,G500);
  dff DFF_519(CK,G518,G105);
  and GNAME520(G520,G518,G521);
  nand GNAME521(G521,G80,G523);
  buf GNAME522(G522,G518);
  buf GNAME523(G523,G513);
  dff DFF_532(CK,G531,G106);
  and GNAME533(G533,G531,G534);
  nand GNAME534(G534,G80,G536);
  buf GNAME535(G535,G531);
  buf GNAME536(G536,G526);
  dff DFF_545(CK,G544,G107);
  and GNAME546(G546,G544,G547);
  nand GNAME547(G547,G80,G549);
  buf GNAME548(G548,G544);
  buf GNAME549(G549,G539);
  dff DFF_558(CK,G557,G102);
  and GNAME559(G559,G557,G560);
  nand GNAME560(G560,G80,G562);
  buf GNAME561(G561,G557);
  buf GNAME562(G562,G552);
  dff DFF_571(CK,G570,G103);
  and GNAME572(G572,G570,G573);
  nand GNAME573(G573,G80,G575);
  buf GNAME574(G574,G570);
  buf GNAME575(G575,G565);
  dff DFF_584(CK,G583,G387);
  and GNAME585(G585,G583,G586);
  nand GNAME586(G586,G80,G588);
  buf GNAME587(G587,G583);
  buf GNAME588(G588,G578);
  dff DFF_597(CK,G596,G390);
  and GNAME598(G598,G596,G599);
  nand GNAME599(G599,G80,G601);
  buf GNAME600(G600,G596);
  buf GNAME601(G601,G591);
  dff DFF_610(CK,G609,G585);
  and GNAME611(G611,G609,G612);
  nand GNAME612(G612,G80,G614);
  buf GNAME613(G613,G609);
  buf GNAME614(G614,G604);
  dff DFF_623(CK,G622,G101);
  and GNAME624(G624,G622,G625);
  nand GNAME625(G625,G80,G627);
  buf GNAME626(G626,G622);
  buf GNAME627(G627,G617);
  buf GNAME628(G628,G479);
  buf GNAME629(G629,G479);
  buf GNAME630(G630,G465);
  buf GNAME631(G631,G466);
  buf GNAME632(G632,G464);
  buf GNAME633(G633,G465);
  buf GNAME634(G634,G466);
  buf GNAME635(G635,G464);
  or GNAME1298(G1298,G1300,G1299);
  and GNAME1299(G1299,G93,G390);
  and GNAME1300(G1300,G1302,G1301);
  not GNAME1301(G1301,G390);
  dff DFF_1303(CK,G1302,G1298);
  and GNAME1304(G1304,G1302,G1305);
  nand GNAME1305(G1305,G80,G1307);
  buf GNAME1306(G1306,G1302);
  buf GNAME1307(G1307,G1289);
  or GNAME1319(G1319,G1321,G1320);
  and GNAME1320(G1320,G100,G390);
  and GNAME1321(G1321,G1323,G1322);
  not GNAME1322(G1322,G390);
  dff DFF_1324(CK,G1323,G1319);
  and GNAME1325(G1325,G1323,G1326);
  nand GNAME1326(G1326,G80,G1328);
  buf GNAME1327(G1327,G1323);
  buf GNAME1328(G1328,G1310);
  or GNAME1340(G1340,G1342,G1341);
  and GNAME1341(G1341,G99,G390);
  and GNAME1342(G1342,G1344,G1343);
  not GNAME1343(G1343,G390);
  dff DFF_1345(CK,G1344,G1340);
  and GNAME1346(G1346,G1344,G1347);
  nand GNAME1347(G1347,G80,G1349);
  buf GNAME1348(G1348,G1344);
  buf GNAME1349(G1349,G1331);
  or GNAME1361(G1361,G1363,G1362);
  and GNAME1362(G1362,G98,G390);
  and GNAME1363(G1363,G1365,G1364);
  not GNAME1364(G1364,G390);
  dff DFF_1366(CK,G1365,G1361);
  and GNAME1367(G1367,G1365,G1368);
  nand GNAME1368(G1368,G80,G1370);
  buf GNAME1369(G1369,G1365);
  buf GNAME1370(G1370,G1352);
  or GNAME1382(G1382,G1384,G1383);
  and GNAME1383(G1383,G97,G390);
  and GNAME1384(G1384,G1386,G1385);
  not GNAME1385(G1385,G390);
  dff DFF_1387(CK,G1386,G1382);
  and GNAME1388(G1388,G1386,G1389);
  nand GNAME1389(G1389,G80,G1391);
  buf GNAME1390(G1390,G1386);
  buf GNAME1391(G1391,G1373);
  or GNAME1403(G1403,G1405,G1404);
  and GNAME1404(G1404,G96,G390);
  and GNAME1405(G1405,G1407,G1406);
  not GNAME1406(G1406,G390);
  dff DFF_1408(CK,G1407,G1403);
  and GNAME1409(G1409,G1407,G1410);
  nand GNAME1410(G1410,G80,G1412);
  buf GNAME1411(G1411,G1407);
  buf GNAME1412(G1412,G1394);
  or GNAME1424(G1424,G1426,G1425);
  and GNAME1425(G1425,G95,G390);
  and GNAME1426(G1426,G1428,G1427);
  not GNAME1427(G1427,G390);
  dff DFF_1429(CK,G1428,G1424);
  and GNAME1430(G1430,G1428,G1431);
  nand GNAME1431(G1431,G80,G1433);
  buf GNAME1432(G1432,G1428);
  buf GNAME1433(G1433,G1415);
  or GNAME1445(G1445,G1447,G1446);
  and GNAME1446(G1446,G94,G390);
  and GNAME1447(G1447,G1449,G1448);
  not GNAME1448(G1448,G390);
  dff DFF_1450(CK,G1449,G1445);
  and GNAME1451(G1451,G1449,G1452);
  nand GNAME1452(G1452,G80,G1454);
  buf GNAME1453(G1453,G1449);
  buf GNAME1454(G1454,G1436);
  or GNAME1506(G1506,G1508,G1507);
  and GNAME1507(G1507,G11522,G435);
  and GNAME1508(G1508,G1510,G1509);
  not GNAME1509(G1509,G435);
  dff DFF_1511(CK,G1510,G1506);
  and GNAME1512(G1512,G1510,G1513);
  nand GNAME1513(G1513,G80,G1515);
  buf GNAME1514(G1514,G1510);
  buf GNAME1515(G1515,G1497);
  or GNAME1527(G1527,G1529,G1528);
  and GNAME1528(G1528,G11521,G435);
  and GNAME1529(G1529,G1531,G1530);
  not GNAME1530(G1530,G435);
  dff DFF_1532(CK,G1531,G1527);
  and GNAME1533(G1533,G1531,G1534);
  nand GNAME1534(G1534,G80,G1536);
  buf GNAME1535(G1535,G1531);
  buf GNAME1536(G1536,G1518);
  or GNAME1548(G1548,G1550,G1549);
  and GNAME1549(G1549,G11520,G435);
  and GNAME1550(G1550,G1552,G1551);
  not GNAME1551(G1551,G435);
  dff DFF_1553(CK,G1552,G1548);
  and GNAME1554(G1554,G1552,G1555);
  nand GNAME1555(G1555,G80,G1557);
  buf GNAME1556(G1556,G1552);
  buf GNAME1557(G1557,G1539);
  or GNAME1569(G1569,G1571,G1570);
  and GNAME1570(G1570,G11519,G435);
  and GNAME1571(G1571,G1573,G1572);
  not GNAME1572(G1572,G435);
  dff DFF_1574(CK,G1573,G1569);
  and GNAME1575(G1575,G1573,G1576);
  nand GNAME1576(G1576,G80,G1578);
  buf GNAME1577(G1577,G1573);
  buf GNAME1578(G1578,G1560);
  or GNAME1590(G1590,G1592,G1591);
  and GNAME1591(G1591,G11518,G435);
  and GNAME1592(G1592,G1594,G1593);
  not GNAME1593(G1593,G435);
  dff DFF_1595(CK,G1594,G1590);
  and GNAME1596(G1596,G1594,G1597);
  nand GNAME1597(G1597,G80,G1599);
  buf GNAME1598(G1598,G1594);
  buf GNAME1599(G1599,G1581);
  or GNAME1611(G1611,G1613,G1612);
  and GNAME1612(G1612,G11517,G435);
  and GNAME1613(G1613,G1615,G1614);
  not GNAME1614(G1614,G435);
  dff DFF_1616(CK,G1615,G1611);
  and GNAME1617(G1617,G1615,G1618);
  nand GNAME1618(G1618,G80,G1620);
  buf GNAME1619(G1619,G1615);
  buf GNAME1620(G1620,G1602);
  or GNAME1632(G1632,G1634,G1633);
  and GNAME1633(G1633,G11516,G435);
  and GNAME1634(G1634,G1636,G1635);
  not GNAME1635(G1635,G435);
  dff DFF_1637(CK,G1636,G1632);
  and GNAME1638(G1638,G1636,G1639);
  nand GNAME1639(G1639,G80,G1641);
  buf GNAME1640(G1640,G1636);
  buf GNAME1641(G1641,G1623);
  or GNAME1653(G1653,G1655,G1654);
  and GNAME1654(G1654,G11515,G435);
  and GNAME1655(G1655,G1657,G1656);
  not GNAME1656(G1656,G435);
  dff DFF_1658(CK,G1657,G1653);
  and GNAME1659(G1659,G1657,G1660);
  nand GNAME1660(G1660,G80,G1662);
  buf GNAME1661(G1661,G1657);
  buf GNAME1662(G1662,G1644);
  or GNAME1714(G1714,G1716,G1715);
  and GNAME1715(G1715,G11546,G436);
  and GNAME1716(G1716,G1718,G1717);
  not GNAME1717(G1717,G436);
  dff DFF_1719(CK,G1718,G1714);
  and GNAME1720(G1720,G1718,G1721);
  nand GNAME1721(G1721,G80,G1723);
  buf GNAME1722(G1722,G1718);
  buf GNAME1723(G1723,G1705);
  or GNAME1735(G1735,G1737,G1736);
  and GNAME1736(G1736,G11545,G436);
  and GNAME1737(G1737,G1739,G1738);
  not GNAME1738(G1738,G436);
  dff DFF_1740(CK,G1739,G1735);
  and GNAME1741(G1741,G1739,G1742);
  nand GNAME1742(G1742,G80,G1744);
  buf GNAME1743(G1743,G1739);
  buf GNAME1744(G1744,G1726);
  or GNAME1756(G1756,G1758,G1757);
  and GNAME1757(G1757,G11544,G436);
  and GNAME1758(G1758,G1760,G1759);
  not GNAME1759(G1759,G436);
  dff DFF_1761(CK,G1760,G1756);
  and GNAME1762(G1762,G1760,G1763);
  nand GNAME1763(G1763,G80,G1765);
  buf GNAME1764(G1764,G1760);
  buf GNAME1765(G1765,G1747);
  or GNAME1777(G1777,G1779,G1778);
  and GNAME1778(G1778,G11543,G436);
  and GNAME1779(G1779,G1781,G1780);
  not GNAME1780(G1780,G436);
  dff DFF_1782(CK,G1781,G1777);
  and GNAME1783(G1783,G1781,G1784);
  nand GNAME1784(G1784,G80,G1786);
  buf GNAME1785(G1785,G1781);
  buf GNAME1786(G1786,G1768);
  or GNAME1798(G1798,G1800,G1799);
  and GNAME1799(G1799,G11542,G436);
  and GNAME1800(G1800,G1802,G1801);
  not GNAME1801(G1801,G436);
  dff DFF_1803(CK,G1802,G1798);
  and GNAME1804(G1804,G1802,G1805);
  nand GNAME1805(G1805,G80,G1807);
  buf GNAME1806(G1806,G1802);
  buf GNAME1807(G1807,G1789);
  or GNAME1819(G1819,G1821,G1820);
  and GNAME1820(G1820,G11541,G436);
  and GNAME1821(G1821,G1823,G1822);
  not GNAME1822(G1822,G436);
  dff DFF_1824(CK,G1823,G1819);
  and GNAME1825(G1825,G1823,G1826);
  nand GNAME1826(G1826,G80,G1828);
  buf GNAME1827(G1827,G1823);
  buf GNAME1828(G1828,G1810);
  or GNAME1840(G1840,G1842,G1841);
  and GNAME1841(G1841,G11540,G436);
  and GNAME1842(G1842,G1844,G1843);
  not GNAME1843(G1843,G436);
  dff DFF_1845(CK,G1844,G1840);
  and GNAME1846(G1846,G1844,G1847);
  nand GNAME1847(G1847,G80,G1849);
  buf GNAME1848(G1848,G1844);
  buf GNAME1849(G1849,G1831);
  or GNAME1861(G1861,G1863,G1862);
  and GNAME1862(G1862,G11539,G436);
  and GNAME1863(G1863,G1865,G1864);
  not GNAME1864(G1864,G436);
  dff DFF_1866(CK,G1865,G1861);
  and GNAME1867(G1867,G1865,G1868);
  nand GNAME1868(G1868,G80,G1870);
  buf GNAME1869(G1869,G1865);
  buf GNAME1870(G1870,G1852);
  or GNAME1922(G1922,G1924,G1923);
  and GNAME1923(G1923,G11546,G439);
  and GNAME1924(G1924,G1926,G1925);
  not GNAME1925(G1925,G439);
  dff DFF_1927(CK,G1926,G1922);
  and GNAME1928(G1928,G1926,G1929);
  nand GNAME1929(G1929,G80,G1931);
  buf GNAME1930(G1930,G1926);
  buf GNAME1931(G1931,G1913);
  or GNAME1943(G1943,G1945,G1944);
  and GNAME1944(G1944,G11545,G439);
  and GNAME1945(G1945,G1947,G1946);
  not GNAME1946(G1946,G439);
  dff DFF_1948(CK,G1947,G1943);
  and GNAME1949(G1949,G1947,G1950);
  nand GNAME1950(G1950,G80,G1952);
  buf GNAME1951(G1951,G1947);
  buf GNAME1952(G1952,G1934);
  or GNAME1964(G1964,G1966,G1965);
  and GNAME1965(G1965,G11544,G439);
  and GNAME1966(G1966,G1968,G1967);
  not GNAME1967(G1967,G439);
  dff DFF_1969(CK,G1968,G1964);
  and GNAME1970(G1970,G1968,G1971);
  nand GNAME1971(G1971,G80,G1973);
  buf GNAME1972(G1972,G1968);
  buf GNAME1973(G1973,G1955);
  or GNAME1985(G1985,G1987,G1986);
  and GNAME1986(G1986,G11543,G439);
  and GNAME1987(G1987,G1989,G1988);
  not GNAME1988(G1988,G439);
  dff DFF_1990(CK,G1989,G1985);
  and GNAME1991(G1991,G1989,G1992);
  nand GNAME1992(G1992,G80,G1994);
  buf GNAME1993(G1993,G1989);
  buf GNAME1994(G1994,G1976);
  or GNAME2006(G2006,G2008,G2007);
  and GNAME2007(G2007,G11542,G439);
  and GNAME2008(G2008,G2010,G2009);
  not GNAME2009(G2009,G439);
  dff DFF_2011(CK,G2010,G2006);
  and GNAME2012(G2012,G2010,G2013);
  nand GNAME2013(G2013,G80,G2015);
  buf GNAME2014(G2014,G2010);
  buf GNAME2015(G2015,G1997);
  or GNAME2027(G2027,G2029,G2028);
  and GNAME2028(G2028,G11541,G439);
  and GNAME2029(G2029,G2031,G2030);
  not GNAME2030(G2030,G439);
  dff DFF_2032(CK,G2031,G2027);
  and GNAME2033(G2033,G2031,G2034);
  nand GNAME2034(G2034,G80,G2036);
  buf GNAME2035(G2035,G2031);
  buf GNAME2036(G2036,G2018);
  or GNAME2048(G2048,G2050,G2049);
  and GNAME2049(G2049,G11540,G439);
  and GNAME2050(G2050,G2052,G2051);
  not GNAME2051(G2051,G439);
  dff DFF_2053(CK,G2052,G2048);
  and GNAME2054(G2054,G2052,G2055);
  nand GNAME2055(G2055,G80,G2057);
  buf GNAME2056(G2056,G2052);
  buf GNAME2057(G2057,G2039);
  or GNAME2069(G2069,G2071,G2070);
  and GNAME2070(G2070,G11539,G439);
  and GNAME2071(G2071,G2073,G2072);
  not GNAME2072(G2072,G439);
  dff DFF_2074(CK,G2073,G2069);
  and GNAME2075(G2075,G2073,G2076);
  nand GNAME2076(G2076,G80,G2078);
  buf GNAME2077(G2077,G2073);
  buf GNAME2078(G2078,G2060);
  or GNAME2130(G2130,G2132,G2131);
  and GNAME2131(G2131,G11546,G438);
  and GNAME2132(G2132,G2134,G2133);
  not GNAME2133(G2133,G438);
  dff DFF_2135(CK,G2134,G2130);
  and GNAME2136(G2136,G2134,G2137);
  nand GNAME2137(G2137,G80,G2139);
  buf GNAME2138(G2138,G2134);
  buf GNAME2139(G2139,G2121);
  or GNAME2151(G2151,G2153,G2152);
  and GNAME2152(G2152,G11545,G438);
  and GNAME2153(G2153,G2155,G2154);
  not GNAME2154(G2154,G438);
  dff DFF_2156(CK,G2155,G2151);
  and GNAME2157(G2157,G2155,G2158);
  nand GNAME2158(G2158,G80,G2160);
  buf GNAME2159(G2159,G2155);
  buf GNAME2160(G2160,G2142);
  or GNAME2172(G2172,G2174,G2173);
  and GNAME2173(G2173,G11544,G438);
  and GNAME2174(G2174,G2176,G2175);
  not GNAME2175(G2175,G438);
  dff DFF_2177(CK,G2176,G2172);
  and GNAME2178(G2178,G2176,G2179);
  nand GNAME2179(G2179,G80,G2181);
  buf GNAME2180(G2180,G2176);
  buf GNAME2181(G2181,G2163);
  or GNAME2193(G2193,G2195,G2194);
  and GNAME2194(G2194,G11543,G438);
  and GNAME2195(G2195,G2197,G2196);
  not GNAME2196(G2196,G438);
  dff DFF_2198(CK,G2197,G2193);
  and GNAME2199(G2199,G2197,G2200);
  nand GNAME2200(G2200,G80,G2202);
  buf GNAME2201(G2201,G2197);
  buf GNAME2202(G2202,G2184);
  or GNAME2214(G2214,G2216,G2215);
  and GNAME2215(G2215,G11542,G438);
  and GNAME2216(G2216,G2218,G2217);
  not GNAME2217(G2217,G438);
  dff DFF_2219(CK,G2218,G2214);
  and GNAME2220(G2220,G2218,G2221);
  nand GNAME2221(G2221,G80,G2223);
  buf GNAME2222(G2222,G2218);
  buf GNAME2223(G2223,G2205);
  or GNAME2235(G2235,G2237,G2236);
  and GNAME2236(G2236,G11541,G438);
  and GNAME2237(G2237,G2239,G2238);
  not GNAME2238(G2238,G438);
  dff DFF_2240(CK,G2239,G2235);
  and GNAME2241(G2241,G2239,G2242);
  nand GNAME2242(G2242,G80,G2244);
  buf GNAME2243(G2243,G2239);
  buf GNAME2244(G2244,G2226);
  or GNAME2256(G2256,G2258,G2257);
  and GNAME2257(G2257,G11540,G438);
  and GNAME2258(G2258,G2260,G2259);
  not GNAME2259(G2259,G438);
  dff DFF_2261(CK,G2260,G2256);
  and GNAME2262(G2262,G2260,G2263);
  nand GNAME2263(G2263,G80,G2265);
  buf GNAME2264(G2264,G2260);
  buf GNAME2265(G2265,G2247);
  or GNAME2277(G2277,G2279,G2278);
  and GNAME2278(G2278,G11539,G438);
  and GNAME2279(G2279,G2281,G2280);
  not GNAME2280(G2280,G438);
  dff DFF_2282(CK,G2281,G2277);
  and GNAME2283(G2283,G2281,G2284);
  nand GNAME2284(G2284,G80,G2286);
  buf GNAME2285(G2285,G2281);
  buf GNAME2286(G2286,G2268);
  or GNAME2338(G2338,G2340,G2339);
  and GNAME2339(G2339,G11546,G442);
  and GNAME2340(G2340,G2342,G2341);
  not GNAME2341(G2341,G442);
  dff DFF_2343(CK,G2342,G2338);
  and GNAME2344(G2344,G2342,G2345);
  nand GNAME2345(G2345,G80,G2347);
  buf GNAME2346(G2346,G2342);
  buf GNAME2347(G2347,G2329);
  or GNAME2359(G2359,G2361,G2360);
  and GNAME2360(G2360,G11545,G442);
  and GNAME2361(G2361,G2363,G2362);
  not GNAME2362(G2362,G442);
  dff DFF_2364(CK,G2363,G2359);
  and GNAME2365(G2365,G2363,G2366);
  nand GNAME2366(G2366,G80,G2368);
  buf GNAME2367(G2367,G2363);
  buf GNAME2368(G2368,G2350);
  or GNAME2380(G2380,G2382,G2381);
  and GNAME2381(G2381,G11544,G442);
  and GNAME2382(G2382,G2384,G2383);
  not GNAME2383(G2383,G442);
  dff DFF_2385(CK,G2384,G2380);
  and GNAME2386(G2386,G2384,G2387);
  nand GNAME2387(G2387,G80,G2389);
  buf GNAME2388(G2388,G2384);
  buf GNAME2389(G2389,G2371);
  or GNAME2401(G2401,G2403,G2402);
  and GNAME2402(G2402,G11543,G442);
  and GNAME2403(G2403,G2405,G2404);
  not GNAME2404(G2404,G442);
  dff DFF_2406(CK,G2405,G2401);
  and GNAME2407(G2407,G2405,G2408);
  nand GNAME2408(G2408,G80,G2410);
  buf GNAME2409(G2409,G2405);
  buf GNAME2410(G2410,G2392);
  or GNAME2422(G2422,G2424,G2423);
  and GNAME2423(G2423,G11542,G442);
  and GNAME2424(G2424,G2426,G2425);
  not GNAME2425(G2425,G442);
  dff DFF_2427(CK,G2426,G2422);
  and GNAME2428(G2428,G2426,G2429);
  nand GNAME2429(G2429,G80,G2431);
  buf GNAME2430(G2430,G2426);
  buf GNAME2431(G2431,G2413);
  or GNAME2443(G2443,G2445,G2444);
  and GNAME2444(G2444,G11541,G442);
  and GNAME2445(G2445,G2447,G2446);
  not GNAME2446(G2446,G442);
  dff DFF_2448(CK,G2447,G2443);
  and GNAME2449(G2449,G2447,G2450);
  nand GNAME2450(G2450,G80,G2452);
  buf GNAME2451(G2451,G2447);
  buf GNAME2452(G2452,G2434);
  or GNAME2464(G2464,G2466,G2465);
  and GNAME2465(G2465,G11540,G442);
  and GNAME2466(G2466,G2468,G2467);
  not GNAME2467(G2467,G442);
  dff DFF_2469(CK,G2468,G2464);
  and GNAME2470(G2470,G2468,G2471);
  nand GNAME2471(G2471,G80,G2473);
  buf GNAME2472(G2472,G2468);
  buf GNAME2473(G2473,G2455);
  or GNAME2485(G2485,G2487,G2486);
  and GNAME2486(G2486,G11539,G442);
  and GNAME2487(G2487,G2489,G2488);
  not GNAME2488(G2488,G442);
  dff DFF_2490(CK,G2489,G2485);
  and GNAME2491(G2491,G2489,G2492);
  nand GNAME2492(G2492,G80,G2494);
  buf GNAME2493(G2493,G2489);
  buf GNAME2494(G2494,G2476);
  or GNAME2546(G2546,G2548,G2547);
  and GNAME2547(G2547,G11546,G437);
  and GNAME2548(G2548,G2550,G2549);
  not GNAME2549(G2549,G437);
  dff DFF_2551(CK,G2550,G2546);
  and GNAME2552(G2552,G2550,G2553);
  nand GNAME2553(G2553,G80,G2555);
  buf GNAME2554(G2554,G2550);
  buf GNAME2555(G2555,G2537);
  or GNAME2567(G2567,G2569,G2568);
  and GNAME2568(G2568,G11545,G437);
  and GNAME2569(G2569,G2571,G2570);
  not GNAME2570(G2570,G437);
  dff DFF_2572(CK,G2571,G2567);
  and GNAME2573(G2573,G2571,G2574);
  nand GNAME2574(G2574,G80,G2576);
  buf GNAME2575(G2575,G2571);
  buf GNAME2576(G2576,G2558);
  or GNAME2588(G2588,G2590,G2589);
  and GNAME2589(G2589,G11544,G437);
  and GNAME2590(G2590,G2592,G2591);
  not GNAME2591(G2591,G437);
  dff DFF_2593(CK,G2592,G2588);
  and GNAME2594(G2594,G2592,G2595);
  nand GNAME2595(G2595,G80,G2597);
  buf GNAME2596(G2596,G2592);
  buf GNAME2597(G2597,G2579);
  or GNAME2609(G2609,G2611,G2610);
  and GNAME2610(G2610,G11543,G437);
  and GNAME2611(G2611,G2613,G2612);
  not GNAME2612(G2612,G437);
  dff DFF_2614(CK,G2613,G2609);
  and GNAME2615(G2615,G2613,G2616);
  nand GNAME2616(G2616,G80,G2618);
  buf GNAME2617(G2617,G2613);
  buf GNAME2618(G2618,G2600);
  or GNAME2630(G2630,G2632,G2631);
  and GNAME2631(G2631,G11542,G437);
  and GNAME2632(G2632,G2634,G2633);
  not GNAME2633(G2633,G437);
  dff DFF_2635(CK,G2634,G2630);
  and GNAME2636(G2636,G2634,G2637);
  nand GNAME2637(G2637,G80,G2639);
  buf GNAME2638(G2638,G2634);
  buf GNAME2639(G2639,G2621);
  or GNAME2651(G2651,G2653,G2652);
  and GNAME2652(G2652,G11541,G437);
  and GNAME2653(G2653,G2655,G2654);
  not GNAME2654(G2654,G437);
  dff DFF_2656(CK,G2655,G2651);
  and GNAME2657(G2657,G2655,G2658);
  nand GNAME2658(G2658,G80,G2660);
  buf GNAME2659(G2659,G2655);
  buf GNAME2660(G2660,G2642);
  or GNAME2672(G2672,G2674,G2673);
  and GNAME2673(G2673,G11540,G437);
  and GNAME2674(G2674,G2676,G2675);
  not GNAME2675(G2675,G437);
  dff DFF_2677(CK,G2676,G2672);
  and GNAME2678(G2678,G2676,G2679);
  nand GNAME2679(G2679,G80,G2681);
  buf GNAME2680(G2680,G2676);
  buf GNAME2681(G2681,G2663);
  or GNAME2693(G2693,G2695,G2694);
  and GNAME2694(G2694,G11539,G437);
  and GNAME2695(G2695,G2697,G2696);
  not GNAME2696(G2696,G437);
  dff DFF_2698(CK,G2697,G2693);
  and GNAME2699(G2699,G2697,G2700);
  nand GNAME2700(G2700,G80,G2702);
  buf GNAME2701(G2701,G2697);
  buf GNAME2702(G2702,G2684);
  or GNAME2754(G2754,G2756,G2755);
  and GNAME2755(G2755,G11546,G441);
  and GNAME2756(G2756,G2758,G2757);
  not GNAME2757(G2757,G441);
  dff DFF_2759(CK,G2758,G2754);
  and GNAME2760(G2760,G2758,G2761);
  nand GNAME2761(G2761,G80,G2763);
  buf GNAME2762(G2762,G2758);
  buf GNAME2763(G2763,G2745);
  or GNAME2775(G2775,G2777,G2776);
  and GNAME2776(G2776,G11545,G441);
  and GNAME2777(G2777,G2779,G2778);
  not GNAME2778(G2778,G441);
  dff DFF_2780(CK,G2779,G2775);
  and GNAME2781(G2781,G2779,G2782);
  nand GNAME2782(G2782,G80,G2784);
  buf GNAME2783(G2783,G2779);
  buf GNAME2784(G2784,G2766);
  or GNAME2796(G2796,G2798,G2797);
  and GNAME2797(G2797,G11544,G441);
  and GNAME2798(G2798,G2800,G2799);
  not GNAME2799(G2799,G441);
  dff DFF_2801(CK,G2800,G2796);
  and GNAME2802(G2802,G2800,G2803);
  nand GNAME2803(G2803,G80,G2805);
  buf GNAME2804(G2804,G2800);
  buf GNAME2805(G2805,G2787);
  or GNAME2817(G2817,G2819,G2818);
  and GNAME2818(G2818,G11543,G441);
  and GNAME2819(G2819,G2821,G2820);
  not GNAME2820(G2820,G441);
  dff DFF_2822(CK,G2821,G2817);
  and GNAME2823(G2823,G2821,G2824);
  nand GNAME2824(G2824,G80,G2826);
  buf GNAME2825(G2825,G2821);
  buf GNAME2826(G2826,G2808);
  or GNAME2838(G2838,G2840,G2839);
  and GNAME2839(G2839,G11542,G441);
  and GNAME2840(G2840,G2842,G2841);
  not GNAME2841(G2841,G441);
  dff DFF_2843(CK,G2842,G2838);
  and GNAME2844(G2844,G2842,G2845);
  nand GNAME2845(G2845,G80,G2847);
  buf GNAME2846(G2846,G2842);
  buf GNAME2847(G2847,G2829);
  or GNAME2859(G2859,G2861,G2860);
  and GNAME2860(G2860,G11541,G441);
  and GNAME2861(G2861,G2863,G2862);
  not GNAME2862(G2862,G441);
  dff DFF_2864(CK,G2863,G2859);
  and GNAME2865(G2865,G2863,G2866);
  nand GNAME2866(G2866,G80,G2868);
  buf GNAME2867(G2867,G2863);
  buf GNAME2868(G2868,G2850);
  or GNAME2880(G2880,G2882,G2881);
  and GNAME2881(G2881,G11540,G441);
  and GNAME2882(G2882,G2884,G2883);
  not GNAME2883(G2883,G441);
  dff DFF_2885(CK,G2884,G2880);
  and GNAME2886(G2886,G2884,G2887);
  nand GNAME2887(G2887,G80,G2889);
  buf GNAME2888(G2888,G2884);
  buf GNAME2889(G2889,G2871);
  or GNAME2901(G2901,G2903,G2902);
  and GNAME2902(G2902,G11539,G441);
  and GNAME2903(G2903,G2905,G2904);
  not GNAME2904(G2904,G441);
  dff DFF_2906(CK,G2905,G2901);
  and GNAME2907(G2907,G2905,G2908);
  nand GNAME2908(G2908,G80,G2910);
  buf GNAME2909(G2909,G2905);
  buf GNAME2910(G2910,G2892);
  or GNAME2962(G2962,G2964,G2963);
  and GNAME2963(G2963,G11546,G440);
  and GNAME2964(G2964,G2966,G2965);
  not GNAME2965(G2965,G440);
  dff DFF_2967(CK,G2966,G2962);
  and GNAME2968(G2968,G2966,G2969);
  nand GNAME2969(G2969,G80,G2971);
  buf GNAME2970(G2970,G2966);
  buf GNAME2971(G2971,G2953);
  or GNAME2983(G2983,G2985,G2984);
  and GNAME2984(G2984,G11545,G440);
  and GNAME2985(G2985,G2987,G2986);
  not GNAME2986(G2986,G440);
  dff DFF_2988(CK,G2987,G2983);
  and GNAME2989(G2989,G2987,G2990);
  nand GNAME2990(G2990,G80,G2992);
  buf GNAME2991(G2991,G2987);
  buf GNAME2992(G2992,G2974);
  or GNAME3004(G3004,G3006,G3005);
  and GNAME3005(G3005,G11544,G440);
  and GNAME3006(G3006,G3008,G3007);
  not GNAME3007(G3007,G440);
  dff DFF_3009(CK,G3008,G3004);
  and GNAME3010(G3010,G3008,G3011);
  nand GNAME3011(G3011,G80,G3013);
  buf GNAME3012(G3012,G3008);
  buf GNAME3013(G3013,G2995);
  or GNAME3025(G3025,G3027,G3026);
  and GNAME3026(G3026,G11543,G440);
  and GNAME3027(G3027,G3029,G3028);
  not GNAME3028(G3028,G440);
  dff DFF_3030(CK,G3029,G3025);
  and GNAME3031(G3031,G3029,G3032);
  nand GNAME3032(G3032,G80,G3034);
  buf GNAME3033(G3033,G3029);
  buf GNAME3034(G3034,G3016);
  or GNAME3046(G3046,G3048,G3047);
  and GNAME3047(G3047,G11542,G440);
  and GNAME3048(G3048,G3050,G3049);
  not GNAME3049(G3049,G440);
  dff DFF_3051(CK,G3050,G3046);
  and GNAME3052(G3052,G3050,G3053);
  nand GNAME3053(G3053,G80,G3055);
  buf GNAME3054(G3054,G3050);
  buf GNAME3055(G3055,G3037);
  or GNAME3067(G3067,G3069,G3068);
  and GNAME3068(G3068,G11541,G440);
  and GNAME3069(G3069,G3071,G3070);
  not GNAME3070(G3070,G440);
  dff DFF_3072(CK,G3071,G3067);
  and GNAME3073(G3073,G3071,G3074);
  nand GNAME3074(G3074,G80,G3076);
  buf GNAME3075(G3075,G3071);
  buf GNAME3076(G3076,G3058);
  or GNAME3088(G3088,G3090,G3089);
  and GNAME3089(G3089,G11540,G440);
  and GNAME3090(G3090,G3092,G3091);
  not GNAME3091(G3091,G440);
  dff DFF_3093(CK,G3092,G3088);
  and GNAME3094(G3094,G3092,G3095);
  nand GNAME3095(G3095,G80,G3097);
  buf GNAME3096(G3096,G3092);
  buf GNAME3097(G3097,G3079);
  or GNAME3109(G3109,G3111,G3110);
  and GNAME3110(G3110,G11539,G440);
  and GNAME3111(G3111,G3113,G3112);
  not GNAME3112(G3112,G440);
  dff DFF_3114(CK,G3113,G3109);
  and GNAME3115(G3115,G3113,G3116);
  nand GNAME3116(G3116,G80,G3118);
  buf GNAME3117(G3117,G3113);
  buf GNAME3118(G3118,G3100);
  or GNAME3170(G3170,G3172,G3171);
  and GNAME3171(G3171,G11546,G403);
  and GNAME3172(G3172,G3174,G3173);
  not GNAME3173(G3173,G403);
  dff DFF_3175(CK,G3174,G3170);
  and GNAME3176(G3176,G3174,G3177);
  nand GNAME3177(G3177,G80,G3179);
  buf GNAME3178(G3178,G3174);
  buf GNAME3179(G3179,G3161);
  or GNAME3191(G3191,G3193,G3192);
  and GNAME3192(G3192,G11545,G403);
  and GNAME3193(G3193,G3195,G3194);
  not GNAME3194(G3194,G403);
  dff DFF_3196(CK,G3195,G3191);
  and GNAME3197(G3197,G3195,G3198);
  nand GNAME3198(G3198,G80,G3200);
  buf GNAME3199(G3199,G3195);
  buf GNAME3200(G3200,G3182);
  or GNAME3212(G3212,G3214,G3213);
  and GNAME3213(G3213,G11544,G403);
  and GNAME3214(G3214,G3216,G3215);
  not GNAME3215(G3215,G403);
  dff DFF_3217(CK,G3216,G3212);
  and GNAME3218(G3218,G3216,G3219);
  nand GNAME3219(G3219,G80,G3221);
  buf GNAME3220(G3220,G3216);
  buf GNAME3221(G3221,G3203);
  or GNAME3233(G3233,G3235,G3234);
  and GNAME3234(G3234,G11543,G403);
  and GNAME3235(G3235,G3237,G3236);
  not GNAME3236(G3236,G403);
  dff DFF_3238(CK,G3237,G3233);
  and GNAME3239(G3239,G3237,G3240);
  nand GNAME3240(G3240,G80,G3242);
  buf GNAME3241(G3241,G3237);
  buf GNAME3242(G3242,G3224);
  or GNAME3254(G3254,G3256,G3255);
  and GNAME3255(G3255,G11542,G403);
  and GNAME3256(G3256,G3258,G3257);
  not GNAME3257(G3257,G403);
  dff DFF_3259(CK,G3258,G3254);
  and GNAME3260(G3260,G3258,G3261);
  nand GNAME3261(G3261,G80,G3263);
  buf GNAME3262(G3262,G3258);
  buf GNAME3263(G3263,G3245);
  or GNAME3275(G3275,G3277,G3276);
  and GNAME3276(G3276,G11541,G403);
  and GNAME3277(G3277,G3279,G3278);
  not GNAME3278(G3278,G403);
  dff DFF_3280(CK,G3279,G3275);
  and GNAME3281(G3281,G3279,G3282);
  nand GNAME3282(G3282,G80,G3284);
  buf GNAME3283(G3283,G3279);
  buf GNAME3284(G3284,G3266);
  or GNAME3296(G3296,G3298,G3297);
  and GNAME3297(G3297,G11540,G403);
  and GNAME3298(G3298,G3300,G3299);
  not GNAME3299(G3299,G403);
  dff DFF_3301(CK,G3300,G3296);
  and GNAME3302(G3302,G3300,G3303);
  nand GNAME3303(G3303,G80,G3305);
  buf GNAME3304(G3304,G3300);
  buf GNAME3305(G3305,G3287);
  or GNAME3317(G3317,G3319,G3318);
  and GNAME3318(G3318,G11539,G403);
  and GNAME3319(G3319,G3321,G3320);
  not GNAME3320(G3320,G403);
  dff DFF_3322(CK,G3321,G3317);
  and GNAME3323(G3323,G3321,G3324);
  nand GNAME3324(G3324,G80,G3326);
  buf GNAME3325(G3325,G3321);
  buf GNAME3326(G3326,G3308);
  or GNAME3378(G3378,G3380,G3379);
  and GNAME3379(G3379,G11546,G402);
  and GNAME3380(G3380,G3382,G3381);
  not GNAME3381(G3381,G402);
  dff DFF_3383(CK,G3382,G3378);
  and GNAME3384(G3384,G3382,G3385);
  nand GNAME3385(G3385,G80,G3387);
  buf GNAME3386(G3386,G3382);
  buf GNAME3387(G3387,G3369);
  or GNAME3399(G3399,G3401,G3400);
  and GNAME3400(G3400,G11545,G402);
  and GNAME3401(G3401,G3403,G3402);
  not GNAME3402(G3402,G402);
  dff DFF_3404(CK,G3403,G3399);
  and GNAME3405(G3405,G3403,G3406);
  nand GNAME3406(G3406,G80,G3408);
  buf GNAME3407(G3407,G3403);
  buf GNAME3408(G3408,G3390);
  or GNAME3420(G3420,G3422,G3421);
  and GNAME3421(G3421,G11544,G402);
  and GNAME3422(G3422,G3424,G3423);
  not GNAME3423(G3423,G402);
  dff DFF_3425(CK,G3424,G3420);
  and GNAME3426(G3426,G3424,G3427);
  nand GNAME3427(G3427,G80,G3429);
  buf GNAME3428(G3428,G3424);
  buf GNAME3429(G3429,G3411);
  or GNAME3441(G3441,G3443,G3442);
  and GNAME3442(G3442,G11543,G402);
  and GNAME3443(G3443,G3445,G3444);
  not GNAME3444(G3444,G402);
  dff DFF_3446(CK,G3445,G3441);
  and GNAME3447(G3447,G3445,G3448);
  nand GNAME3448(G3448,G80,G3450);
  buf GNAME3449(G3449,G3445);
  buf GNAME3450(G3450,G3432);
  or GNAME3462(G3462,G3464,G3463);
  and GNAME3463(G3463,G11542,G402);
  and GNAME3464(G3464,G3466,G3465);
  not GNAME3465(G3465,G402);
  dff DFF_3467(CK,G3466,G3462);
  and GNAME3468(G3468,G3466,G3469);
  nand GNAME3469(G3469,G80,G3471);
  buf GNAME3470(G3470,G3466);
  buf GNAME3471(G3471,G3453);
  or GNAME3483(G3483,G3485,G3484);
  and GNAME3484(G3484,G11541,G402);
  and GNAME3485(G3485,G3487,G3486);
  not GNAME3486(G3486,G402);
  dff DFF_3488(CK,G3487,G3483);
  and GNAME3489(G3489,G3487,G3490);
  nand GNAME3490(G3490,G80,G3492);
  buf GNAME3491(G3491,G3487);
  buf GNAME3492(G3492,G3474);
  or GNAME3504(G3504,G3506,G3505);
  and GNAME3505(G3505,G11540,G402);
  and GNAME3506(G3506,G3508,G3507);
  not GNAME3507(G3507,G402);
  dff DFF_3509(CK,G3508,G3504);
  and GNAME3510(G3510,G3508,G3511);
  nand GNAME3511(G3511,G80,G3513);
  buf GNAME3512(G3512,G3508);
  buf GNAME3513(G3513,G3495);
  or GNAME3525(G3525,G3527,G3526);
  and GNAME3526(G3526,G11539,G402);
  and GNAME3527(G3527,G3529,G3528);
  not GNAME3528(G3528,G402);
  dff DFF_3530(CK,G3529,G3525);
  and GNAME3531(G3531,G3529,G3532);
  nand GNAME3532(G3532,G80,G3534);
  buf GNAME3533(G3533,G3529);
  buf GNAME3534(G3534,G3516);
  or GNAME3546(G3546,G3548,G3547);
  and GNAME3547(G3547,G11522,G395);
  and GNAME3548(G3548,G3550,G3549);
  not GNAME3549(G3549,G395);
  dff DFF_3551(CK,G3550,G3546);
  and GNAME3552(G3552,G3550,G3553);
  nand GNAME3553(G3553,G80,G3555);
  buf GNAME3554(G3554,G3550);
  buf GNAME3555(G3555,G3537);
  or GNAME3607(G3607,G3609,G3608);
  and GNAME3608(G3608,G11546,G401);
  and GNAME3609(G3609,G3611,G3610);
  not GNAME3610(G3610,G401);
  dff DFF_3612(CK,G3611,G3607);
  and GNAME3613(G3613,G3611,G3614);
  nand GNAME3614(G3614,G80,G3616);
  buf GNAME3615(G3615,G3611);
  buf GNAME3616(G3616,G3598);
  or GNAME3628(G3628,G3630,G3629);
  and GNAME3629(G3629,G11545,G401);
  and GNAME3630(G3630,G3632,G3631);
  not GNAME3631(G3631,G401);
  dff DFF_3633(CK,G3632,G3628);
  and GNAME3634(G3634,G3632,G3635);
  nand GNAME3635(G3635,G80,G3637);
  buf GNAME3636(G3636,G3632);
  buf GNAME3637(G3637,G3619);
  or GNAME3649(G3649,G3651,G3650);
  and GNAME3650(G3650,G11544,G401);
  and GNAME3651(G3651,G3653,G3652);
  not GNAME3652(G3652,G401);
  dff DFF_3654(CK,G3653,G3649);
  and GNAME3655(G3655,G3653,G3656);
  nand GNAME3656(G3656,G80,G3658);
  buf GNAME3657(G3657,G3653);
  buf GNAME3658(G3658,G3640);
  or GNAME3670(G3670,G3672,G3671);
  and GNAME3671(G3671,G11543,G401);
  and GNAME3672(G3672,G3674,G3673);
  not GNAME3673(G3673,G401);
  dff DFF_3675(CK,G3674,G3670);
  and GNAME3676(G3676,G3674,G3677);
  nand GNAME3677(G3677,G80,G3679);
  buf GNAME3678(G3678,G3674);
  buf GNAME3679(G3679,G3661);
  or GNAME3691(G3691,G3693,G3692);
  and GNAME3692(G3692,G11542,G401);
  and GNAME3693(G3693,G3695,G3694);
  not GNAME3694(G3694,G401);
  dff DFF_3696(CK,G3695,G3691);
  and GNAME3697(G3697,G3695,G3698);
  nand GNAME3698(G3698,G80,G3700);
  buf GNAME3699(G3699,G3695);
  buf GNAME3700(G3700,G3682);
  or GNAME3712(G3712,G3714,G3713);
  and GNAME3713(G3713,G11541,G401);
  and GNAME3714(G3714,G3716,G3715);
  not GNAME3715(G3715,G401);
  dff DFF_3717(CK,G3716,G3712);
  and GNAME3718(G3718,G3716,G3719);
  nand GNAME3719(G3719,G80,G3721);
  buf GNAME3720(G3720,G3716);
  buf GNAME3721(G3721,G3703);
  or GNAME3733(G3733,G3735,G3734);
  and GNAME3734(G3734,G11540,G401);
  and GNAME3735(G3735,G3737,G3736);
  not GNAME3736(G3736,G401);
  dff DFF_3738(CK,G3737,G3733);
  and GNAME3739(G3739,G3737,G3740);
  nand GNAME3740(G3740,G80,G3742);
  buf GNAME3741(G3741,G3737);
  buf GNAME3742(G3742,G3724);
  or GNAME3754(G3754,G3756,G3755);
  and GNAME3755(G3755,G11539,G401);
  and GNAME3756(G3756,G3758,G3757);
  not GNAME3757(G3757,G401);
  dff DFF_3759(CK,G3758,G3754);
  and GNAME3760(G3760,G3758,G3761);
  nand GNAME3761(G3761,G80,G3763);
  buf GNAME3762(G3762,G3758);
  buf GNAME3763(G3763,G3745);
  or GNAME3815(G3815,G3817,G3816);
  and GNAME3816(G3816,G11546,G400);
  and GNAME3817(G3817,G3819,G3818);
  not GNAME3818(G3818,G400);
  dff DFF_3820(CK,G3819,G3815);
  and GNAME3821(G3821,G3819,G3822);
  nand GNAME3822(G3822,G80,G3824);
  buf GNAME3823(G3823,G3819);
  buf GNAME3824(G3824,G3806);
  or GNAME3836(G3836,G3838,G3837);
  and GNAME3837(G3837,G11545,G400);
  and GNAME3838(G3838,G3840,G3839);
  not GNAME3839(G3839,G400);
  dff DFF_3841(CK,G3840,G3836);
  and GNAME3842(G3842,G3840,G3843);
  nand GNAME3843(G3843,G80,G3845);
  buf GNAME3844(G3844,G3840);
  buf GNAME3845(G3845,G3827);
  or GNAME3857(G3857,G3859,G3858);
  and GNAME3858(G3858,G11544,G400);
  and GNAME3859(G3859,G3861,G3860);
  not GNAME3860(G3860,G400);
  dff DFF_3862(CK,G3861,G3857);
  and GNAME3863(G3863,G3861,G3864);
  nand GNAME3864(G3864,G80,G3866);
  buf GNAME3865(G3865,G3861);
  buf GNAME3866(G3866,G3848);
  or GNAME3878(G3878,G3880,G3879);
  and GNAME3879(G3879,G11543,G400);
  and GNAME3880(G3880,G3882,G3881);
  not GNAME3881(G3881,G400);
  dff DFF_3883(CK,G3882,G3878);
  and GNAME3884(G3884,G3882,G3885);
  nand GNAME3885(G3885,G80,G3887);
  buf GNAME3886(G3886,G3882);
  buf GNAME3887(G3887,G3869);
  or GNAME3899(G3899,G3901,G3900);
  and GNAME3900(G3900,G11542,G400);
  and GNAME3901(G3901,G3903,G3902);
  not GNAME3902(G3902,G400);
  dff DFF_3904(CK,G3903,G3899);
  and GNAME3905(G3905,G3903,G3906);
  nand GNAME3906(G3906,G80,G3908);
  buf GNAME3907(G3907,G3903);
  buf GNAME3908(G3908,G3890);
  or GNAME3920(G3920,G3922,G3921);
  and GNAME3921(G3921,G11541,G400);
  and GNAME3922(G3922,G3924,G3923);
  not GNAME3923(G3923,G400);
  dff DFF_3925(CK,G3924,G3920);
  and GNAME3926(G3926,G3924,G3927);
  nand GNAME3927(G3927,G80,G3929);
  buf GNAME3928(G3928,G3924);
  buf GNAME3929(G3929,G3911);
  or GNAME3941(G3941,G3943,G3942);
  and GNAME3942(G3942,G11540,G400);
  and GNAME3943(G3943,G3945,G3944);
  not GNAME3944(G3944,G400);
  dff DFF_3946(CK,G3945,G3941);
  and GNAME3947(G3947,G3945,G3948);
  nand GNAME3948(G3948,G80,G3950);
  buf GNAME3949(G3949,G3945);
  buf GNAME3950(G3950,G3932);
  or GNAME3962(G3962,G3964,G3963);
  and GNAME3963(G3963,G11539,G400);
  and GNAME3964(G3964,G3966,G3965);
  not GNAME3965(G3965,G400);
  dff DFF_3967(CK,G3966,G3962);
  and GNAME3968(G3968,G3966,G3969);
  nand GNAME3969(G3969,G80,G3971);
  buf GNAME3970(G3970,G3966);
  buf GNAME3971(G3971,G3953);
  or GNAME4023(G4023,G4025,G4024);
  and GNAME4024(G4024,G11538,G399);
  and GNAME4025(G4025,G4027,G4026);
  not GNAME4026(G4026,G399);
  dff DFF_4028(CK,G4027,G4023);
  and GNAME4029(G4029,G4027,G4030);
  nand GNAME4030(G4030,G80,G4032);
  buf GNAME4031(G4031,G4027);
  buf GNAME4032(G4032,G4014);
  or GNAME4044(G4044,G4046,G4045);
  and GNAME4045(G4045,G11545,G399);
  and GNAME4046(G4046,G4048,G4047);
  not GNAME4047(G4047,G399);
  dff DFF_4049(CK,G4048,G4044);
  and GNAME4050(G4050,G4048,G4051);
  nand GNAME4051(G4051,G80,G4053);
  buf GNAME4052(G4052,G4048);
  buf GNAME4053(G4053,G4035);
  or GNAME4065(G4065,G4067,G4066);
  and GNAME4066(G4066,G11544,G399);
  and GNAME4067(G4067,G4069,G4068);
  not GNAME4068(G4068,G399);
  dff DFF_4070(CK,G4069,G4065);
  and GNAME4071(G4071,G4069,G4072);
  nand GNAME4072(G4072,G80,G4074);
  buf GNAME4073(G4073,G4069);
  buf GNAME4074(G4074,G4056);
  or GNAME4086(G4086,G4088,G4087);
  and GNAME4087(G4087,G11543,G399);
  and GNAME4088(G4088,G4090,G4089);
  not GNAME4089(G4089,G399);
  dff DFF_4091(CK,G4090,G4086);
  and GNAME4092(G4092,G4090,G4093);
  nand GNAME4093(G4093,G80,G4095);
  buf GNAME4094(G4094,G4090);
  buf GNAME4095(G4095,G4077);
  or GNAME4107(G4107,G4109,G4108);
  and GNAME4108(G4108,G11542,G399);
  and GNAME4109(G4109,G4111,G4110);
  not GNAME4110(G4110,G399);
  dff DFF_4112(CK,G4111,G4107);
  and GNAME4113(G4113,G4111,G4114);
  nand GNAME4114(G4114,G80,G4116);
  buf GNAME4115(G4115,G4111);
  buf GNAME4116(G4116,G4098);
  or GNAME4128(G4128,G4130,G4129);
  and GNAME4129(G4129,G11541,G399);
  and GNAME4130(G4130,G4132,G4131);
  not GNAME4131(G4131,G399);
  dff DFF_4133(CK,G4132,G4128);
  and GNAME4134(G4134,G4132,G4135);
  nand GNAME4135(G4135,G80,G4137);
  buf GNAME4136(G4136,G4132);
  buf GNAME4137(G4137,G4119);
  or GNAME4149(G4149,G4151,G4150);
  and GNAME4150(G4150,G11540,G399);
  and GNAME4151(G4151,G4153,G4152);
  not GNAME4152(G4152,G399);
  dff DFF_4154(CK,G4153,G4149);
  and GNAME4155(G4155,G4153,G4156);
  nand GNAME4156(G4156,G80,G4158);
  buf GNAME4157(G4157,G4153);
  buf GNAME4158(G4158,G4140);
  or GNAME4170(G4170,G4172,G4171);
  and GNAME4171(G4171,G11539,G399);
  and GNAME4172(G4172,G4174,G4173);
  not GNAME4173(G4173,G399);
  dff DFF_4175(CK,G4174,G4170);
  and GNAME4176(G4176,G4174,G4177);
  nand GNAME4177(G4177,G80,G4179);
  buf GNAME4178(G4178,G4174);
  buf GNAME4179(G4179,G4161);
  or GNAME4231(G4231,G4233,G4232);
  and GNAME4232(G4232,G11538,G398);
  and GNAME4233(G4233,G4235,G4234);
  not GNAME4234(G4234,G398);
  dff DFF_4236(CK,G4235,G4231);
  and GNAME4237(G4237,G4235,G4238);
  nand GNAME4238(G4238,G80,G4240);
  buf GNAME4239(G4239,G4235);
  buf GNAME4240(G4240,G4222);
  or GNAME4252(G4252,G4254,G4253);
  and GNAME4253(G4253,G11537,G398);
  and GNAME4254(G4254,G4256,G4255);
  not GNAME4255(G4255,G398);
  dff DFF_4257(CK,G4256,G4252);
  and GNAME4258(G4258,G4256,G4259);
  nand GNAME4259(G4259,G80,G4261);
  buf GNAME4260(G4260,G4256);
  buf GNAME4261(G4261,G4243);
  or GNAME4273(G4273,G4275,G4274);
  and GNAME4274(G4274,G11536,G398);
  and GNAME4275(G4275,G4277,G4276);
  not GNAME4276(G4276,G398);
  dff DFF_4278(CK,G4277,G4273);
  and GNAME4279(G4279,G4277,G4280);
  nand GNAME4280(G4280,G80,G4282);
  buf GNAME4281(G4281,G4277);
  buf GNAME4282(G4282,G4264);
  or GNAME4294(G4294,G4296,G4295);
  and GNAME4295(G4295,G11535,G398);
  and GNAME4296(G4296,G4298,G4297);
  not GNAME4297(G4297,G398);
  dff DFF_4299(CK,G4298,G4294);
  and GNAME4300(G4300,G4298,G4301);
  nand GNAME4301(G4301,G80,G4303);
  buf GNAME4302(G4302,G4298);
  buf GNAME4303(G4303,G4285);
  or GNAME4315(G4315,G4317,G4316);
  and GNAME4316(G4316,G11534,G398);
  and GNAME4317(G4317,G4319,G4318);
  not GNAME4318(G4318,G398);
  dff DFF_4320(CK,G4319,G4315);
  and GNAME4321(G4321,G4319,G4322);
  nand GNAME4322(G4322,G80,G4324);
  buf GNAME4323(G4323,G4319);
  buf GNAME4324(G4324,G4306);
  or GNAME4336(G4336,G4338,G4337);
  and GNAME4337(G4337,G11533,G398);
  and GNAME4338(G4338,G4340,G4339);
  not GNAME4339(G4339,G398);
  dff DFF_4341(CK,G4340,G4336);
  and GNAME4342(G4342,G4340,G4343);
  nand GNAME4343(G4343,G80,G4345);
  buf GNAME4344(G4344,G4340);
  buf GNAME4345(G4345,G4327);
  or GNAME4357(G4357,G4359,G4358);
  and GNAME4358(G4358,G11532,G398);
  and GNAME4359(G4359,G4361,G4360);
  not GNAME4360(G4360,G398);
  dff DFF_4362(CK,G4361,G4357);
  and GNAME4363(G4363,G4361,G4364);
  nand GNAME4364(G4364,G80,G4366);
  buf GNAME4365(G4365,G4361);
  buf GNAME4366(G4366,G4348);
  or GNAME4378(G4378,G4380,G4379);
  and GNAME4379(G4379,G11531,G398);
  and GNAME4380(G4380,G4382,G4381);
  not GNAME4381(G4381,G398);
  dff DFF_4383(CK,G4382,G4378);
  and GNAME4384(G4384,G4382,G4385);
  nand GNAME4385(G4385,G80,G4387);
  buf GNAME4386(G4386,G4382);
  buf GNAME4387(G4387,G4369);
  or GNAME4399(G4399,G4401,G4400);
  and GNAME4400(G4400,G11522,G396);
  and GNAME4401(G4401,G4403,G4402);
  not GNAME4402(G4402,G396);
  dff DFF_4404(CK,G4403,G4399);
  and GNAME4405(G4405,G4403,G4406);
  nand GNAME4406(G4406,G80,G4408);
  buf GNAME4407(G4407,G4403);
  buf GNAME4408(G4408,G4390);
  or GNAME4460(G4460,G4462,G4461);
  and GNAME4461(G4461,G11538,G434);
  and GNAME4462(G4462,G4464,G4463);
  not GNAME4463(G4463,G434);
  dff DFF_4465(CK,G4464,G4460);
  and GNAME4466(G4466,G4464,G4467);
  nand GNAME4467(G4467,G80,G4469);
  buf GNAME4468(G4468,G4464);
  buf GNAME4469(G4469,G4451);
  or GNAME4481(G4481,G4483,G4482);
  and GNAME4482(G4482,G11537,G434);
  and GNAME4483(G4483,G4485,G4484);
  not GNAME4484(G4484,G434);
  dff DFF_4486(CK,G4485,G4481);
  and GNAME4487(G4487,G4485,G4488);
  nand GNAME4488(G4488,G80,G4490);
  buf GNAME4489(G4489,G4485);
  buf GNAME4490(G4490,G4472);
  or GNAME4502(G4502,G4504,G4503);
  and GNAME4503(G4503,G11536,G434);
  and GNAME4504(G4504,G4506,G4505);
  not GNAME4505(G4505,G434);
  dff DFF_4507(CK,G4506,G4502);
  and GNAME4508(G4508,G4506,G4509);
  nand GNAME4509(G4509,G80,G4511);
  buf GNAME4510(G4510,G4506);
  buf GNAME4511(G4511,G4493);
  or GNAME4523(G4523,G4525,G4524);
  and GNAME4524(G4524,G11535,G434);
  and GNAME4525(G4525,G4527,G4526);
  not GNAME4526(G4526,G434);
  dff DFF_4528(CK,G4527,G4523);
  and GNAME4529(G4529,G4527,G4530);
  nand GNAME4530(G4530,G80,G4532);
  buf GNAME4531(G4531,G4527);
  buf GNAME4532(G4532,G4514);
  or GNAME4544(G4544,G4546,G4545);
  and GNAME4545(G4545,G11534,G434);
  and GNAME4546(G4546,G4548,G4547);
  not GNAME4547(G4547,G434);
  dff DFF_4549(CK,G4548,G4544);
  and GNAME4550(G4550,G4548,G4551);
  nand GNAME4551(G4551,G80,G4553);
  buf GNAME4552(G4552,G4548);
  buf GNAME4553(G4553,G4535);
  or GNAME4565(G4565,G4567,G4566);
  and GNAME4566(G4566,G11533,G434);
  and GNAME4567(G4567,G4569,G4568);
  not GNAME4568(G4568,G434);
  dff DFF_4570(CK,G4569,G4565);
  and GNAME4571(G4571,G4569,G4572);
  nand GNAME4572(G4572,G80,G4574);
  buf GNAME4573(G4573,G4569);
  buf GNAME4574(G4574,G4556);
  or GNAME4586(G4586,G4588,G4587);
  and GNAME4587(G4587,G11532,G434);
  and GNAME4588(G4588,G4590,G4589);
  not GNAME4589(G4589,G434);
  dff DFF_4591(CK,G4590,G4586);
  and GNAME4592(G4592,G4590,G4593);
  nand GNAME4593(G4593,G80,G4595);
  buf GNAME4594(G4594,G4590);
  buf GNAME4595(G4595,G4577);
  or GNAME4607(G4607,G4609,G4608);
  and GNAME4608(G4608,G11531,G434);
  and GNAME4609(G4609,G4611,G4610);
  not GNAME4610(G4610,G434);
  dff DFF_4612(CK,G4611,G4607);
  and GNAME4613(G4613,G4611,G4614);
  nand GNAME4614(G4614,G80,G4616);
  buf GNAME4615(G4615,G4611);
  buf GNAME4616(G4616,G4598);
  or GNAME4668(G4668,G4670,G4669);
  and GNAME4669(G4669,G11538,G433);
  and GNAME4670(G4670,G4672,G4671);
  not GNAME4671(G4671,G433);
  dff DFF_4673(CK,G4672,G4668);
  and GNAME4674(G4674,G4672,G4675);
  nand GNAME4675(G4675,G80,G4677);
  buf GNAME4676(G4676,G4672);
  buf GNAME4677(G4677,G4659);
  or GNAME4689(G4689,G4691,G4690);
  and GNAME4690(G4690,G11537,G433);
  and GNAME4691(G4691,G4693,G4692);
  not GNAME4692(G4692,G433);
  dff DFF_4694(CK,G4693,G4689);
  and GNAME4695(G4695,G4693,G4696);
  nand GNAME4696(G4696,G80,G4698);
  buf GNAME4697(G4697,G4693);
  buf GNAME4698(G4698,G4680);
  or GNAME4710(G4710,G4712,G4711);
  and GNAME4711(G4711,G11536,G433);
  and GNAME4712(G4712,G4714,G4713);
  not GNAME4713(G4713,G433);
  dff DFF_4715(CK,G4714,G4710);
  and GNAME4716(G4716,G4714,G4717);
  nand GNAME4717(G4717,G80,G4719);
  buf GNAME4718(G4718,G4714);
  buf GNAME4719(G4719,G4701);
  or GNAME4731(G4731,G4733,G4732);
  and GNAME4732(G4732,G11535,G433);
  and GNAME4733(G4733,G4735,G4734);
  not GNAME4734(G4734,G433);
  dff DFF_4736(CK,G4735,G4731);
  and GNAME4737(G4737,G4735,G4738);
  nand GNAME4738(G4738,G80,G4740);
  buf GNAME4739(G4739,G4735);
  buf GNAME4740(G4740,G4722);
  or GNAME4752(G4752,G4754,G4753);
  and GNAME4753(G4753,G11534,G433);
  and GNAME4754(G4754,G4756,G4755);
  not GNAME4755(G4755,G433);
  dff DFF_4757(CK,G4756,G4752);
  and GNAME4758(G4758,G4756,G4759);
  nand GNAME4759(G4759,G80,G4761);
  buf GNAME4760(G4760,G4756);
  buf GNAME4761(G4761,G4743);
  or GNAME4773(G4773,G4775,G4774);
  and GNAME4774(G4774,G11533,G433);
  and GNAME4775(G4775,G4777,G4776);
  not GNAME4776(G4776,G433);
  dff DFF_4778(CK,G4777,G4773);
  and GNAME4779(G4779,G4777,G4780);
  nand GNAME4780(G4780,G80,G4782);
  buf GNAME4781(G4781,G4777);
  buf GNAME4782(G4782,G4764);
  or GNAME4794(G4794,G4796,G4795);
  and GNAME4795(G4795,G11532,G433);
  and GNAME4796(G4796,G4798,G4797);
  not GNAME4797(G4797,G433);
  dff DFF_4799(CK,G4798,G4794);
  and GNAME4800(G4800,G4798,G4801);
  nand GNAME4801(G4801,G80,G4803);
  buf GNAME4802(G4802,G4798);
  buf GNAME4803(G4803,G4785);
  or GNAME4815(G4815,G4817,G4816);
  and GNAME4816(G4816,G11531,G433);
  and GNAME4817(G4817,G4819,G4818);
  not GNAME4818(G4818,G433);
  dff DFF_4820(CK,G4819,G4815);
  and GNAME4821(G4821,G4819,G4822);
  nand GNAME4822(G4822,G80,G4824);
  buf GNAME4823(G4823,G4819);
  buf GNAME4824(G4824,G4806);
  or GNAME4876(G4876,G4878,G4877);
  and GNAME4877(G4877,G11538,G432);
  and GNAME4878(G4878,G4880,G4879);
  not GNAME4879(G4879,G432);
  dff DFF_4881(CK,G4880,G4876);
  and GNAME4882(G4882,G4880,G4883);
  nand GNAME4883(G4883,G80,G4885);
  buf GNAME4884(G4884,G4880);
  buf GNAME4885(G4885,G4867);
  or GNAME4897(G4897,G4899,G4898);
  and GNAME4898(G4898,G11537,G432);
  and GNAME4899(G4899,G4901,G4900);
  not GNAME4900(G4900,G432);
  dff DFF_4902(CK,G4901,G4897);
  and GNAME4903(G4903,G4901,G4904);
  nand GNAME4904(G4904,G80,G4906);
  buf GNAME4905(G4905,G4901);
  buf GNAME4906(G4906,G4888);
  or GNAME4918(G4918,G4920,G4919);
  and GNAME4919(G4919,G11536,G432);
  and GNAME4920(G4920,G4922,G4921);
  not GNAME4921(G4921,G432);
  dff DFF_4923(CK,G4922,G4918);
  and GNAME4924(G4924,G4922,G4925);
  nand GNAME4925(G4925,G80,G4927);
  buf GNAME4926(G4926,G4922);
  buf GNAME4927(G4927,G4909);
  or GNAME4939(G4939,G4941,G4940);
  and GNAME4940(G4940,G11535,G432);
  and GNAME4941(G4941,G4943,G4942);
  not GNAME4942(G4942,G432);
  dff DFF_4944(CK,G4943,G4939);
  and GNAME4945(G4945,G4943,G4946);
  nand GNAME4946(G4946,G80,G4948);
  buf GNAME4947(G4947,G4943);
  buf GNAME4948(G4948,G4930);
  or GNAME4960(G4960,G4962,G4961);
  and GNAME4961(G4961,G11534,G432);
  and GNAME4962(G4962,G4964,G4963);
  not GNAME4963(G4963,G432);
  dff DFF_4965(CK,G4964,G4960);
  and GNAME4966(G4966,G4964,G4967);
  nand GNAME4967(G4967,G80,G4969);
  buf GNAME4968(G4968,G4964);
  buf GNAME4969(G4969,G4951);
  or GNAME4981(G4981,G4983,G4982);
  and GNAME4982(G4982,G11533,G432);
  and GNAME4983(G4983,G4985,G4984);
  not GNAME4984(G4984,G432);
  dff DFF_4986(CK,G4985,G4981);
  and GNAME4987(G4987,G4985,G4988);
  nand GNAME4988(G4988,G80,G4990);
  buf GNAME4989(G4989,G4985);
  buf GNAME4990(G4990,G4972);
  or GNAME5002(G5002,G5004,G5003);
  and GNAME5003(G5003,G11532,G432);
  and GNAME5004(G5004,G5006,G5005);
  not GNAME5005(G5005,G432);
  dff DFF_5007(CK,G5006,G5002);
  and GNAME5008(G5008,G5006,G5009);
  nand GNAME5009(G5009,G80,G5011);
  buf GNAME5010(G5010,G5006);
  buf GNAME5011(G5011,G4993);
  or GNAME5023(G5023,G5025,G5024);
  and GNAME5024(G5024,G11531,G432);
  and GNAME5025(G5025,G5027,G5026);
  not GNAME5026(G5026,G432);
  dff DFF_5028(CK,G5027,G5023);
  and GNAME5029(G5029,G5027,G5030);
  nand GNAME5030(G5030,G80,G5032);
  buf GNAME5031(G5031,G5027);
  buf GNAME5032(G5032,G5014);
  or GNAME5084(G5084,G5086,G5085);
  and GNAME5085(G5085,G11538,G431);
  and GNAME5086(G5086,G5088,G5087);
  not GNAME5087(G5087,G431);
  dff DFF_5089(CK,G5088,G5084);
  and GNAME5090(G5090,G5088,G5091);
  nand GNAME5091(G5091,G80,G5093);
  buf GNAME5092(G5092,G5088);
  buf GNAME5093(G5093,G5075);
  or GNAME5105(G5105,G5107,G5106);
  and GNAME5106(G5106,G11537,G431);
  and GNAME5107(G5107,G5109,G5108);
  not GNAME5108(G5108,G431);
  dff DFF_5110(CK,G5109,G5105);
  and GNAME5111(G5111,G5109,G5112);
  nand GNAME5112(G5112,G80,G5114);
  buf GNAME5113(G5113,G5109);
  buf GNAME5114(G5114,G5096);
  or GNAME5126(G5126,G5128,G5127);
  and GNAME5127(G5127,G11536,G431);
  and GNAME5128(G5128,G5130,G5129);
  not GNAME5129(G5129,G431);
  dff DFF_5131(CK,G5130,G5126);
  and GNAME5132(G5132,G5130,G5133);
  nand GNAME5133(G5133,G80,G5135);
  buf GNAME5134(G5134,G5130);
  buf GNAME5135(G5135,G5117);
  or GNAME5147(G5147,G5149,G5148);
  and GNAME5148(G5148,G11535,G431);
  and GNAME5149(G5149,G5151,G5150);
  not GNAME5150(G5150,G431);
  dff DFF_5152(CK,G5151,G5147);
  and GNAME5153(G5153,G5151,G5154);
  nand GNAME5154(G5154,G80,G5156);
  buf GNAME5155(G5155,G5151);
  buf GNAME5156(G5156,G5138);
  or GNAME5168(G5168,G5170,G5169);
  and GNAME5169(G5169,G11534,G431);
  and GNAME5170(G5170,G5172,G5171);
  not GNAME5171(G5171,G431);
  dff DFF_5173(CK,G5172,G5168);
  and GNAME5174(G5174,G5172,G5175);
  nand GNAME5175(G5175,G80,G5177);
  buf GNAME5176(G5176,G5172);
  buf GNAME5177(G5177,G5159);
  or GNAME5189(G5189,G5191,G5190);
  and GNAME5190(G5190,G11533,G431);
  and GNAME5191(G5191,G5193,G5192);
  not GNAME5192(G5192,G431);
  dff DFF_5194(CK,G5193,G5189);
  and GNAME5195(G5195,G5193,G5196);
  nand GNAME5196(G5196,G80,G5198);
  buf GNAME5197(G5197,G5193);
  buf GNAME5198(G5198,G5180);
  or GNAME5210(G5210,G5212,G5211);
  and GNAME5211(G5211,G11532,G431);
  and GNAME5212(G5212,G5214,G5213);
  not GNAME5213(G5213,G431);
  dff DFF_5215(CK,G5214,G5210);
  and GNAME5216(G5216,G5214,G5217);
  nand GNAME5217(G5217,G80,G5219);
  buf GNAME5218(G5218,G5214);
  buf GNAME5219(G5219,G5201);
  or GNAME5231(G5231,G5233,G5232);
  and GNAME5232(G5232,G11531,G431);
  and GNAME5233(G5233,G5235,G5234);
  not GNAME5234(G5234,G431);
  dff DFF_5236(CK,G5235,G5231);
  and GNAME5237(G5237,G5235,G5238);
  nand GNAME5238(G5238,G80,G5240);
  buf GNAME5239(G5239,G5235);
  buf GNAME5240(G5240,G5222);
  or GNAME5252(G5252,G5254,G5253);
  and GNAME5253(G5253,G11546,G397);
  and GNAME5254(G5254,G5256,G5255);
  not GNAME5255(G5255,G397);
  dff DFF_5257(CK,G5256,G5252);
  and GNAME5258(G5258,G5256,G5259);
  nand GNAME5259(G5259,G80,G5261);
  buf GNAME5260(G5260,G5256);
  buf GNAME5261(G5261,G5243);
  or GNAME5313(G5313,G5315,G5314);
  and GNAME5314(G5314,G11538,G430);
  and GNAME5315(G5315,G5317,G5316);
  not GNAME5316(G5316,G430);
  dff DFF_5318(CK,G5317,G5313);
  and GNAME5319(G5319,G5317,G5320);
  nand GNAME5320(G5320,G80,G5322);
  buf GNAME5321(G5321,G5317);
  buf GNAME5322(G5322,G5304);
  or GNAME5334(G5334,G5336,G5335);
  and GNAME5335(G5335,G11537,G430);
  and GNAME5336(G5336,G5338,G5337);
  not GNAME5337(G5337,G430);
  dff DFF_5339(CK,G5338,G5334);
  and GNAME5340(G5340,G5338,G5341);
  nand GNAME5341(G5341,G80,G5343);
  buf GNAME5342(G5342,G5338);
  buf GNAME5343(G5343,G5325);
  or GNAME5355(G5355,G5357,G5356);
  and GNAME5356(G5356,G11536,G430);
  and GNAME5357(G5357,G5359,G5358);
  not GNAME5358(G5358,G430);
  dff DFF_5360(CK,G5359,G5355);
  and GNAME5361(G5361,G5359,G5362);
  nand GNAME5362(G5362,G80,G5364);
  buf GNAME5363(G5363,G5359);
  buf GNAME5364(G5364,G5346);
  or GNAME5376(G5376,G5378,G5377);
  and GNAME5377(G5377,G11535,G430);
  and GNAME5378(G5378,G5380,G5379);
  not GNAME5379(G5379,G430);
  dff DFF_5381(CK,G5380,G5376);
  and GNAME5382(G5382,G5380,G5383);
  nand GNAME5383(G5383,G80,G5385);
  buf GNAME5384(G5384,G5380);
  buf GNAME5385(G5385,G5367);
  or GNAME5397(G5397,G5399,G5398);
  and GNAME5398(G5398,G11534,G430);
  and GNAME5399(G5399,G5401,G5400);
  not GNAME5400(G5400,G430);
  dff DFF_5402(CK,G5401,G5397);
  and GNAME5403(G5403,G5401,G5404);
  nand GNAME5404(G5404,G80,G5406);
  buf GNAME5405(G5405,G5401);
  buf GNAME5406(G5406,G5388);
  or GNAME5418(G5418,G5420,G5419);
  and GNAME5419(G5419,G11533,G430);
  and GNAME5420(G5420,G5422,G5421);
  not GNAME5421(G5421,G430);
  dff DFF_5423(CK,G5422,G5418);
  and GNAME5424(G5424,G5422,G5425);
  nand GNAME5425(G5425,G80,G5427);
  buf GNAME5426(G5426,G5422);
  buf GNAME5427(G5427,G5409);
  or GNAME5439(G5439,G5441,G5440);
  and GNAME5440(G5440,G11532,G430);
  and GNAME5441(G5441,G5443,G5442);
  not GNAME5442(G5442,G430);
  dff DFF_5444(CK,G5443,G5439);
  and GNAME5445(G5445,G5443,G5446);
  nand GNAME5446(G5446,G80,G5448);
  buf GNAME5447(G5447,G5443);
  buf GNAME5448(G5448,G5430);
  or GNAME5460(G5460,G5462,G5461);
  and GNAME5461(G5461,G11531,G430);
  and GNAME5462(G5462,G5464,G5463);
  not GNAME5463(G5463,G430);
  dff DFF_5465(CK,G5464,G5460);
  and GNAME5466(G5466,G5464,G5467);
  nand GNAME5467(G5467,G80,G5469);
  buf GNAME5468(G5468,G5464);
  buf GNAME5469(G5469,G5451);
  or GNAME5521(G5521,G5523,G5522);
  and GNAME5522(G5522,G11538,G429);
  and GNAME5523(G5523,G5525,G5524);
  not GNAME5524(G5524,G429);
  dff DFF_5526(CK,G5525,G5521);
  and GNAME5527(G5527,G5525,G5528);
  nand GNAME5528(G5528,G80,G5530);
  buf GNAME5529(G5529,G5525);
  buf GNAME5530(G5530,G5512);
  or GNAME5542(G5542,G5544,G5543);
  and GNAME5543(G5543,G11537,G429);
  and GNAME5544(G5544,G5546,G5545);
  not GNAME5545(G5545,G429);
  dff DFF_5547(CK,G5546,G5542);
  and GNAME5548(G5548,G5546,G5549);
  nand GNAME5549(G5549,G80,G5551);
  buf GNAME5550(G5550,G5546);
  buf GNAME5551(G5551,G5533);
  or GNAME5563(G5563,G5565,G5564);
  and GNAME5564(G5564,G11536,G429);
  and GNAME5565(G5565,G5567,G5566);
  not GNAME5566(G5566,G429);
  dff DFF_5568(CK,G5567,G5563);
  and GNAME5569(G5569,G5567,G5570);
  nand GNAME5570(G5570,G80,G5572);
  buf GNAME5571(G5571,G5567);
  buf GNAME5572(G5572,G5554);
  or GNAME5584(G5584,G5586,G5585);
  and GNAME5585(G5585,G11535,G429);
  and GNAME5586(G5586,G5588,G5587);
  not GNAME5587(G5587,G429);
  dff DFF_5589(CK,G5588,G5584);
  and GNAME5590(G5590,G5588,G5591);
  nand GNAME5591(G5591,G80,G5593);
  buf GNAME5592(G5592,G5588);
  buf GNAME5593(G5593,G5575);
  or GNAME5605(G5605,G5607,G5606);
  and GNAME5606(G5606,G11534,G429);
  and GNAME5607(G5607,G5609,G5608);
  not GNAME5608(G5608,G429);
  dff DFF_5610(CK,G5609,G5605);
  and GNAME5611(G5611,G5609,G5612);
  nand GNAME5612(G5612,G80,G5614);
  buf GNAME5613(G5613,G5609);
  buf GNAME5614(G5614,G5596);
  or GNAME5626(G5626,G5628,G5627);
  and GNAME5627(G5627,G11533,G429);
  and GNAME5628(G5628,G5630,G5629);
  not GNAME5629(G5629,G429);
  dff DFF_5631(CK,G5630,G5626);
  and GNAME5632(G5632,G5630,G5633);
  nand GNAME5633(G5633,G80,G5635);
  buf GNAME5634(G5634,G5630);
  buf GNAME5635(G5635,G5617);
  or GNAME5647(G5647,G5649,G5648);
  and GNAME5648(G5648,G11532,G429);
  and GNAME5649(G5649,G5651,G5650);
  not GNAME5650(G5650,G429);
  dff DFF_5652(CK,G5651,G5647);
  and GNAME5653(G5653,G5651,G5654);
  nand GNAME5654(G5654,G80,G5656);
  buf GNAME5655(G5655,G5651);
  buf GNAME5656(G5656,G5638);
  or GNAME5668(G5668,G5670,G5669);
  and GNAME5669(G5669,G11531,G429);
  and GNAME5670(G5670,G5672,G5671);
  not GNAME5671(G5671,G429);
  dff DFF_5673(CK,G5672,G5668);
  and GNAME5674(G5674,G5672,G5675);
  nand GNAME5675(G5675,G80,G5677);
  buf GNAME5676(G5676,G5672);
  buf GNAME5677(G5677,G5659);
  or GNAME5729(G5729,G5731,G5730);
  and GNAME5730(G5730,G11538,G428);
  and GNAME5731(G5731,G5733,G5732);
  not GNAME5732(G5732,G428);
  dff DFF_5734(CK,G5733,G5729);
  and GNAME5735(G5735,G5733,G5736);
  nand GNAME5736(G5736,G80,G5738);
  buf GNAME5737(G5737,G5733);
  buf GNAME5738(G5738,G5720);
  or GNAME5750(G5750,G5752,G5751);
  and GNAME5751(G5751,G11537,G428);
  and GNAME5752(G5752,G5754,G5753);
  not GNAME5753(G5753,G428);
  dff DFF_5755(CK,G5754,G5750);
  and GNAME5756(G5756,G5754,G5757);
  nand GNAME5757(G5757,G80,G5759);
  buf GNAME5758(G5758,G5754);
  buf GNAME5759(G5759,G5741);
  or GNAME5771(G5771,G5773,G5772);
  and GNAME5772(G5772,G11536,G428);
  and GNAME5773(G5773,G5775,G5774);
  not GNAME5774(G5774,G428);
  dff DFF_5776(CK,G5775,G5771);
  and GNAME5777(G5777,G5775,G5778);
  nand GNAME5778(G5778,G80,G5780);
  buf GNAME5779(G5779,G5775);
  buf GNAME5780(G5780,G5762);
  or GNAME5792(G5792,G5794,G5793);
  and GNAME5793(G5793,G11535,G428);
  and GNAME5794(G5794,G5796,G5795);
  not GNAME5795(G5795,G428);
  dff DFF_5797(CK,G5796,G5792);
  and GNAME5798(G5798,G5796,G5799);
  nand GNAME5799(G5799,G80,G5801);
  buf GNAME5800(G5800,G5796);
  buf GNAME5801(G5801,G5783);
  or GNAME5813(G5813,G5815,G5814);
  and GNAME5814(G5814,G11534,G428);
  and GNAME5815(G5815,G5817,G5816);
  not GNAME5816(G5816,G428);
  dff DFF_5818(CK,G5817,G5813);
  and GNAME5819(G5819,G5817,G5820);
  nand GNAME5820(G5820,G80,G5822);
  buf GNAME5821(G5821,G5817);
  buf GNAME5822(G5822,G5804);
  or GNAME5834(G5834,G5836,G5835);
  and GNAME5835(G5835,G11533,G428);
  and GNAME5836(G5836,G5838,G5837);
  not GNAME5837(G5837,G428);
  dff DFF_5839(CK,G5838,G5834);
  and GNAME5840(G5840,G5838,G5841);
  nand GNAME5841(G5841,G80,G5843);
  buf GNAME5842(G5842,G5838);
  buf GNAME5843(G5843,G5825);
  or GNAME5855(G5855,G5857,G5856);
  and GNAME5856(G5856,G11532,G428);
  and GNAME5857(G5857,G5859,G5858);
  not GNAME5858(G5858,G428);
  dff DFF_5860(CK,G5859,G5855);
  and GNAME5861(G5861,G5859,G5862);
  nand GNAME5862(G5862,G80,G5864);
  buf GNAME5863(G5863,G5859);
  buf GNAME5864(G5864,G5846);
  or GNAME5876(G5876,G5878,G5877);
  and GNAME5877(G5877,G11531,G428);
  and GNAME5878(G5878,G5880,G5879);
  not GNAME5879(G5879,G428);
  dff DFF_5881(CK,G5880,G5876);
  and GNAME5882(G5882,G5880,G5883);
  nand GNAME5883(G5883,G80,G5885);
  buf GNAME5884(G5884,G5880);
  buf GNAME5885(G5885,G5867);
  or GNAME5937(G5937,G5939,G5938);
  and GNAME5938(G5938,G11538,G411);
  and GNAME5939(G5939,G5941,G5940);
  not GNAME5940(G5940,G411);
  dff DFF_5942(CK,G5941,G5937);
  and GNAME5943(G5943,G5941,G5944);
  nand GNAME5944(G5944,G80,G5946);
  buf GNAME5945(G5945,G5941);
  buf GNAME5946(G5946,G5928);
  or GNAME5958(G5958,G5960,G5959);
  and GNAME5959(G5959,G11537,G411);
  and GNAME5960(G5960,G5962,G5961);
  not GNAME5961(G5961,G411);
  dff DFF_5963(CK,G5962,G5958);
  and GNAME5964(G5964,G5962,G5965);
  nand GNAME5965(G5965,G80,G5967);
  buf GNAME5966(G5966,G5962);
  buf GNAME5967(G5967,G5949);
  or GNAME5979(G5979,G5981,G5980);
  and GNAME5980(G5980,G11536,G411);
  and GNAME5981(G5981,G5983,G5982);
  not GNAME5982(G5982,G411);
  dff DFF_5984(CK,G5983,G5979);
  and GNAME5985(G5985,G5983,G5986);
  nand GNAME5986(G5986,G80,G5988);
  buf GNAME5987(G5987,G5983);
  buf GNAME5988(G5988,G5970);
  or GNAME6000(G6000,G6002,G6001);
  and GNAME6001(G6001,G11535,G411);
  and GNAME6002(G6002,G6004,G6003);
  not GNAME6003(G6003,G411);
  dff DFF_6005(CK,G6004,G6000);
  and GNAME6006(G6006,G6004,G6007);
  nand GNAME6007(G6007,G80,G6009);
  buf GNAME6008(G6008,G6004);
  buf GNAME6009(G6009,G5991);
  or GNAME6021(G6021,G6023,G6022);
  and GNAME6022(G6022,G11534,G411);
  and GNAME6023(G6023,G6025,G6024);
  not GNAME6024(G6024,G411);
  dff DFF_6026(CK,G6025,G6021);
  and GNAME6027(G6027,G6025,G6028);
  nand GNAME6028(G6028,G80,G6030);
  buf GNAME6029(G6029,G6025);
  buf GNAME6030(G6030,G6012);
  or GNAME6042(G6042,G6044,G6043);
  and GNAME6043(G6043,G11533,G411);
  and GNAME6044(G6044,G6046,G6045);
  not GNAME6045(G6045,G411);
  dff DFF_6047(CK,G6046,G6042);
  and GNAME6048(G6048,G6046,G6049);
  nand GNAME6049(G6049,G80,G6051);
  buf GNAME6050(G6050,G6046);
  buf GNAME6051(G6051,G6033);
  or GNAME6063(G6063,G6065,G6064);
  and GNAME6064(G6064,G11532,G411);
  and GNAME6065(G6065,G6067,G6066);
  not GNAME6066(G6066,G411);
  dff DFF_6068(CK,G6067,G6063);
  and GNAME6069(G6069,G6067,G6070);
  nand GNAME6070(G6070,G80,G6072);
  buf GNAME6071(G6071,G6067);
  buf GNAME6072(G6072,G6054);
  or GNAME6084(G6084,G6086,G6085);
  and GNAME6085(G6085,G11531,G411);
  and GNAME6086(G6086,G6088,G6087);
  not GNAME6087(G6087,G411);
  dff DFF_6089(CK,G6088,G6084);
  and GNAME6090(G6090,G6088,G6091);
  nand GNAME6091(G6091,G80,G6093);
  buf GNAME6092(G6092,G6088);
  buf GNAME6093(G6093,G6075);
  or GNAME6145(G6145,G6147,G6146);
  and GNAME6146(G6146,G11538,G410);
  and GNAME6147(G6147,G6149,G6148);
  not GNAME6148(G6148,G410);
  dff DFF_6150(CK,G6149,G6145);
  and GNAME6151(G6151,G6149,G6152);
  nand GNAME6152(G6152,G80,G6154);
  buf GNAME6153(G6153,G6149);
  buf GNAME6154(G6154,G6136);
  or GNAME6166(G6166,G6168,G6167);
  and GNAME6167(G6167,G11537,G410);
  and GNAME6168(G6168,G6170,G6169);
  not GNAME6169(G6169,G410);
  dff DFF_6171(CK,G6170,G6166);
  and GNAME6172(G6172,G6170,G6173);
  nand GNAME6173(G6173,G80,G6175);
  buf GNAME6174(G6174,G6170);
  buf GNAME6175(G6175,G6157);
  or GNAME6187(G6187,G6189,G6188);
  and GNAME6188(G6188,G11536,G410);
  and GNAME6189(G6189,G6191,G6190);
  not GNAME6190(G6190,G410);
  dff DFF_6192(CK,G6191,G6187);
  and GNAME6193(G6193,G6191,G6194);
  nand GNAME6194(G6194,G80,G6196);
  buf GNAME6195(G6195,G6191);
  buf GNAME6196(G6196,G6178);
  or GNAME6208(G6208,G6210,G6209);
  and GNAME6209(G6209,G11535,G410);
  and GNAME6210(G6210,G6212,G6211);
  not GNAME6211(G6211,G410);
  dff DFF_6213(CK,G6212,G6208);
  and GNAME6214(G6214,G6212,G6215);
  nand GNAME6215(G6215,G80,G6217);
  buf GNAME6216(G6216,G6212);
  buf GNAME6217(G6217,G6199);
  or GNAME6229(G6229,G6231,G6230);
  and GNAME6230(G6230,G11534,G410);
  and GNAME6231(G6231,G6233,G6232);
  not GNAME6232(G6232,G410);
  dff DFF_6234(CK,G6233,G6229);
  and GNAME6235(G6235,G6233,G6236);
  nand GNAME6236(G6236,G80,G6238);
  buf GNAME6237(G6237,G6233);
  buf GNAME6238(G6238,G6220);
  or GNAME6250(G6250,G6252,G6251);
  and GNAME6251(G6251,G11533,G410);
  and GNAME6252(G6252,G6254,G6253);
  not GNAME6253(G6253,G410);
  dff DFF_6255(CK,G6254,G6250);
  and GNAME6256(G6256,G6254,G6257);
  nand GNAME6257(G6257,G80,G6259);
  buf GNAME6258(G6258,G6254);
  buf GNAME6259(G6259,G6241);
  or GNAME6271(G6271,G6273,G6272);
  and GNAME6272(G6272,G11532,G410);
  and GNAME6273(G6273,G6275,G6274);
  not GNAME6274(G6274,G410);
  dff DFF_6276(CK,G6275,G6271);
  and GNAME6277(G6277,G6275,G6278);
  nand GNAME6278(G6278,G80,G6280);
  buf GNAME6279(G6279,G6275);
  buf GNAME6280(G6280,G6262);
  or GNAME6292(G6292,G6294,G6293);
  and GNAME6293(G6293,G11531,G410);
  and GNAME6294(G6294,G6296,G6295);
  not GNAME6295(G6295,G410);
  dff DFF_6297(CK,G6296,G6292);
  and GNAME6298(G6298,G6296,G6299);
  nand GNAME6299(G6299,G80,G6301);
  buf GNAME6300(G6300,G6296);
  buf GNAME6301(G6301,G6283);
  or GNAME6353(G6353,G6355,G6354);
  and GNAME6354(G6354,G11538,G409);
  and GNAME6355(G6355,G6357,G6356);
  not GNAME6356(G6356,G409);
  dff DFF_6358(CK,G6357,G6353);
  and GNAME6359(G6359,G6357,G6360);
  nand GNAME6360(G6360,G80,G6362);
  buf GNAME6361(G6361,G6357);
  buf GNAME6362(G6362,G6344);
  or GNAME6374(G6374,G6376,G6375);
  and GNAME6375(G6375,G11537,G409);
  and GNAME6376(G6376,G6378,G6377);
  not GNAME6377(G6377,G409);
  dff DFF_6379(CK,G6378,G6374);
  and GNAME6380(G6380,G6378,G6381);
  nand GNAME6381(G6381,G80,G6383);
  buf GNAME6382(G6382,G6378);
  buf GNAME6383(G6383,G6365);
  or GNAME6395(G6395,G6397,G6396);
  and GNAME6396(G6396,G11536,G409);
  and GNAME6397(G6397,G6399,G6398);
  not GNAME6398(G6398,G409);
  dff DFF_6400(CK,G6399,G6395);
  and GNAME6401(G6401,G6399,G6402);
  nand GNAME6402(G6402,G80,G6404);
  buf GNAME6403(G6403,G6399);
  buf GNAME6404(G6404,G6386);
  or GNAME6416(G6416,G6418,G6417);
  and GNAME6417(G6417,G11535,G409);
  and GNAME6418(G6418,G6420,G6419);
  not GNAME6419(G6419,G409);
  dff DFF_6421(CK,G6420,G6416);
  and GNAME6422(G6422,G6420,G6423);
  nand GNAME6423(G6423,G80,G6425);
  buf GNAME6424(G6424,G6420);
  buf GNAME6425(G6425,G6407);
  or GNAME6437(G6437,G6439,G6438);
  and GNAME6438(G6438,G11534,G409);
  and GNAME6439(G6439,G6441,G6440);
  not GNAME6440(G6440,G409);
  dff DFF_6442(CK,G6441,G6437);
  and GNAME6443(G6443,G6441,G6444);
  nand GNAME6444(G6444,G80,G6446);
  buf GNAME6445(G6445,G6441);
  buf GNAME6446(G6446,G6428);
  or GNAME6458(G6458,G6460,G6459);
  and GNAME6459(G6459,G11533,G409);
  and GNAME6460(G6460,G6462,G6461);
  not GNAME6461(G6461,G409);
  dff DFF_6463(CK,G6462,G6458);
  and GNAME6464(G6464,G6462,G6465);
  nand GNAME6465(G6465,G80,G6467);
  buf GNAME6466(G6466,G6462);
  buf GNAME6467(G6467,G6449);
  or GNAME6479(G6479,G6481,G6480);
  and GNAME6480(G6480,G11532,G409);
  and GNAME6481(G6481,G6483,G6482);
  not GNAME6482(G6482,G409);
  dff DFF_6484(CK,G6483,G6479);
  and GNAME6485(G6485,G6483,G6486);
  nand GNAME6486(G6486,G80,G6488);
  buf GNAME6487(G6487,G6483);
  buf GNAME6488(G6488,G6470);
  or GNAME6500(G6500,G6502,G6501);
  and GNAME6501(G6501,G11531,G409);
  and GNAME6502(G6502,G6504,G6503);
  not GNAME6503(G6503,G409);
  dff DFF_6505(CK,G6504,G6500);
  and GNAME6506(G6506,G6504,G6507);
  nand GNAME6507(G6507,G80,G6509);
  buf GNAME6508(G6508,G6504);
  buf GNAME6509(G6509,G6491);
  or GNAME6561(G6561,G6563,G6562);
  and GNAME6562(G6562,G11530,G408);
  and GNAME6563(G6563,G6565,G6564);
  not GNAME6564(G6564,G408);
  dff DFF_6566(CK,G6565,G6561);
  and GNAME6567(G6567,G6565,G6568);
  nand GNAME6568(G6568,G80,G6570);
  buf GNAME6569(G6569,G6565);
  buf GNAME6570(G6570,G6552);
  or GNAME6582(G6582,G6584,G6583);
  and GNAME6583(G6583,G11537,G408);
  and GNAME6584(G6584,G6586,G6585);
  not GNAME6585(G6585,G408);
  dff DFF_6587(CK,G6586,G6582);
  and GNAME6588(G6588,G6586,G6589);
  nand GNAME6589(G6589,G80,G6591);
  buf GNAME6590(G6590,G6586);
  buf GNAME6591(G6591,G6573);
  or GNAME6603(G6603,G6605,G6604);
  and GNAME6604(G6604,G11536,G408);
  and GNAME6605(G6605,G6607,G6606);
  not GNAME6606(G6606,G408);
  dff DFF_6608(CK,G6607,G6603);
  and GNAME6609(G6609,G6607,G6610);
  nand GNAME6610(G6610,G80,G6612);
  buf GNAME6611(G6611,G6607);
  buf GNAME6612(G6612,G6594);
  or GNAME6624(G6624,G6626,G6625);
  and GNAME6625(G6625,G11535,G408);
  and GNAME6626(G6626,G6628,G6627);
  not GNAME6627(G6627,G408);
  dff DFF_6629(CK,G6628,G6624);
  and GNAME6630(G6630,G6628,G6631);
  nand GNAME6631(G6631,G80,G6633);
  buf GNAME6632(G6632,G6628);
  buf GNAME6633(G6633,G6615);
  or GNAME6645(G6645,G6647,G6646);
  and GNAME6646(G6646,G11534,G408);
  and GNAME6647(G6647,G6649,G6648);
  not GNAME6648(G6648,G408);
  dff DFF_6650(CK,G6649,G6645);
  and GNAME6651(G6651,G6649,G6652);
  nand GNAME6652(G6652,G80,G6654);
  buf GNAME6653(G6653,G6649);
  buf GNAME6654(G6654,G6636);
  or GNAME6666(G6666,G6668,G6667);
  and GNAME6667(G6667,G11533,G408);
  and GNAME6668(G6668,G6670,G6669);
  not GNAME6669(G6669,G408);
  dff DFF_6671(CK,G6670,G6666);
  and GNAME6672(G6672,G6670,G6673);
  nand GNAME6673(G6673,G80,G6675);
  buf GNAME6674(G6674,G6670);
  buf GNAME6675(G6675,G6657);
  or GNAME6687(G6687,G6689,G6688);
  and GNAME6688(G6688,G11532,G408);
  and GNAME6689(G6689,G6691,G6690);
  not GNAME6690(G6690,G408);
  dff DFF_6692(CK,G6691,G6687);
  and GNAME6693(G6693,G6691,G6694);
  nand GNAME6694(G6694,G80,G6696);
  buf GNAME6695(G6695,G6691);
  buf GNAME6696(G6696,G6678);
  or GNAME6708(G6708,G6710,G6709);
  and GNAME6709(G6709,G11531,G408);
  and GNAME6710(G6710,G6712,G6711);
  not GNAME6711(G6711,G408);
  dff DFF_6713(CK,G6712,G6708);
  and GNAME6714(G6714,G6712,G6715);
  nand GNAME6715(G6715,G80,G6717);
  buf GNAME6716(G6716,G6712);
  buf GNAME6717(G6717,G6699);
  or GNAME6769(G6769,G6771,G6770);
  and GNAME6770(G6770,G11530,G427);
  and GNAME6771(G6771,G6773,G6772);
  not GNAME6772(G6772,G427);
  dff DFF_6774(CK,G6773,G6769);
  and GNAME6775(G6775,G6773,G6776);
  nand GNAME6776(G6776,G80,G6778);
  buf GNAME6777(G6777,G6773);
  buf GNAME6778(G6778,G6760);
  or GNAME6790(G6790,G6792,G6791);
  and GNAME6791(G6791,G11529,G427);
  and GNAME6792(G6792,G6794,G6793);
  not GNAME6793(G6793,G427);
  dff DFF_6795(CK,G6794,G6790);
  and GNAME6796(G6796,G6794,G6797);
  nand GNAME6797(G6797,G80,G6799);
  buf GNAME6798(G6798,G6794);
  buf GNAME6799(G6799,G6781);
  or GNAME6811(G6811,G6813,G6812);
  and GNAME6812(G6812,G11528,G427);
  and GNAME6813(G6813,G6815,G6814);
  not GNAME6814(G6814,G427);
  dff DFF_6816(CK,G6815,G6811);
  and GNAME6817(G6817,G6815,G6818);
  nand GNAME6818(G6818,G80,G6820);
  buf GNAME6819(G6819,G6815);
  buf GNAME6820(G6820,G6802);
  or GNAME6832(G6832,G6834,G6833);
  and GNAME6833(G6833,G11527,G427);
  and GNAME6834(G6834,G6836,G6835);
  not GNAME6835(G6835,G427);
  dff DFF_6837(CK,G6836,G6832);
  and GNAME6838(G6838,G6836,G6839);
  nand GNAME6839(G6839,G80,G6841);
  buf GNAME6840(G6840,G6836);
  buf GNAME6841(G6841,G6823);
  or GNAME6853(G6853,G6855,G6854);
  and GNAME6854(G6854,G11526,G427);
  and GNAME6855(G6855,G6857,G6856);
  not GNAME6856(G6856,G427);
  dff DFF_6858(CK,G6857,G6853);
  and GNAME6859(G6859,G6857,G6860);
  nand GNAME6860(G6860,G80,G6862);
  buf GNAME6861(G6861,G6857);
  buf GNAME6862(G6862,G6844);
  or GNAME6874(G6874,G6876,G6875);
  and GNAME6875(G6875,G11525,G427);
  and GNAME6876(G6876,G6878,G6877);
  not GNAME6877(G6877,G427);
  dff DFF_6879(CK,G6878,G6874);
  and GNAME6880(G6880,G6878,G6881);
  nand GNAME6881(G6881,G80,G6883);
  buf GNAME6882(G6882,G6878);
  buf GNAME6883(G6883,G6865);
  or GNAME6895(G6895,G6897,G6896);
  and GNAME6896(G6896,G11524,G427);
  and GNAME6897(G6897,G6899,G6898);
  not GNAME6898(G6898,G427);
  dff DFF_6900(CK,G6899,G6895);
  and GNAME6901(G6901,G6899,G6902);
  nand GNAME6902(G6902,G80,G6904);
  buf GNAME6903(G6903,G6899);
  buf GNAME6904(G6904,G6886);
  or GNAME6916(G6916,G6918,G6917);
  and GNAME6917(G6917,G11523,G427);
  and GNAME6918(G6918,G6920,G6919);
  not GNAME6919(G6919,G427);
  dff DFF_6921(CK,G6920,G6916);
  and GNAME6922(G6922,G6920,G6923);
  nand GNAME6923(G6923,G80,G6925);
  buf GNAME6924(G6924,G6920);
  buf GNAME6925(G6925,G6907);
  or GNAME6977(G6977,G6979,G6978);
  and GNAME6978(G6978,G11530,G426);
  and GNAME6979(G6979,G6981,G6980);
  not GNAME6980(G6980,G426);
  dff DFF_6982(CK,G6981,G6977);
  and GNAME6983(G6983,G6981,G6984);
  nand GNAME6984(G6984,G80,G6986);
  buf GNAME6985(G6985,G6981);
  buf GNAME6986(G6986,G6968);
  or GNAME6998(G6998,G7000,G6999);
  and GNAME6999(G6999,G11529,G426);
  and GNAME7000(G7000,G7002,G7001);
  not GNAME7001(G7001,G426);
  dff DFF_7003(CK,G7002,G6998);
  and GNAME7004(G7004,G7002,G7005);
  nand GNAME7005(G7005,G80,G7007);
  buf GNAME7006(G7006,G7002);
  buf GNAME7007(G7007,G6989);
  or GNAME7019(G7019,G7021,G7020);
  and GNAME7020(G7020,G11528,G426);
  and GNAME7021(G7021,G7023,G7022);
  not GNAME7022(G7022,G426);
  dff DFF_7024(CK,G7023,G7019);
  and GNAME7025(G7025,G7023,G7026);
  nand GNAME7026(G7026,G80,G7028);
  buf GNAME7027(G7027,G7023);
  buf GNAME7028(G7028,G7010);
  or GNAME7040(G7040,G7042,G7041);
  and GNAME7041(G7041,G11527,G426);
  and GNAME7042(G7042,G7044,G7043);
  not GNAME7043(G7043,G426);
  dff DFF_7045(CK,G7044,G7040);
  and GNAME7046(G7046,G7044,G7047);
  nand GNAME7047(G7047,G80,G7049);
  buf GNAME7048(G7048,G7044);
  buf GNAME7049(G7049,G7031);
  or GNAME7061(G7061,G7063,G7062);
  and GNAME7062(G7062,G11526,G426);
  and GNAME7063(G7063,G7065,G7064);
  not GNAME7064(G7064,G426);
  dff DFF_7066(CK,G7065,G7061);
  and GNAME7067(G7067,G7065,G7068);
  nand GNAME7068(G7068,G80,G7070);
  buf GNAME7069(G7069,G7065);
  buf GNAME7070(G7070,G7052);
  or GNAME7082(G7082,G7084,G7083);
  and GNAME7083(G7083,G11525,G426);
  and GNAME7084(G7084,G7086,G7085);
  not GNAME7085(G7085,G426);
  dff DFF_7087(CK,G7086,G7082);
  and GNAME7088(G7088,G7086,G7089);
  nand GNAME7089(G7089,G80,G7091);
  buf GNAME7090(G7090,G7086);
  buf GNAME7091(G7091,G7073);
  or GNAME7103(G7103,G7105,G7104);
  and GNAME7104(G7104,G11524,G426);
  and GNAME7105(G7105,G7107,G7106);
  not GNAME7106(G7106,G426);
  dff DFF_7108(CK,G7107,G7103);
  and GNAME7109(G7109,G7107,G7110);
  nand GNAME7110(G7110,G80,G7112);
  buf GNAME7111(G7111,G7107);
  buf GNAME7112(G7112,G7094);
  or GNAME7124(G7124,G7126,G7125);
  and GNAME7125(G7125,G11523,G426);
  and GNAME7126(G7126,G7128,G7127);
  not GNAME7127(G7127,G426);
  dff DFF_7129(CK,G7128,G7124);
  and GNAME7130(G7130,G7128,G7131);
  nand GNAME7131(G7131,G80,G7133);
  buf GNAME7132(G7132,G7128);
  buf GNAME7133(G7133,G7115);
  or GNAME7185(G7185,G7187,G7186);
  and GNAME7186(G7186,G11530,G425);
  and GNAME7187(G7187,G7189,G7188);
  not GNAME7188(G7188,G425);
  dff DFF_7190(CK,G7189,G7185);
  and GNAME7191(G7191,G7189,G7192);
  nand GNAME7192(G7192,G80,G7194);
  buf GNAME7193(G7193,G7189);
  buf GNAME7194(G7194,G7176);
  or GNAME7206(G7206,G7208,G7207);
  and GNAME7207(G7207,G11529,G425);
  and GNAME7208(G7208,G7210,G7209);
  not GNAME7209(G7209,G425);
  dff DFF_7211(CK,G7210,G7206);
  and GNAME7212(G7212,G7210,G7213);
  nand GNAME7213(G7213,G80,G7215);
  buf GNAME7214(G7214,G7210);
  buf GNAME7215(G7215,G7197);
  or GNAME7227(G7227,G7229,G7228);
  and GNAME7228(G7228,G11528,G425);
  and GNAME7229(G7229,G7231,G7230);
  not GNAME7230(G7230,G425);
  dff DFF_7232(CK,G7231,G7227);
  and GNAME7233(G7233,G7231,G7234);
  nand GNAME7234(G7234,G80,G7236);
  buf GNAME7235(G7235,G7231);
  buf GNAME7236(G7236,G7218);
  or GNAME7248(G7248,G7250,G7249);
  and GNAME7249(G7249,G11527,G425);
  and GNAME7250(G7250,G7252,G7251);
  not GNAME7251(G7251,G425);
  dff DFF_7253(CK,G7252,G7248);
  and GNAME7254(G7254,G7252,G7255);
  nand GNAME7255(G7255,G80,G7257);
  buf GNAME7256(G7256,G7252);
  buf GNAME7257(G7257,G7239);
  or GNAME7269(G7269,G7271,G7270);
  and GNAME7270(G7270,G11526,G425);
  and GNAME7271(G7271,G7273,G7272);
  not GNAME7272(G7272,G425);
  dff DFF_7274(CK,G7273,G7269);
  and GNAME7275(G7275,G7273,G7276);
  nand GNAME7276(G7276,G80,G7278);
  buf GNAME7277(G7277,G7273);
  buf GNAME7278(G7278,G7260);
  or GNAME7290(G7290,G7292,G7291);
  and GNAME7291(G7291,G11525,G425);
  and GNAME7292(G7292,G7294,G7293);
  not GNAME7293(G7293,G425);
  dff DFF_7295(CK,G7294,G7290);
  and GNAME7296(G7296,G7294,G7297);
  nand GNAME7297(G7297,G80,G7299);
  buf GNAME7298(G7298,G7294);
  buf GNAME7299(G7299,G7281);
  or GNAME7311(G7311,G7313,G7312);
  and GNAME7312(G7312,G11524,G425);
  and GNAME7313(G7313,G7315,G7314);
  not GNAME7314(G7314,G425);
  dff DFF_7316(CK,G7315,G7311);
  and GNAME7317(G7317,G7315,G7318);
  nand GNAME7318(G7318,G80,G7320);
  buf GNAME7319(G7319,G7315);
  buf GNAME7320(G7320,G7302);
  or GNAME7332(G7332,G7334,G7333);
  and GNAME7333(G7333,G11523,G425);
  and GNAME7334(G7334,G7336,G7335);
  not GNAME7335(G7335,G425);
  dff DFF_7337(CK,G7336,G7332);
  and GNAME7338(G7338,G7336,G7339);
  nand GNAME7339(G7339,G80,G7341);
  buf GNAME7340(G7340,G7336);
  buf GNAME7341(G7341,G7323);
  or GNAME7393(G7393,G7395,G7394);
  and GNAME7394(G7394,G11530,G424);
  and GNAME7395(G7395,G7397,G7396);
  not GNAME7396(G7396,G424);
  dff DFF_7398(CK,G7397,G7393);
  and GNAME7399(G7399,G7397,G7400);
  nand GNAME7400(G7400,G80,G7402);
  buf GNAME7401(G7401,G7397);
  buf GNAME7402(G7402,G7384);
  or GNAME7414(G7414,G7416,G7415);
  and GNAME7415(G7415,G11529,G424);
  and GNAME7416(G7416,G7418,G7417);
  not GNAME7417(G7417,G424);
  dff DFF_7419(CK,G7418,G7414);
  and GNAME7420(G7420,G7418,G7421);
  nand GNAME7421(G7421,G80,G7423);
  buf GNAME7422(G7422,G7418);
  buf GNAME7423(G7423,G7405);
  or GNAME7435(G7435,G7437,G7436);
  and GNAME7436(G7436,G11528,G424);
  and GNAME7437(G7437,G7439,G7438);
  not GNAME7438(G7438,G424);
  dff DFF_7440(CK,G7439,G7435);
  and GNAME7441(G7441,G7439,G7442);
  nand GNAME7442(G7442,G80,G7444);
  buf GNAME7443(G7443,G7439);
  buf GNAME7444(G7444,G7426);
  or GNAME7456(G7456,G7458,G7457);
  and GNAME7457(G7457,G11527,G424);
  and GNAME7458(G7458,G7460,G7459);
  not GNAME7459(G7459,G424);
  dff DFF_7461(CK,G7460,G7456);
  and GNAME7462(G7462,G7460,G7463);
  nand GNAME7463(G7463,G80,G7465);
  buf GNAME7464(G7464,G7460);
  buf GNAME7465(G7465,G7447);
  or GNAME7477(G7477,G7479,G7478);
  and GNAME7478(G7478,G11526,G424);
  and GNAME7479(G7479,G7481,G7480);
  not GNAME7480(G7480,G424);
  dff DFF_7482(CK,G7481,G7477);
  and GNAME7483(G7483,G7481,G7484);
  nand GNAME7484(G7484,G80,G7486);
  buf GNAME7485(G7485,G7481);
  buf GNAME7486(G7486,G7468);
  or GNAME7498(G7498,G7500,G7499);
  and GNAME7499(G7499,G11525,G424);
  and GNAME7500(G7500,G7502,G7501);
  not GNAME7501(G7501,G424);
  dff DFF_7503(CK,G7502,G7498);
  and GNAME7504(G7504,G7502,G7505);
  nand GNAME7505(G7505,G80,G7507);
  buf GNAME7506(G7506,G7502);
  buf GNAME7507(G7507,G7489);
  or GNAME7519(G7519,G7521,G7520);
  and GNAME7520(G7520,G11524,G424);
  and GNAME7521(G7521,G7523,G7522);
  not GNAME7522(G7522,G424);
  dff DFF_7524(CK,G7523,G7519);
  and GNAME7525(G7525,G7523,G7526);
  nand GNAME7526(G7526,G80,G7528);
  buf GNAME7527(G7527,G7523);
  buf GNAME7528(G7528,G7510);
  or GNAME7540(G7540,G7542,G7541);
  and GNAME7541(G7541,G11523,G424);
  and GNAME7542(G7542,G7544,G7543);
  not GNAME7543(G7543,G424);
  dff DFF_7545(CK,G7544,G7540);
  and GNAME7546(G7546,G7544,G7547);
  nand GNAME7547(G7547,G80,G7549);
  buf GNAME7548(G7548,G7544);
  buf GNAME7549(G7549,G7531);
  or GNAME7601(G7601,G7603,G7602);
  and GNAME7602(G7602,G11530,G423);
  and GNAME7603(G7603,G7605,G7604);
  not GNAME7604(G7604,G423);
  dff DFF_7606(CK,G7605,G7601);
  and GNAME7607(G7607,G7605,G7608);
  nand GNAME7608(G7608,G80,G7610);
  buf GNAME7609(G7609,G7605);
  buf GNAME7610(G7610,G7592);
  or GNAME7622(G7622,G7624,G7623);
  and GNAME7623(G7623,G11529,G423);
  and GNAME7624(G7624,G7626,G7625);
  not GNAME7625(G7625,G423);
  dff DFF_7627(CK,G7626,G7622);
  and GNAME7628(G7628,G7626,G7629);
  nand GNAME7629(G7629,G80,G7631);
  buf GNAME7630(G7630,G7626);
  buf GNAME7631(G7631,G7613);
  or GNAME7643(G7643,G7645,G7644);
  and GNAME7644(G7644,G11528,G423);
  and GNAME7645(G7645,G7647,G7646);
  not GNAME7646(G7646,G423);
  dff DFF_7648(CK,G7647,G7643);
  and GNAME7649(G7649,G7647,G7650);
  nand GNAME7650(G7650,G80,G7652);
  buf GNAME7651(G7651,G7647);
  buf GNAME7652(G7652,G7634);
  or GNAME7664(G7664,G7666,G7665);
  and GNAME7665(G7665,G11527,G423);
  and GNAME7666(G7666,G7668,G7667);
  not GNAME7667(G7667,G423);
  dff DFF_7669(CK,G7668,G7664);
  and GNAME7670(G7670,G7668,G7671);
  nand GNAME7671(G7671,G80,G7673);
  buf GNAME7672(G7672,G7668);
  buf GNAME7673(G7673,G7655);
  or GNAME7685(G7685,G7687,G7686);
  and GNAME7686(G7686,G11526,G423);
  and GNAME7687(G7687,G7689,G7688);
  not GNAME7688(G7688,G423);
  dff DFF_7690(CK,G7689,G7685);
  and GNAME7691(G7691,G7689,G7692);
  nand GNAME7692(G7692,G80,G7694);
  buf GNAME7693(G7693,G7689);
  buf GNAME7694(G7694,G7676);
  or GNAME7706(G7706,G7708,G7707);
  and GNAME7707(G7707,G11525,G423);
  and GNAME7708(G7708,G7710,G7709);
  not GNAME7709(G7709,G423);
  dff DFF_7711(CK,G7710,G7706);
  and GNAME7712(G7712,G7710,G7713);
  nand GNAME7713(G7713,G80,G7715);
  buf GNAME7714(G7714,G7710);
  buf GNAME7715(G7715,G7697);
  or GNAME7727(G7727,G7729,G7728);
  and GNAME7728(G7728,G11524,G423);
  and GNAME7729(G7729,G7731,G7730);
  not GNAME7730(G7730,G423);
  dff DFF_7732(CK,G7731,G7727);
  and GNAME7733(G7733,G7731,G7734);
  nand GNAME7734(G7734,G80,G7736);
  buf GNAME7735(G7735,G7731);
  buf GNAME7736(G7736,G7718);
  or GNAME7748(G7748,G7750,G7749);
  and GNAME7749(G7749,G11523,G423);
  and GNAME7750(G7750,G7752,G7751);
  not GNAME7751(G7751,G423);
  dff DFF_7753(CK,G7752,G7748);
  and GNAME7754(G7754,G7752,G7755);
  nand GNAME7755(G7755,G80,G7757);
  buf GNAME7756(G7756,G7752);
  buf GNAME7757(G7757,G7739);
  or GNAME7809(G7809,G7811,G7810);
  and GNAME7810(G7810,G11530,G422);
  and GNAME7811(G7811,G7813,G7812);
  not GNAME7812(G7812,G422);
  dff DFF_7814(CK,G7813,G7809);
  and GNAME7815(G7815,G7813,G7816);
  nand GNAME7816(G7816,G80,G7818);
  buf GNAME7817(G7817,G7813);
  buf GNAME7818(G7818,G7800);
  or GNAME7830(G7830,G7832,G7831);
  and GNAME7831(G7831,G11529,G422);
  and GNAME7832(G7832,G7834,G7833);
  not GNAME7833(G7833,G422);
  dff DFF_7835(CK,G7834,G7830);
  and GNAME7836(G7836,G7834,G7837);
  nand GNAME7837(G7837,G80,G7839);
  buf GNAME7838(G7838,G7834);
  buf GNAME7839(G7839,G7821);
  or GNAME7851(G7851,G7853,G7852);
  and GNAME7852(G7852,G11528,G422);
  and GNAME7853(G7853,G7855,G7854);
  not GNAME7854(G7854,G422);
  dff DFF_7856(CK,G7855,G7851);
  and GNAME7857(G7857,G7855,G7858);
  nand GNAME7858(G7858,G80,G7860);
  buf GNAME7859(G7859,G7855);
  buf GNAME7860(G7860,G7842);
  or GNAME7872(G7872,G7874,G7873);
  and GNAME7873(G7873,G11527,G422);
  and GNAME7874(G7874,G7876,G7875);
  not GNAME7875(G7875,G422);
  dff DFF_7877(CK,G7876,G7872);
  and GNAME7878(G7878,G7876,G7879);
  nand GNAME7879(G7879,G80,G7881);
  buf GNAME7880(G7880,G7876);
  buf GNAME7881(G7881,G7863);
  or GNAME7893(G7893,G7895,G7894);
  and GNAME7894(G7894,G11526,G422);
  and GNAME7895(G7895,G7897,G7896);
  not GNAME7896(G7896,G422);
  dff DFF_7898(CK,G7897,G7893);
  and GNAME7899(G7899,G7897,G7900);
  nand GNAME7900(G7900,G80,G7902);
  buf GNAME7901(G7901,G7897);
  buf GNAME7902(G7902,G7884);
  or GNAME7914(G7914,G7916,G7915);
  and GNAME7915(G7915,G11525,G422);
  and GNAME7916(G7916,G7918,G7917);
  not GNAME7917(G7917,G422);
  dff DFF_7919(CK,G7918,G7914);
  and GNAME7920(G7920,G7918,G7921);
  nand GNAME7921(G7921,G80,G7923);
  buf GNAME7922(G7922,G7918);
  buf GNAME7923(G7923,G7905);
  or GNAME7935(G7935,G7937,G7936);
  and GNAME7936(G7936,G11524,G422);
  and GNAME7937(G7937,G7939,G7938);
  not GNAME7938(G7938,G422);
  dff DFF_7940(CK,G7939,G7935);
  and GNAME7941(G7941,G7939,G7942);
  nand GNAME7942(G7942,G80,G7944);
  buf GNAME7943(G7943,G7939);
  buf GNAME7944(G7944,G7926);
  or GNAME7956(G7956,G7958,G7957);
  and GNAME7957(G7957,G11523,G422);
  and GNAME7958(G7958,G7960,G7959);
  not GNAME7959(G7959,G422);
  dff DFF_7961(CK,G7960,G7956);
  and GNAME7962(G7962,G7960,G7963);
  nand GNAME7963(G7963,G80,G7965);
  buf GNAME7964(G7964,G7960);
  buf GNAME7965(G7965,G7947);
  or GNAME8017(G8017,G8019,G8018);
  and GNAME8018(G8018,G11530,G421);
  and GNAME8019(G8019,G8021,G8020);
  not GNAME8020(G8020,G421);
  dff DFF_8022(CK,G8021,G8017);
  and GNAME8023(G8023,G8021,G8024);
  nand GNAME8024(G8024,G80,G8026);
  buf GNAME8025(G8025,G8021);
  buf GNAME8026(G8026,G8008);
  or GNAME8038(G8038,G8040,G8039);
  and GNAME8039(G8039,G11529,G421);
  and GNAME8040(G8040,G8042,G8041);
  not GNAME8041(G8041,G421);
  dff DFF_8043(CK,G8042,G8038);
  and GNAME8044(G8044,G8042,G8045);
  nand GNAME8045(G8045,G80,G8047);
  buf GNAME8046(G8046,G8042);
  buf GNAME8047(G8047,G8029);
  or GNAME8059(G8059,G8061,G8060);
  and GNAME8060(G8060,G11528,G421);
  and GNAME8061(G8061,G8063,G8062);
  not GNAME8062(G8062,G421);
  dff DFF_8064(CK,G8063,G8059);
  and GNAME8065(G8065,G8063,G8066);
  nand GNAME8066(G8066,G80,G8068);
  buf GNAME8067(G8067,G8063);
  buf GNAME8068(G8068,G8050);
  or GNAME8080(G8080,G8082,G8081);
  and GNAME8081(G8081,G11527,G421);
  and GNAME8082(G8082,G8084,G8083);
  not GNAME8083(G8083,G421);
  dff DFF_8085(CK,G8084,G8080);
  and GNAME8086(G8086,G8084,G8087);
  nand GNAME8087(G8087,G80,G8089);
  buf GNAME8088(G8088,G8084);
  buf GNAME8089(G8089,G8071);
  or GNAME8101(G8101,G8103,G8102);
  and GNAME8102(G8102,G11526,G421);
  and GNAME8103(G8103,G8105,G8104);
  not GNAME8104(G8104,G421);
  dff DFF_8106(CK,G8105,G8101);
  and GNAME8107(G8107,G8105,G8108);
  nand GNAME8108(G8108,G80,G8110);
  buf GNAME8109(G8109,G8105);
  buf GNAME8110(G8110,G8092);
  or GNAME8122(G8122,G8124,G8123);
  and GNAME8123(G8123,G11525,G421);
  and GNAME8124(G8124,G8126,G8125);
  not GNAME8125(G8125,G421);
  dff DFF_8127(CK,G8126,G8122);
  and GNAME8128(G8128,G8126,G8129);
  nand GNAME8129(G8129,G80,G8131);
  buf GNAME8130(G8130,G8126);
  buf GNAME8131(G8131,G8113);
  or GNAME8143(G8143,G8145,G8144);
  and GNAME8144(G8144,G11524,G421);
  and GNAME8145(G8145,G8147,G8146);
  not GNAME8146(G8146,G421);
  dff DFF_8148(CK,G8147,G8143);
  and GNAME8149(G8149,G8147,G8150);
  nand GNAME8150(G8150,G80,G8152);
  buf GNAME8151(G8151,G8147);
  buf GNAME8152(G8152,G8134);
  or GNAME8164(G8164,G8166,G8165);
  and GNAME8165(G8165,G11523,G421);
  and GNAME8166(G8166,G8168,G8167);
  not GNAME8167(G8167,G421);
  dff DFF_8169(CK,G8168,G8164);
  and GNAME8170(G8170,G8168,G8171);
  nand GNAME8171(G8171,G80,G8173);
  buf GNAME8172(G8172,G8168);
  buf GNAME8173(G8173,G8155);
  or GNAME8225(G8225,G8227,G8226);
  and GNAME8226(G8226,G11530,G420);
  and GNAME8227(G8227,G8229,G8228);
  not GNAME8228(G8228,G420);
  dff DFF_8230(CK,G8229,G8225);
  and GNAME8231(G8231,G8229,G8232);
  nand GNAME8232(G8232,G80,G8234);
  buf GNAME8233(G8233,G8229);
  buf GNAME8234(G8234,G8216);
  or GNAME8246(G8246,G8248,G8247);
  and GNAME8247(G8247,G11529,G420);
  and GNAME8248(G8248,G8250,G8249);
  not GNAME8249(G8249,G420);
  dff DFF_8251(CK,G8250,G8246);
  and GNAME8252(G8252,G8250,G8253);
  nand GNAME8253(G8253,G80,G8255);
  buf GNAME8254(G8254,G8250);
  buf GNAME8255(G8255,G8237);
  or GNAME8267(G8267,G8269,G8268);
  and GNAME8268(G8268,G11528,G420);
  and GNAME8269(G8269,G8271,G8270);
  not GNAME8270(G8270,G420);
  dff DFF_8272(CK,G8271,G8267);
  and GNAME8273(G8273,G8271,G8274);
  nand GNAME8274(G8274,G80,G8276);
  buf GNAME8275(G8275,G8271);
  buf GNAME8276(G8276,G8258);
  or GNAME8288(G8288,G8290,G8289);
  and GNAME8289(G8289,G11527,G420);
  and GNAME8290(G8290,G8292,G8291);
  not GNAME8291(G8291,G420);
  dff DFF_8293(CK,G8292,G8288);
  and GNAME8294(G8294,G8292,G8295);
  nand GNAME8295(G8295,G80,G8297);
  buf GNAME8296(G8296,G8292);
  buf GNAME8297(G8297,G8279);
  or GNAME8309(G8309,G8311,G8310);
  and GNAME8310(G8310,G11526,G420);
  and GNAME8311(G8311,G8313,G8312);
  not GNAME8312(G8312,G420);
  dff DFF_8314(CK,G8313,G8309);
  and GNAME8315(G8315,G8313,G8316);
  nand GNAME8316(G8316,G80,G8318);
  buf GNAME8317(G8317,G8313);
  buf GNAME8318(G8318,G8300);
  or GNAME8330(G8330,G8332,G8331);
  and GNAME8331(G8331,G11525,G420);
  and GNAME8332(G8332,G8334,G8333);
  not GNAME8333(G8333,G420);
  dff DFF_8335(CK,G8334,G8330);
  and GNAME8336(G8336,G8334,G8337);
  nand GNAME8337(G8337,G80,G8339);
  buf GNAME8338(G8338,G8334);
  buf GNAME8339(G8339,G8321);
  or GNAME8351(G8351,G8353,G8352);
  and GNAME8352(G8352,G11524,G420);
  and GNAME8353(G8353,G8355,G8354);
  not GNAME8354(G8354,G420);
  dff DFF_8356(CK,G8355,G8351);
  and GNAME8357(G8357,G8355,G8358);
  nand GNAME8358(G8358,G80,G8360);
  buf GNAME8359(G8359,G8355);
  buf GNAME8360(G8360,G8342);
  or GNAME8372(G8372,G8374,G8373);
  and GNAME8373(G8373,G11523,G420);
  and GNAME8374(G8374,G8376,G8375);
  not GNAME8375(G8375,G420);
  dff DFF_8377(CK,G8376,G8372);
  and GNAME8378(G8378,G8376,G8379);
  nand GNAME8379(G8379,G80,G8381);
  buf GNAME8380(G8380,G8376);
  buf GNAME8381(G8381,G8363);
  or GNAME8433(G8433,G8435,G8434);
  and GNAME8434(G8434,G11530,G419);
  and GNAME8435(G8435,G8437,G8436);
  not GNAME8436(G8436,G419);
  dff DFF_8438(CK,G8437,G8433);
  and GNAME8439(G8439,G8437,G8440);
  nand GNAME8440(G8440,G80,G8442);
  buf GNAME8441(G8441,G8437);
  buf GNAME8442(G8442,G8424);
  or GNAME8454(G8454,G8456,G8455);
  and GNAME8455(G8455,G11529,G419);
  and GNAME8456(G8456,G8458,G8457);
  not GNAME8457(G8457,G419);
  dff DFF_8459(CK,G8458,G8454);
  and GNAME8460(G8460,G8458,G8461);
  nand GNAME8461(G8461,G80,G8463);
  buf GNAME8462(G8462,G8458);
  buf GNAME8463(G8463,G8445);
  or GNAME8475(G8475,G8477,G8476);
  and GNAME8476(G8476,G11528,G419);
  and GNAME8477(G8477,G8479,G8478);
  not GNAME8478(G8478,G419);
  dff DFF_8480(CK,G8479,G8475);
  and GNAME8481(G8481,G8479,G8482);
  nand GNAME8482(G8482,G80,G8484);
  buf GNAME8483(G8483,G8479);
  buf GNAME8484(G8484,G8466);
  or GNAME8496(G8496,G8498,G8497);
  and GNAME8497(G8497,G11527,G419);
  and GNAME8498(G8498,G8500,G8499);
  not GNAME8499(G8499,G419);
  dff DFF_8501(CK,G8500,G8496);
  and GNAME8502(G8502,G8500,G8503);
  nand GNAME8503(G8503,G80,G8505);
  buf GNAME8504(G8504,G8500);
  buf GNAME8505(G8505,G8487);
  or GNAME8517(G8517,G8519,G8518);
  and GNAME8518(G8518,G11526,G419);
  and GNAME8519(G8519,G8521,G8520);
  not GNAME8520(G8520,G419);
  dff DFF_8522(CK,G8521,G8517);
  and GNAME8523(G8523,G8521,G8524);
  nand GNAME8524(G8524,G80,G8526);
  buf GNAME8525(G8525,G8521);
  buf GNAME8526(G8526,G8508);
  or GNAME8538(G8538,G8540,G8539);
  and GNAME8539(G8539,G11525,G419);
  and GNAME8540(G8540,G8542,G8541);
  not GNAME8541(G8541,G419);
  dff DFF_8543(CK,G8542,G8538);
  and GNAME8544(G8544,G8542,G8545);
  nand GNAME8545(G8545,G80,G8547);
  buf GNAME8546(G8546,G8542);
  buf GNAME8547(G8547,G8529);
  or GNAME8559(G8559,G8561,G8560);
  and GNAME8560(G8560,G11524,G419);
  and GNAME8561(G8561,G8563,G8562);
  not GNAME8562(G8562,G419);
  dff DFF_8564(CK,G8563,G8559);
  and GNAME8565(G8565,G8563,G8566);
  nand GNAME8566(G8566,G80,G8568);
  buf GNAME8567(G8567,G8563);
  buf GNAME8568(G8568,G8550);
  or GNAME8580(G8580,G8582,G8581);
  and GNAME8581(G8581,G11523,G419);
  and GNAME8582(G8582,G8584,G8583);
  not GNAME8583(G8583,G419);
  dff DFF_8585(CK,G8584,G8580);
  and GNAME8586(G8586,G8584,G8587);
  nand GNAME8587(G8587,G80,G8589);
  buf GNAME8588(G8588,G8584);
  buf GNAME8589(G8589,G8571);
  or GNAME8641(G8641,G8643,G8642);
  and GNAME8642(G8642,G11530,G418);
  and GNAME8643(G8643,G8645,G8644);
  not GNAME8644(G8644,G418);
  dff DFF_8646(CK,G8645,G8641);
  and GNAME8647(G8647,G8645,G8648);
  nand GNAME8648(G8648,G80,G8650);
  buf GNAME8649(G8649,G8645);
  buf GNAME8650(G8650,G8632);
  or GNAME8662(G8662,G8664,G8663);
  and GNAME8663(G8663,G11529,G418);
  and GNAME8664(G8664,G8666,G8665);
  not GNAME8665(G8665,G418);
  dff DFF_8667(CK,G8666,G8662);
  and GNAME8668(G8668,G8666,G8669);
  nand GNAME8669(G8669,G80,G8671);
  buf GNAME8670(G8670,G8666);
  buf GNAME8671(G8671,G8653);
  or GNAME8683(G8683,G8685,G8684);
  and GNAME8684(G8684,G11528,G418);
  and GNAME8685(G8685,G8687,G8686);
  not GNAME8686(G8686,G418);
  dff DFF_8688(CK,G8687,G8683);
  and GNAME8689(G8689,G8687,G8690);
  nand GNAME8690(G8690,G80,G8692);
  buf GNAME8691(G8691,G8687);
  buf GNAME8692(G8692,G8674);
  or GNAME8704(G8704,G8706,G8705);
  and GNAME8705(G8705,G11527,G418);
  and GNAME8706(G8706,G8708,G8707);
  not GNAME8707(G8707,G418);
  dff DFF_8709(CK,G8708,G8704);
  and GNAME8710(G8710,G8708,G8711);
  nand GNAME8711(G8711,G80,G8713);
  buf GNAME8712(G8712,G8708);
  buf GNAME8713(G8713,G8695);
  or GNAME8725(G8725,G8727,G8726);
  and GNAME8726(G8726,G11526,G418);
  and GNAME8727(G8727,G8729,G8728);
  not GNAME8728(G8728,G418);
  dff DFF_8730(CK,G8729,G8725);
  and GNAME8731(G8731,G8729,G8732);
  nand GNAME8732(G8732,G80,G8734);
  buf GNAME8733(G8733,G8729);
  buf GNAME8734(G8734,G8716);
  or GNAME8746(G8746,G8748,G8747);
  and GNAME8747(G8747,G11525,G418);
  and GNAME8748(G8748,G8750,G8749);
  not GNAME8749(G8749,G418);
  dff DFF_8751(CK,G8750,G8746);
  and GNAME8752(G8752,G8750,G8753);
  nand GNAME8753(G8753,G80,G8755);
  buf GNAME8754(G8754,G8750);
  buf GNAME8755(G8755,G8737);
  or GNAME8767(G8767,G8769,G8768);
  and GNAME8768(G8768,G11524,G418);
  and GNAME8769(G8769,G8771,G8770);
  not GNAME8770(G8770,G418);
  dff DFF_8772(CK,G8771,G8767);
  and GNAME8773(G8773,G8771,G8774);
  nand GNAME8774(G8774,G80,G8776);
  buf GNAME8775(G8775,G8771);
  buf GNAME8776(G8776,G8758);
  or GNAME8788(G8788,G8790,G8789);
  and GNAME8789(G8789,G11523,G418);
  and GNAME8790(G8790,G8792,G8791);
  not GNAME8791(G8791,G418);
  dff DFF_8793(CK,G8792,G8788);
  and GNAME8794(G8794,G8792,G8795);
  nand GNAME8795(G8795,G80,G8797);
  buf GNAME8796(G8796,G8792);
  buf GNAME8797(G8797,G8779);
  or GNAME8849(G8849,G8851,G8850);
  and GNAME8850(G8850,G11530,G417);
  and GNAME8851(G8851,G8853,G8852);
  not GNAME8852(G8852,G417);
  dff DFF_8854(CK,G8853,G8849);
  and GNAME8855(G8855,G8853,G8856);
  nand GNAME8856(G8856,G80,G8858);
  buf GNAME8857(G8857,G8853);
  buf GNAME8858(G8858,G8840);
  or GNAME8870(G8870,G8872,G8871);
  and GNAME8871(G8871,G11529,G417);
  and GNAME8872(G8872,G8874,G8873);
  not GNAME8873(G8873,G417);
  dff DFF_8875(CK,G8874,G8870);
  and GNAME8876(G8876,G8874,G8877);
  nand GNAME8877(G8877,G80,G8879);
  buf GNAME8878(G8878,G8874);
  buf GNAME8879(G8879,G8861);
  or GNAME8891(G8891,G8893,G8892);
  and GNAME8892(G8892,G11528,G417);
  and GNAME8893(G8893,G8895,G8894);
  not GNAME8894(G8894,G417);
  dff DFF_8896(CK,G8895,G8891);
  and GNAME8897(G8897,G8895,G8898);
  nand GNAME8898(G8898,G80,G8900);
  buf GNAME8899(G8899,G8895);
  buf GNAME8900(G8900,G8882);
  or GNAME8912(G8912,G8914,G8913);
  and GNAME8913(G8913,G11527,G417);
  and GNAME8914(G8914,G8916,G8915);
  not GNAME8915(G8915,G417);
  dff DFF_8917(CK,G8916,G8912);
  and GNAME8918(G8918,G8916,G8919);
  nand GNAME8919(G8919,G80,G8921);
  buf GNAME8920(G8920,G8916);
  buf GNAME8921(G8921,G8903);
  or GNAME8933(G8933,G8935,G8934);
  and GNAME8934(G8934,G11526,G417);
  and GNAME8935(G8935,G8937,G8936);
  not GNAME8936(G8936,G417);
  dff DFF_8938(CK,G8937,G8933);
  and GNAME8939(G8939,G8937,G8940);
  nand GNAME8940(G8940,G80,G8942);
  buf GNAME8941(G8941,G8937);
  buf GNAME8942(G8942,G8924);
  or GNAME8954(G8954,G8956,G8955);
  and GNAME8955(G8955,G11525,G417);
  and GNAME8956(G8956,G8958,G8957);
  not GNAME8957(G8957,G417);
  dff DFF_8959(CK,G8958,G8954);
  and GNAME8960(G8960,G8958,G8961);
  nand GNAME8961(G8961,G80,G8963);
  buf GNAME8962(G8962,G8958);
  buf GNAME8963(G8963,G8945);
  or GNAME8975(G8975,G8977,G8976);
  and GNAME8976(G8976,G11524,G417);
  and GNAME8977(G8977,G8979,G8978);
  not GNAME8978(G8978,G417);
  dff DFF_8980(CK,G8979,G8975);
  and GNAME8981(G8981,G8979,G8982);
  nand GNAME8982(G8982,G80,G8984);
  buf GNAME8983(G8983,G8979);
  buf GNAME8984(G8984,G8966);
  or GNAME8996(G8996,G8998,G8997);
  and GNAME8997(G8997,G11523,G417);
  and GNAME8998(G8998,G9000,G8999);
  not GNAME8999(G8999,G417);
  dff DFF_9001(CK,G9000,G8996);
  and GNAME9002(G9002,G9000,G9003);
  nand GNAME9003(G9003,G80,G9005);
  buf GNAME9004(G9004,G9000);
  buf GNAME9005(G9005,G8987);
  or GNAME9057(G9057,G9059,G9058);
  and GNAME9058(G9058,G11522,G416);
  and GNAME9059(G9059,G9061,G9060);
  not GNAME9060(G9060,G416);
  dff DFF_9062(CK,G9061,G9057);
  and GNAME9063(G9063,G9061,G9064);
  nand GNAME9064(G9064,G80,G9066);
  buf GNAME9065(G9065,G9061);
  buf GNAME9066(G9066,G9048);
  or GNAME9078(G9078,G9080,G9079);
  and GNAME9079(G9079,G11529,G416);
  and GNAME9080(G9080,G9082,G9081);
  not GNAME9081(G9081,G416);
  dff DFF_9083(CK,G9082,G9078);
  and GNAME9084(G9084,G9082,G9085);
  nand GNAME9085(G9085,G80,G9087);
  buf GNAME9086(G9086,G9082);
  buf GNAME9087(G9087,G9069);
  or GNAME9099(G9099,G9101,G9100);
  and GNAME9100(G9100,G11528,G416);
  and GNAME9101(G9101,G9103,G9102);
  not GNAME9102(G9102,G416);
  dff DFF_9104(CK,G9103,G9099);
  and GNAME9105(G9105,G9103,G9106);
  nand GNAME9106(G9106,G80,G9108);
  buf GNAME9107(G9107,G9103);
  buf GNAME9108(G9108,G9090);
  or GNAME9120(G9120,G9122,G9121);
  and GNAME9121(G9121,G11527,G416);
  and GNAME9122(G9122,G9124,G9123);
  not GNAME9123(G9123,G416);
  dff DFF_9125(CK,G9124,G9120);
  and GNAME9126(G9126,G9124,G9127);
  nand GNAME9127(G9127,G80,G9129);
  buf GNAME9128(G9128,G9124);
  buf GNAME9129(G9129,G9111);
  or GNAME9141(G9141,G9143,G9142);
  and GNAME9142(G9142,G11526,G416);
  and GNAME9143(G9143,G9145,G9144);
  not GNAME9144(G9144,G416);
  dff DFF_9146(CK,G9145,G9141);
  and GNAME9147(G9147,G9145,G9148);
  nand GNAME9148(G9148,G80,G9150);
  buf GNAME9149(G9149,G9145);
  buf GNAME9150(G9150,G9132);
  or GNAME9162(G9162,G9164,G9163);
  and GNAME9163(G9163,G11525,G416);
  and GNAME9164(G9164,G9166,G9165);
  not GNAME9165(G9165,G416);
  dff DFF_9167(CK,G9166,G9162);
  and GNAME9168(G9168,G9166,G9169);
  nand GNAME9169(G9169,G80,G9171);
  buf GNAME9170(G9170,G9166);
  buf GNAME9171(G9171,G9153);
  or GNAME9183(G9183,G9185,G9184);
  and GNAME9184(G9184,G11524,G416);
  and GNAME9185(G9185,G9187,G9186);
  not GNAME9186(G9186,G416);
  dff DFF_9188(CK,G9187,G9183);
  and GNAME9189(G9189,G9187,G9190);
  nand GNAME9190(G9190,G80,G9192);
  buf GNAME9191(G9191,G9187);
  buf GNAME9192(G9192,G9174);
  or GNAME9204(G9204,G9206,G9205);
  and GNAME9205(G9205,G11523,G416);
  and GNAME9206(G9206,G9208,G9207);
  not GNAME9207(G9207,G416);
  dff DFF_9209(CK,G9208,G9204);
  and GNAME9210(G9210,G9208,G9211);
  nand GNAME9211(G9211,G80,G9213);
  buf GNAME9212(G9212,G9208);
  buf GNAME9213(G9213,G9195);
  or GNAME9265(G9265,G9267,G9266);
  and GNAME9266(G9266,G11522,G407);
  and GNAME9267(G9267,G9269,G9268);
  not GNAME9268(G9268,G407);
  dff DFF_9270(CK,G9269,G9265);
  and GNAME9271(G9271,G9269,G9272);
  nand GNAME9272(G9272,G80,G9274);
  buf GNAME9273(G9273,G9269);
  buf GNAME9274(G9274,G9256);
  or GNAME9286(G9286,G9288,G9287);
  and GNAME9287(G9287,G11521,G407);
  and GNAME9288(G9288,G9290,G9289);
  not GNAME9289(G9289,G407);
  dff DFF_9291(CK,G9290,G9286);
  and GNAME9292(G9292,G9290,G9293);
  nand GNAME9293(G9293,G80,G9295);
  buf GNAME9294(G9294,G9290);
  buf GNAME9295(G9295,G9277);
  or GNAME9307(G9307,G9309,G9308);
  and GNAME9308(G9308,G11520,G407);
  and GNAME9309(G9309,G9311,G9310);
  not GNAME9310(G9310,G407);
  dff DFF_9312(CK,G9311,G9307);
  and GNAME9313(G9313,G9311,G9314);
  nand GNAME9314(G9314,G80,G9316);
  buf GNAME9315(G9315,G9311);
  buf GNAME9316(G9316,G9298);
  or GNAME9328(G9328,G9330,G9329);
  and GNAME9329(G9329,G11519,G407);
  and GNAME9330(G9330,G9332,G9331);
  not GNAME9331(G9331,G407);
  dff DFF_9333(CK,G9332,G9328);
  and GNAME9334(G9334,G9332,G9335);
  nand GNAME9335(G9335,G80,G9337);
  buf GNAME9336(G9336,G9332);
  buf GNAME9337(G9337,G9319);
  or GNAME9349(G9349,G9351,G9350);
  and GNAME9350(G9350,G11518,G407);
  and GNAME9351(G9351,G9353,G9352);
  not GNAME9352(G9352,G407);
  dff DFF_9354(CK,G9353,G9349);
  and GNAME9355(G9355,G9353,G9356);
  nand GNAME9356(G9356,G80,G9358);
  buf GNAME9357(G9357,G9353);
  buf GNAME9358(G9358,G9340);
  or GNAME9370(G9370,G9372,G9371);
  and GNAME9371(G9371,G11517,G407);
  and GNAME9372(G9372,G9374,G9373);
  not GNAME9373(G9373,G407);
  dff DFF_9375(CK,G9374,G9370);
  and GNAME9376(G9376,G9374,G9377);
  nand GNAME9377(G9377,G80,G9379);
  buf GNAME9378(G9378,G9374);
  buf GNAME9379(G9379,G9361);
  or GNAME9391(G9391,G9393,G9392);
  and GNAME9392(G9392,G11516,G407);
  and GNAME9393(G9393,G9395,G9394);
  not GNAME9394(G9394,G407);
  dff DFF_9396(CK,G9395,G9391);
  and GNAME9397(G9397,G9395,G9398);
  nand GNAME9398(G9398,G80,G9400);
  buf GNAME9399(G9399,G9395);
  buf GNAME9400(G9400,G9382);
  or GNAME9412(G9412,G9414,G9413);
  and GNAME9413(G9413,G11515,G407);
  and GNAME9414(G9414,G9416,G9415);
  not GNAME9415(G9415,G407);
  dff DFF_9417(CK,G9416,G9412);
  and GNAME9418(G9418,G9416,G9419);
  nand GNAME9419(G9419,G80,G9421);
  buf GNAME9420(G9420,G9416);
  buf GNAME9421(G9421,G9403);
  or GNAME9473(G9473,G9475,G9474);
  and GNAME9474(G9474,G11522,G406);
  and GNAME9475(G9475,G9477,G9476);
  not GNAME9476(G9476,G406);
  dff DFF_9478(CK,G9477,G9473);
  and GNAME9479(G9479,G9477,G9480);
  nand GNAME9480(G9480,G80,G9482);
  buf GNAME9481(G9481,G9477);
  buf GNAME9482(G9482,G9464);
  or GNAME9494(G9494,G9496,G9495);
  and GNAME9495(G9495,G11521,G406);
  and GNAME9496(G9496,G9498,G9497);
  not GNAME9497(G9497,G406);
  dff DFF_9499(CK,G9498,G9494);
  and GNAME9500(G9500,G9498,G9501);
  nand GNAME9501(G9501,G80,G9503);
  buf GNAME9502(G9502,G9498);
  buf GNAME9503(G9503,G9485);
  or GNAME9515(G9515,G9517,G9516);
  and GNAME9516(G9516,G11520,G406);
  and GNAME9517(G9517,G9519,G9518);
  not GNAME9518(G9518,G406);
  dff DFF_9520(CK,G9519,G9515);
  and GNAME9521(G9521,G9519,G9522);
  nand GNAME9522(G9522,G80,G9524);
  buf GNAME9523(G9523,G9519);
  buf GNAME9524(G9524,G9506);
  or GNAME9536(G9536,G9538,G9537);
  and GNAME9537(G9537,G11519,G406);
  and GNAME9538(G9538,G9540,G9539);
  not GNAME9539(G9539,G406);
  dff DFF_9541(CK,G9540,G9536);
  and GNAME9542(G9542,G9540,G9543);
  nand GNAME9543(G9543,G80,G9545);
  buf GNAME9544(G9544,G9540);
  buf GNAME9545(G9545,G9527);
  or GNAME9557(G9557,G9559,G9558);
  and GNAME9558(G9558,G11518,G406);
  and GNAME9559(G9559,G9561,G9560);
  not GNAME9560(G9560,G406);
  dff DFF_9562(CK,G9561,G9557);
  and GNAME9563(G9563,G9561,G9564);
  nand GNAME9564(G9564,G80,G9566);
  buf GNAME9565(G9565,G9561);
  buf GNAME9566(G9566,G9548);
  or GNAME9578(G9578,G9580,G9579);
  and GNAME9579(G9579,G11517,G406);
  and GNAME9580(G9580,G9582,G9581);
  not GNAME9581(G9581,G406);
  dff DFF_9583(CK,G9582,G9578);
  and GNAME9584(G9584,G9582,G9585);
  nand GNAME9585(G9585,G80,G9587);
  buf GNAME9586(G9586,G9582);
  buf GNAME9587(G9587,G9569);
  or GNAME9599(G9599,G9601,G9600);
  and GNAME9600(G9600,G11516,G406);
  and GNAME9601(G9601,G9603,G9602);
  not GNAME9602(G9602,G406);
  dff DFF_9604(CK,G9603,G9599);
  and GNAME9605(G9605,G9603,G9606);
  nand GNAME9606(G9606,G80,G9608);
  buf GNAME9607(G9607,G9603);
  buf GNAME9608(G9608,G9590);
  or GNAME9620(G9620,G9622,G9621);
  and GNAME9621(G9621,G11515,G406);
  and GNAME9622(G9622,G9624,G9623);
  not GNAME9623(G9623,G406);
  dff DFF_9625(CK,G9624,G9620);
  and GNAME9626(G9626,G9624,G9627);
  nand GNAME9627(G9627,G80,G9629);
  buf GNAME9628(G9628,G9624);
  buf GNAME9629(G9629,G9611);
  or GNAME9681(G9681,G9683,G9682);
  and GNAME9682(G9682,G11522,G405);
  and GNAME9683(G9683,G9685,G9684);
  not GNAME9684(G9684,G405);
  dff DFF_9686(CK,G9685,G9681);
  and GNAME9687(G9687,G9685,G9688);
  nand GNAME9688(G9688,G80,G9690);
  buf GNAME9689(G9689,G9685);
  buf GNAME9690(G9690,G9672);
  or GNAME9702(G9702,G9704,G9703);
  and GNAME9703(G9703,G11521,G405);
  and GNAME9704(G9704,G9706,G9705);
  not GNAME9705(G9705,G405);
  dff DFF_9707(CK,G9706,G9702);
  and GNAME9708(G9708,G9706,G9709);
  nand GNAME9709(G9709,G80,G9711);
  buf GNAME9710(G9710,G9706);
  buf GNAME9711(G9711,G9693);
  or GNAME9723(G9723,G9725,G9724);
  and GNAME9724(G9724,G11520,G405);
  and GNAME9725(G9725,G9727,G9726);
  not GNAME9726(G9726,G405);
  dff DFF_9728(CK,G9727,G9723);
  and GNAME9729(G9729,G9727,G9730);
  nand GNAME9730(G9730,G80,G9732);
  buf GNAME9731(G9731,G9727);
  buf GNAME9732(G9732,G9714);
  or GNAME9744(G9744,G9746,G9745);
  and GNAME9745(G9745,G11519,G405);
  and GNAME9746(G9746,G9748,G9747);
  not GNAME9747(G9747,G405);
  dff DFF_9749(CK,G9748,G9744);
  and GNAME9750(G9750,G9748,G9751);
  nand GNAME9751(G9751,G80,G9753);
  buf GNAME9752(G9752,G9748);
  buf GNAME9753(G9753,G9735);
  or GNAME9765(G9765,G9767,G9766);
  and GNAME9766(G9766,G11518,G405);
  and GNAME9767(G9767,G9769,G9768);
  not GNAME9768(G9768,G405);
  dff DFF_9770(CK,G9769,G9765);
  and GNAME9771(G9771,G9769,G9772);
  nand GNAME9772(G9772,G80,G9774);
  buf GNAME9773(G9773,G9769);
  buf GNAME9774(G9774,G9756);
  or GNAME9786(G9786,G9788,G9787);
  and GNAME9787(G9787,G11517,G405);
  and GNAME9788(G9788,G9790,G9789);
  not GNAME9789(G9789,G405);
  dff DFF_9791(CK,G9790,G9786);
  and GNAME9792(G9792,G9790,G9793);
  nand GNAME9793(G9793,G80,G9795);
  buf GNAME9794(G9794,G9790);
  buf GNAME9795(G9795,G9777);
  or GNAME9807(G9807,G9809,G9808);
  and GNAME9808(G9808,G11516,G405);
  and GNAME9809(G9809,G9811,G9810);
  not GNAME9810(G9810,G405);
  dff DFF_9812(CK,G9811,G9807);
  and GNAME9813(G9813,G9811,G9814);
  nand GNAME9814(G9814,G80,G9816);
  buf GNAME9815(G9815,G9811);
  buf GNAME9816(G9816,G9798);
  or GNAME9828(G9828,G9830,G9829);
  and GNAME9829(G9829,G11515,G405);
  and GNAME9830(G9830,G9832,G9831);
  not GNAME9831(G9831,G405);
  dff DFF_9833(CK,G9832,G9828);
  and GNAME9834(G9834,G9832,G9835);
  nand GNAME9835(G9835,G80,G9837);
  buf GNAME9836(G9836,G9832);
  buf GNAME9837(G9837,G9819);
  or GNAME9889(G9889,G9891,G9890);
  and GNAME9890(G9890,G11522,G404);
  and GNAME9891(G9891,G9893,G9892);
  not GNAME9892(G9892,G404);
  dff DFF_9894(CK,G9893,G9889);
  and GNAME9895(G9895,G9893,G9896);
  nand GNAME9896(G9896,G80,G9898);
  buf GNAME9897(G9897,G9893);
  buf GNAME9898(G9898,G9880);
  or GNAME9910(G9910,G9912,G9911);
  and GNAME9911(G9911,G11521,G404);
  and GNAME9912(G9912,G9914,G9913);
  not GNAME9913(G9913,G404);
  dff DFF_9915(CK,G9914,G9910);
  and GNAME9916(G9916,G9914,G9917);
  nand GNAME9917(G9917,G80,G9919);
  buf GNAME9918(G9918,G9914);
  buf GNAME9919(G9919,G9901);
  or GNAME9931(G9931,G9933,G9932);
  and GNAME9932(G9932,G11520,G404);
  and GNAME9933(G9933,G9935,G9934);
  not GNAME9934(G9934,G404);
  dff DFF_9936(CK,G9935,G9931);
  and GNAME9937(G9937,G9935,G9938);
  nand GNAME9938(G9938,G80,G9940);
  buf GNAME9939(G9939,G9935);
  buf GNAME9940(G9940,G9922);
  or GNAME9952(G9952,G9954,G9953);
  and GNAME9953(G9953,G11519,G404);
  and GNAME9954(G9954,G9956,G9955);
  not GNAME9955(G9955,G404);
  dff DFF_9957(CK,G9956,G9952);
  and GNAME9958(G9958,G9956,G9959);
  nand GNAME9959(G9959,G80,G9961);
  buf GNAME9960(G9960,G9956);
  buf GNAME9961(G9961,G9943);
  or GNAME9973(G9973,G9975,G9974);
  and GNAME9974(G9974,G11518,G404);
  and GNAME9975(G9975,G9977,G9976);
  not GNAME9976(G9976,G404);
  dff DFF_9978(CK,G9977,G9973);
  and GNAME9979(G9979,G9977,G9980);
  nand GNAME9980(G9980,G80,G9982);
  buf GNAME9981(G9981,G9977);
  buf GNAME9982(G9982,G9964);
  or GNAME9994(G9994,G9996,G9995);
  and GNAME9995(G9995,G11517,G404);
  and GNAME9996(G9996,G9998,G9997);
  not GNAME9997(G9997,G404);
  dff DFF_9999(CK,G9998,G9994);
  and GNAME10000(G10000,G9998,G10001);
  nand GNAME10001(G10001,G80,G10003);
  buf GNAME10002(G10002,G9998);
  buf GNAME10003(G10003,G9985);
  or GNAME10015(G10015,G10017,G10016);
  and GNAME10016(G10016,G11516,G404);
  and GNAME10017(G10017,G10019,G10018);
  not GNAME10018(G10018,G404);
  dff DFF_10020(CK,G10019,G10015);
  and GNAME10021(G10021,G10019,G10022);
  nand GNAME10022(G10022,G80,G10024);
  buf GNAME10023(G10023,G10019);
  buf GNAME10024(G10024,G10006);
  or GNAME10036(G10036,G10038,G10037);
  and GNAME10037(G10037,G11515,G404);
  and GNAME10038(G10038,G10040,G10039);
  not GNAME10039(G10039,G404);
  dff DFF_10041(CK,G10040,G10036);
  and GNAME10042(G10042,G10040,G10043);
  nand GNAME10043(G10043,G80,G10045);
  buf GNAME10044(G10044,G10040);
  buf GNAME10045(G10045,G10027);
  or GNAME10097(G10097,G10099,G10098);
  and GNAME10098(G10098,G11522,G415);
  and GNAME10099(G10099,G10101,G10100);
  not GNAME10100(G10100,G415);
  dff DFF_10102(CK,G10101,G10097);
  and GNAME10103(G10103,G10101,G10104);
  nand GNAME10104(G10104,G80,G10106);
  buf GNAME10105(G10105,G10101);
  buf GNAME10106(G10106,G10088);
  or GNAME10118(G10118,G10120,G10119);
  and GNAME10119(G10119,G11521,G415);
  and GNAME10120(G10120,G10122,G10121);
  not GNAME10121(G10121,G415);
  dff DFF_10123(CK,G10122,G10118);
  and GNAME10124(G10124,G10122,G10125);
  nand GNAME10125(G10125,G80,G10127);
  buf GNAME10126(G10126,G10122);
  buf GNAME10127(G10127,G10109);
  or GNAME10139(G10139,G10141,G10140);
  and GNAME10140(G10140,G11520,G415);
  and GNAME10141(G10141,G10143,G10142);
  not GNAME10142(G10142,G415);
  dff DFF_10144(CK,G10143,G10139);
  and GNAME10145(G10145,G10143,G10146);
  nand GNAME10146(G10146,G80,G10148);
  buf GNAME10147(G10147,G10143);
  buf GNAME10148(G10148,G10130);
  or GNAME10160(G10160,G10162,G10161);
  and GNAME10161(G10161,G11519,G415);
  and GNAME10162(G10162,G10164,G10163);
  not GNAME10163(G10163,G415);
  dff DFF_10165(CK,G10164,G10160);
  and GNAME10166(G10166,G10164,G10167);
  nand GNAME10167(G10167,G80,G10169);
  buf GNAME10168(G10168,G10164);
  buf GNAME10169(G10169,G10151);
  or GNAME10181(G10181,G10183,G10182);
  and GNAME10182(G10182,G11518,G415);
  and GNAME10183(G10183,G10185,G10184);
  not GNAME10184(G10184,G415);
  dff DFF_10186(CK,G10185,G10181);
  and GNAME10187(G10187,G10185,G10188);
  nand GNAME10188(G10188,G80,G10190);
  buf GNAME10189(G10189,G10185);
  buf GNAME10190(G10190,G10172);
  or GNAME10202(G10202,G10204,G10203);
  and GNAME10203(G10203,G11517,G415);
  and GNAME10204(G10204,G10206,G10205);
  not GNAME10205(G10205,G415);
  dff DFF_10207(CK,G10206,G10202);
  and GNAME10208(G10208,G10206,G10209);
  nand GNAME10209(G10209,G80,G10211);
  buf GNAME10210(G10210,G10206);
  buf GNAME10211(G10211,G10193);
  or GNAME10223(G10223,G10225,G10224);
  and GNAME10224(G10224,G11516,G415);
  and GNAME10225(G10225,G10227,G10226);
  not GNAME10226(G10226,G415);
  dff DFF_10228(CK,G10227,G10223);
  and GNAME10229(G10229,G10227,G10230);
  nand GNAME10230(G10230,G80,G10232);
  buf GNAME10231(G10231,G10227);
  buf GNAME10232(G10232,G10214);
  or GNAME10244(G10244,G10246,G10245);
  and GNAME10245(G10245,G11515,G415);
  and GNAME10246(G10246,G10248,G10247);
  not GNAME10247(G10247,G415);
  dff DFF_10249(CK,G10248,G10244);
  and GNAME10250(G10250,G10248,G10251);
  nand GNAME10251(G10251,G80,G10253);
  buf GNAME10252(G10252,G10248);
  buf GNAME10253(G10253,G10235);
  or GNAME10305(G10305,G10307,G10306);
  and GNAME10306(G10306,G11522,G414);
  and GNAME10307(G10307,G10309,G10308);
  not GNAME10308(G10308,G414);
  dff DFF_10310(CK,G10309,G10305);
  and GNAME10311(G10311,G10309,G10312);
  nand GNAME10312(G10312,G80,G10314);
  buf GNAME10313(G10313,G10309);
  buf GNAME10314(G10314,G10296);
  or GNAME10326(G10326,G10328,G10327);
  and GNAME10327(G10327,G11521,G414);
  and GNAME10328(G10328,G10330,G10329);
  not GNAME10329(G10329,G414);
  dff DFF_10331(CK,G10330,G10326);
  and GNAME10332(G10332,G10330,G10333);
  nand GNAME10333(G10333,G80,G10335);
  buf GNAME10334(G10334,G10330);
  buf GNAME10335(G10335,G10317);
  or GNAME10347(G10347,G10349,G10348);
  and GNAME10348(G10348,G11520,G414);
  and GNAME10349(G10349,G10351,G10350);
  not GNAME10350(G10350,G414);
  dff DFF_10352(CK,G10351,G10347);
  and GNAME10353(G10353,G10351,G10354);
  nand GNAME10354(G10354,G80,G10356);
  buf GNAME10355(G10355,G10351);
  buf GNAME10356(G10356,G10338);
  or GNAME10368(G10368,G10370,G10369);
  and GNAME10369(G10369,G11519,G414);
  and GNAME10370(G10370,G10372,G10371);
  not GNAME10371(G10371,G414);
  dff DFF_10373(CK,G10372,G10368);
  and GNAME10374(G10374,G10372,G10375);
  nand GNAME10375(G10375,G80,G10377);
  buf GNAME10376(G10376,G10372);
  buf GNAME10377(G10377,G10359);
  or GNAME10389(G10389,G10391,G10390);
  and GNAME10390(G10390,G11518,G414);
  and GNAME10391(G10391,G10393,G10392);
  not GNAME10392(G10392,G414);
  dff DFF_10394(CK,G10393,G10389);
  and GNAME10395(G10395,G10393,G10396);
  nand GNAME10396(G10396,G80,G10398);
  buf GNAME10397(G10397,G10393);
  buf GNAME10398(G10398,G10380);
  or GNAME10410(G10410,G10412,G10411);
  and GNAME10411(G10411,G11517,G414);
  and GNAME10412(G10412,G10414,G10413);
  not GNAME10413(G10413,G414);
  dff DFF_10415(CK,G10414,G10410);
  and GNAME10416(G10416,G10414,G10417);
  nand GNAME10417(G10417,G80,G10419);
  buf GNAME10418(G10418,G10414);
  buf GNAME10419(G10419,G10401);
  or GNAME10431(G10431,G10433,G10432);
  and GNAME10432(G10432,G11516,G414);
  and GNAME10433(G10433,G10435,G10434);
  not GNAME10434(G10434,G414);
  dff DFF_10436(CK,G10435,G10431);
  and GNAME10437(G10437,G10435,G10438);
  nand GNAME10438(G10438,G80,G10440);
  buf GNAME10439(G10439,G10435);
  buf GNAME10440(G10440,G10422);
  or GNAME10452(G10452,G10454,G10453);
  and GNAME10453(G10453,G11515,G414);
  and GNAME10454(G10454,G10456,G10455);
  not GNAME10455(G10455,G414);
  dff DFF_10457(CK,G10456,G10452);
  and GNAME10458(G10458,G10456,G10459);
  nand GNAME10459(G10459,G80,G10461);
  buf GNAME10460(G10460,G10456);
  buf GNAME10461(G10461,G10443);
  or GNAME10513(G10513,G10515,G10514);
  and GNAME10514(G10514,G11522,G413);
  and GNAME10515(G10515,G10517,G10516);
  not GNAME10516(G10516,G413);
  dff DFF_10518(CK,G10517,G10513);
  and GNAME10519(G10519,G10517,G10520);
  nand GNAME10520(G10520,G80,G10522);
  buf GNAME10521(G10521,G10517);
  buf GNAME10522(G10522,G10504);
  or GNAME10534(G10534,G10536,G10535);
  and GNAME10535(G10535,G11521,G413);
  and GNAME10536(G10536,G10538,G10537);
  not GNAME10537(G10537,G413);
  dff DFF_10539(CK,G10538,G10534);
  and GNAME10540(G10540,G10538,G10541);
  nand GNAME10541(G10541,G80,G10543);
  buf GNAME10542(G10542,G10538);
  buf GNAME10543(G10543,G10525);
  or GNAME10555(G10555,G10557,G10556);
  and GNAME10556(G10556,G11520,G413);
  and GNAME10557(G10557,G10559,G10558);
  not GNAME10558(G10558,G413);
  dff DFF_10560(CK,G10559,G10555);
  and GNAME10561(G10561,G10559,G10562);
  nand GNAME10562(G10562,G80,G10564);
  buf GNAME10563(G10563,G10559);
  buf GNAME10564(G10564,G10546);
  or GNAME10576(G10576,G10578,G10577);
  and GNAME10577(G10577,G11519,G413);
  and GNAME10578(G10578,G10580,G10579);
  not GNAME10579(G10579,G413);
  dff DFF_10581(CK,G10580,G10576);
  and GNAME10582(G10582,G10580,G10583);
  nand GNAME10583(G10583,G80,G10585);
  buf GNAME10584(G10584,G10580);
  buf GNAME10585(G10585,G10567);
  or GNAME10597(G10597,G10599,G10598);
  and GNAME10598(G10598,G11518,G413);
  and GNAME10599(G10599,G10601,G10600);
  not GNAME10600(G10600,G413);
  dff DFF_10602(CK,G10601,G10597);
  and GNAME10603(G10603,G10601,G10604);
  nand GNAME10604(G10604,G80,G10606);
  buf GNAME10605(G10605,G10601);
  buf GNAME10606(G10606,G10588);
  or GNAME10618(G10618,G10620,G10619);
  and GNAME10619(G10619,G11517,G413);
  and GNAME10620(G10620,G10622,G10621);
  not GNAME10621(G10621,G413);
  dff DFF_10623(CK,G10622,G10618);
  and GNAME10624(G10624,G10622,G10625);
  nand GNAME10625(G10625,G80,G10627);
  buf GNAME10626(G10626,G10622);
  buf GNAME10627(G10627,G10609);
  or GNAME10639(G10639,G10641,G10640);
  and GNAME10640(G10640,G11516,G413);
  and GNAME10641(G10641,G10643,G10642);
  not GNAME10642(G10642,G413);
  dff DFF_10644(CK,G10643,G10639);
  and GNAME10645(G10645,G10643,G10646);
  nand GNAME10646(G10646,G80,G10648);
  buf GNAME10647(G10647,G10643);
  buf GNAME10648(G10648,G10630);
  or GNAME10660(G10660,G10662,G10661);
  and GNAME10661(G10661,G11515,G413);
  and GNAME10662(G10662,G10664,G10663);
  not GNAME10663(G10663,G413);
  dff DFF_10665(CK,G10664,G10660);
  and GNAME10666(G10666,G10664,G10667);
  nand GNAME10667(G10667,G80,G10669);
  buf GNAME10668(G10668,G10664);
  buf GNAME10669(G10669,G10651);
  or GNAME10721(G10721,G10723,G10722);
  and GNAME10722(G10722,G11522,G412);
  and GNAME10723(G10723,G10725,G10724);
  not GNAME10724(G10724,G412);
  dff DFF_10726(CK,G10725,G10721);
  and GNAME10727(G10727,G10725,G10728);
  nand GNAME10728(G10728,G80,G10730);
  buf GNAME10729(G10729,G10725);
  buf GNAME10730(G10730,G10712);
  or GNAME10742(G10742,G10744,G10743);
  and GNAME10743(G10743,G11521,G412);
  and GNAME10744(G10744,G10746,G10745);
  not GNAME10745(G10745,G412);
  dff DFF_10747(CK,G10746,G10742);
  and GNAME10748(G10748,G10746,G10749);
  nand GNAME10749(G10749,G80,G10751);
  buf GNAME10750(G10750,G10746);
  buf GNAME10751(G10751,G10733);
  or GNAME10763(G10763,G10765,G10764);
  and GNAME10764(G10764,G11520,G412);
  and GNAME10765(G10765,G10767,G10766);
  not GNAME10766(G10766,G412);
  dff DFF_10768(CK,G10767,G10763);
  and GNAME10769(G10769,G10767,G10770);
  nand GNAME10770(G10770,G80,G10772);
  buf GNAME10771(G10771,G10767);
  buf GNAME10772(G10772,G10754);
  or GNAME10784(G10784,G10786,G10785);
  and GNAME10785(G10785,G11519,G412);
  and GNAME10786(G10786,G10788,G10787);
  not GNAME10787(G10787,G412);
  dff DFF_10789(CK,G10788,G10784);
  and GNAME10790(G10790,G10788,G10791);
  nand GNAME10791(G10791,G80,G10793);
  buf GNAME10792(G10792,G10788);
  buf GNAME10793(G10793,G10775);
  or GNAME10805(G10805,G10807,G10806);
  and GNAME10806(G10806,G11518,G412);
  and GNAME10807(G10807,G10809,G10808);
  not GNAME10808(G10808,G412);
  dff DFF_10810(CK,G10809,G10805);
  and GNAME10811(G10811,G10809,G10812);
  nand GNAME10812(G10812,G80,G10814);
  buf GNAME10813(G10813,G10809);
  buf GNAME10814(G10814,G10796);
  or GNAME10826(G10826,G10828,G10827);
  and GNAME10827(G10827,G11517,G412);
  and GNAME10828(G10828,G10830,G10829);
  not GNAME10829(G10829,G412);
  dff DFF_10831(CK,G10830,G10826);
  and GNAME10832(G10832,G10830,G10833);
  nand GNAME10833(G10833,G80,G10835);
  buf GNAME10834(G10834,G10830);
  buf GNAME10835(G10835,G10817);
  or GNAME10847(G10847,G10849,G10848);
  and GNAME10848(G10848,G11516,G412);
  and GNAME10849(G10849,G10851,G10850);
  not GNAME10850(G10850,G412);
  dff DFF_10852(CK,G10851,G10847);
  and GNAME10853(G10853,G10851,G10854);
  nand GNAME10854(G10854,G80,G10856);
  buf GNAME10855(G10855,G10851);
  buf GNAME10856(G10856,G10838);
  or GNAME10868(G10868,G10870,G10869);
  and GNAME10869(G10869,G11515,G412);
  and GNAME10870(G10870,G10872,G10871);
  not GNAME10871(G10871,G412);
  dff DFF_10873(CK,G10872,G10868);
  and GNAME10874(G10874,G10872,G10875);
  nand GNAME10875(G10875,G80,G10877);
  buf GNAME10876(G10876,G10872);
  buf GNAME10877(G10877,G10859);
  nor GNAME11072(G11072,G11495,G454,G11298);
  nor GNAME11073(G11073,G11494,G11072,G11281);
  nor GNAME11074(G11074,G11187,G11186,G11497);
  not GNAME11075(G11075,G11078);
  not GNAME11076(G11076,G11188);
  not GNAME11077(G11077,G11130);
  and GNAME11078(G11078,G11246,G11290,G11077,G11076);
  not GNAME11079(G11079,G11082);
  not GNAME11080(G11080,G11189);
  not GNAME11081(G11081,G11135);
  and GNAME11082(G11082,G11249,G11291,G11081,G11080);
  not GNAME11083(G11083,G11086);
  not GNAME11084(G11084,G11190);
  not GNAME11085(G11085,G11140);
  and GNAME11086(G11086,G11252,G11292,G11085,G11084);
  not GNAME11087(G11087,G11090);
  not GNAME11088(G11088,G11191);
  not GNAME11089(G11089,G11145);
  and GNAME11090(G11090,G11255,G11293,G11089,G11088);
  not GNAME11091(G11091,G11094);
  not GNAME11092(G11092,G11192);
  not GNAME11093(G11093,G11150);
  and GNAME11094(G11094,G11258,G11294,G11093,G11092);
  not GNAME11095(G11095,G11098);
  not GNAME11096(G11096,G11193);
  not GNAME11097(G11097,G11155);
  and GNAME11098(G11098,G11261,G11295,G11097,G11096);
  not GNAME11099(G11099,G11102);
  not GNAME11100(G11100,G11194);
  not GNAME11101(G11101,G11160);
  and GNAME11102(G11102,G11264,G11296,G11101,G11100);
  not GNAME11103(G11103,G11106);
  not GNAME11104(G11104,G11195);
  not GNAME11105(G11105,G11165);
  and GNAME11106(G11106,G11267,G11297,G11105,G11104);
  not GNAME11107(G11107,G11110);
  not GNAME11108(G11108,G11122);
  not GNAME11109(G11109,G11184);
  and GNAME11110(G11110,G11300,G11074,G11109,G11108);
  not GNAME11111(G11111,G11114);
  not GNAME11112(G11112,G11107);
  not GNAME11113(G11113,G11272);
  and GNAME11114(G11114,G11073,G11280,G11113,G11112);
  not GNAME11115(G11115,G11117);
  not GNAME11116(G11116,G11170);
  or GNAME11117(G11117,G445,G11116);
  not GNAME11118(G11118,G11121);
  not GNAME11119(G11119,G448);
  not GNAME11120(G11120,G11276);
  or GNAME11121(G11121,G451,G11120,G11119);
  not GNAME11122(G11122,G11125);
  not GNAME11123(G11123,G444);
  not GNAME11124(G11124,G11115);
  or GNAME11125(G11125,G447,G11124,G11123);
  not GNAME11126(G11126,G11129);
  not GNAME11127(G11127,G443);
  not GNAME11128(G11128,G11173);
  or GNAME11129(G11129,G446,G11128,G11127);
  not GNAME11130(G11130,G11134);
  not GNAME11131(G11131,G34579);
  not GNAME11132(G11132,G11272);
  or GNAME11133(G11133,G11132,G11131);
  and GNAME11134(G11134,G11198,G11133);
  not GNAME11135(G11135,G11139);
  not GNAME11136(G11136,G34566);
  not GNAME11137(G11137,G11272);
  or GNAME11138(G11138,G11137,G11136);
  and GNAME11139(G11139,G11201,G11138);
  not GNAME11140(G11140,G11144);
  not GNAME11141(G11141,G34553);
  not GNAME11142(G11142,G11272);
  or GNAME11143(G11143,G11142,G11141);
  and GNAME11144(G11144,G11204,G11143);
  not GNAME11145(G11145,G11149);
  not GNAME11146(G11146,G34540);
  not GNAME11147(G11147,G11272);
  or GNAME11148(G11148,G11147,G11146);
  and GNAME11149(G11149,G11207,G11148);
  not GNAME11150(G11150,G11154);
  not GNAME11151(G11151,G34527);
  not GNAME11152(G11152,G11272);
  or GNAME11153(G11153,G11152,G11151);
  and GNAME11154(G11154,G11210,G11153);
  not GNAME11155(G11155,G11159);
  not GNAME11156(G11156,G34514);
  not GNAME11157(G11157,G11272);
  or GNAME11158(G11158,G11157,G11156);
  and GNAME11159(G11159,G11213,G11158);
  not GNAME11160(G11160,G11164);
  not GNAME11161(G11161,G34501);
  not GNAME11162(G11162,G11272);
  or GNAME11163(G11163,G11162,G11161);
  and GNAME11164(G11164,G11216,G11163);
  not GNAME11165(G11165,G11169);
  not GNAME11166(G11166,G34488);
  not GNAME11167(G11167,G11272);
  or GNAME11168(G11168,G11167,G11166);
  and GNAME11169(G11169,G11219,G11168);
  not GNAME11170(G11170,G11172);
  not GNAME11171(G11171,G11276);
  or GNAME11172(G11172,G451,G448,G11171);
  not GNAME11173(G11173,G11175);
  not GNAME11174(G11174,G11115);
  or GNAME11175(G11175,G447,G444,G11174);
  and GNAME11176(G11176,G57238,G11187);
  and GNAME11177(G11177,G57225,G11187);
  and GNAME11178(G11178,G57212,G11187);
  and GNAME11179(G11179,G57199,G11187);
  and GNAME11180(G11180,G57186,G11187);
  and GNAME11181(G11181,G57173,G11187);
  and GNAME11182(G11182,G57160,G11187);
  and GNAME11183(G11183,G57147,G11187);
  and GNAME11184(G11184,G445,G11170);
  and GNAME11185(G11185,G446,G11173);
  and GNAME11186(G11186,G11115,G447);
  and GNAME11187(G11187,G11276,G451);
  nand GNAME11188(G11188,G11222,G11282,G11303);
  nand GNAME11189(G11189,G11225,G11289,G11306);
  nand GNAME11190(G11190,G11228,G11283,G11309);
  nand GNAME11191(G11191,G11231,G11284,G11312);
  nand GNAME11192(G11192,G11234,G11285,G11315);
  nand GNAME11193(G11193,G11237,G11286,G11318);
  nand GNAME11194(G11194,G11240,G11287,G11321);
  nand GNAME11195(G11195,G11243,G11288,G11324);
  and GNAME11196(G11196,G34319,G11072);
  and GNAME11197(G11197,G34215,G11281);
  nor GNAME11198(G11198,G11197,G11196);
  and GNAME11199(G11199,G34306,G11072);
  and GNAME11200(G11200,G34202,G11281);
  nor GNAME11201(G11201,G11200,G11199);
  and GNAME11202(G11202,G34293,G11072);
  and GNAME11203(G11203,G34189,G11281);
  nor GNAME11204(G11204,G11203,G11202);
  and GNAME11205(G11205,G34280,G11072);
  and GNAME11206(G11206,G34176,G11281);
  nor GNAME11207(G11207,G11206,G11205);
  and GNAME11208(G11208,G34267,G11072);
  and GNAME11209(G11209,G34163,G11281);
  nor GNAME11210(G11210,G11209,G11208);
  and GNAME11211(G11211,G34254,G11072);
  and GNAME11212(G11212,G34150,G11281);
  nor GNAME11213(G11213,G11212,G11211);
  and GNAME11214(G11214,G34241,G11072);
  and GNAME11215(G11215,G34137,G11281);
  nor GNAME11216(G11216,G11215,G11214);
  and GNAME11217(G11217,G34228,G11072);
  and GNAME11218(G11218,G34124,G11281);
  nor GNAME11219(G11219,G11218,G11217);
  and GNAME11220(G11220,G57446,G11184);
  and GNAME11221(G11221,G80365,G11122);
  nor GNAME11222(G11222,G11221,G11220);
  and GNAME11223(G11223,G57433,G11184);
  and GNAME11224(G11224,G80352,G11122);
  nor GNAME11225(G11225,G11224,G11223);
  and GNAME11226(G11226,G57420,G11184);
  and GNAME11227(G11227,G80339,G11122);
  nor GNAME11228(G11228,G11227,G11226);
  and GNAME11229(G11229,G57407,G11184);
  and GNAME11230(G11230,G80326,G11122);
  nor GNAME11231(G11231,G11230,G11229);
  and GNAME11232(G11232,G57394,G11184);
  and GNAME11233(G11233,G80313,G11122);
  nor GNAME11234(G11234,G11233,G11232);
  and GNAME11235(G11235,G57381,G11184);
  and GNAME11236(G11236,G80300,G11122);
  nor GNAME11237(G11237,G11236,G11235);
  and GNAME11238(G11238,G57368,G11184);
  and GNAME11239(G11239,G80287,G11122);
  nor GNAME11240(G11240,G11239,G11238);
  and GNAME11241(G11241,G57355,G11184);
  and GNAME11242(G11242,G80274,G11122);
  nor GNAME11243(G11243,G11242,G11241);
  and GNAME11244(G11244,G80573,G11498);
  and GNAME11245(G11245,G80469,G11185);
  nor GNAME11246(G11246,G11245,G11244);
  and GNAME11247(G11247,G80560,G11498);
  and GNAME11248(G11248,G80456,G11185);
  nor GNAME11249(G11249,G11248,G11247);
  and GNAME11250(G11250,G80547,G11498);
  and GNAME11251(G11251,G80443,G11185);
  nor GNAME11252(G11252,G11251,G11250);
  and GNAME11253(G11253,G80534,G11498);
  and GNAME11254(G11254,G80430,G11185);
  nor GNAME11255(G11255,G11254,G11253);
  and GNAME11256(G11256,G80521,G11498);
  and GNAME11257(G11257,G80417,G11185);
  nor GNAME11258(G11258,G11257,G11256);
  and GNAME11259(G11259,G80508,G11498);
  and GNAME11260(G11260,G80404,G11185);
  nor GNAME11261(G11261,G11260,G11259);
  and GNAME11262(G11262,G80495,G11498);
  and GNAME11263(G11263,G80391,G11185);
  nor GNAME11264(G11264,G11263,G11262);
  and GNAME11265(G11265,G80482,G11498);
  and GNAME11266(G11266,G80378,G11185);
  nor GNAME11267(G11267,G11266,G11265);
  not GNAME11268(G11268,G11271);
  not GNAME11269(G11269,G11173);
  not GNAME11270(G11270,G453);
  or GNAME11271(G11271,G443,G446,G11270,G11269);
  not GNAME11272(G11272,G11275);
  not GNAME11273(G11273,G449);
  not GNAME11274(G11274,G11300);
  or GNAME11275(G11275,G452,G454,G11274,G11273);
  not GNAME11276(G11276,G11279);
  not GNAME11277(G11277,G11298);
  not GNAME11278(G11278,G11299);
  or GNAME11279(G11279,G11496,G449,G11278,G11277);
  nor GNAME11280(G11280,G11498,G11185);
  nor GNAME11281(G11281,G11299,G11495);
  nand GNAME11282(G11282,G34098,G11496);
  nand GNAME11283(G11283,G34085,G11496);
  nand GNAME11284(G11284,G34072,G11496);
  nand GNAME11285(G11285,G34059,G11496);
  nand GNAME11286(G11286,G34046,G11496);
  nand GNAME11287(G11287,G34033,G11496);
  nand GNAME11288(G11288,G34020,G11495);
  nand GNAME11289(G11289,G11495,G34111);
  nand GNAME11290(G11290,G80833,G11494);
  nand GNAME11291(G11291,G80820,G11494);
  nand GNAME11292(G11292,G80807,G11494);
  nand GNAME11293(G11293,G80794,G11494);
  nand GNAME11294(G11294,G80781,G11494);
  nand GNAME11295(G11295,G80768,G11494);
  nand GNAME11296(G11296,G80755,G11494);
  nand GNAME11297(G11297,G80742,G11494);
  not GNAME11298(G11298,G452);
  not GNAME11299(G11299,G454);
  not GNAME11300(G11300,G11495);
  and GNAME11301(G11301,G57550,G11497);
  and GNAME11302(G11302,G57342,G11186);
  nor GNAME11303(G11303,G11176,G11302,G11301);
  and GNAME11304(G11304,G57537,G11497);
  and GNAME11305(G11305,G57329,G11186);
  nor GNAME11306(G11306,G11177,G11305,G11304);
  and GNAME11307(G11307,G57524,G11497);
  and GNAME11308(G11308,G57316,G11186);
  nor GNAME11309(G11309,G11178,G11308,G11307);
  and GNAME11310(G11310,G57511,G11497);
  and GNAME11311(G11311,G57303,G11186);
  nor GNAME11312(G11312,G11179,G11311,G11310);
  and GNAME11313(G11313,G57498,G11497);
  and GNAME11314(G11314,G57290,G11186);
  nor GNAME11315(G11315,G11180,G11314,G11313);
  and GNAME11316(G11316,G57485,G11497);
  and GNAME11317(G11317,G57277,G11186);
  nor GNAME11318(G11318,G11181,G11317,G11316);
  and GNAME11319(G11319,G57472,G11497);
  and GNAME11320(G11320,G57264,G11186);
  nor GNAME11321(G11321,G11182,G11320,G11319);
  and GNAME11322(G11322,G57459,G11497);
  and GNAME11323(G11323,G57251,G11186);
  nor GNAME11324(G11324,G11183,G11323,G11322);
  or GNAME11336(G11336,G11338,G11337);
  and GNAME11337(G11337,G11103,G11111);
  and GNAME11338(G11338,G11340,G11339);
  not GNAME11339(G11339,G11111);
  dff DFF_11341(CK,G11340,G11336);
  and GNAME11342(G11342,G11340,G11343);
  nand GNAME11343(G11343,G80,G11345);
  buf GNAME11344(G11344,G11340);
  buf GNAME11345(G11345,G11327);
  or GNAME11357(G11357,G11359,G11358);
  and GNAME11358(G11358,G11099,G11111);
  and GNAME11359(G11359,G11361,G11360);
  not GNAME11360(G11360,G11111);
  dff DFF_11362(CK,G11361,G11357);
  and GNAME11363(G11363,G11361,G11364);
  nand GNAME11364(G11364,G80,G11366);
  buf GNAME11365(G11365,G11361);
  buf GNAME11366(G11366,G11348);
  or GNAME11378(G11378,G11380,G11379);
  and GNAME11379(G11379,G11095,G11111);
  and GNAME11380(G11380,G11382,G11381);
  not GNAME11381(G11381,G11111);
  dff DFF_11383(CK,G11382,G11378);
  and GNAME11384(G11384,G11382,G11385);
  nand GNAME11385(G11385,G80,G11387);
  buf GNAME11386(G11386,G11382);
  buf GNAME11387(G11387,G11369);
  or GNAME11399(G11399,G11401,G11400);
  and GNAME11400(G11400,G11091,G11111);
  and GNAME11401(G11401,G11403,G11402);
  not GNAME11402(G11402,G11111);
  dff DFF_11404(CK,G11403,G11399);
  and GNAME11405(G11405,G11403,G11406);
  nand GNAME11406(G11406,G80,G11408);
  buf GNAME11407(G11407,G11403);
  buf GNAME11408(G11408,G11390);
  or GNAME11420(G11420,G11422,G11421);
  and GNAME11421(G11421,G11087,G11111);
  and GNAME11422(G11422,G11424,G11423);
  not GNAME11423(G11423,G11111);
  dff DFF_11425(CK,G11424,G11420);
  and GNAME11426(G11426,G11424,G11427);
  nand GNAME11427(G11427,G80,G11429);
  buf GNAME11428(G11428,G11424);
  buf GNAME11429(G11429,G11411);
  or GNAME11441(G11441,G11443,G11442);
  and GNAME11442(G11442,G11083,G11111);
  and GNAME11443(G11443,G11445,G11444);
  not GNAME11444(G11444,G11111);
  dff DFF_11446(CK,G11445,G11441);
  and GNAME11447(G11447,G11445,G11448);
  nand GNAME11448(G11448,G80,G11450);
  buf GNAME11449(G11449,G11445);
  buf GNAME11450(G11450,G11432);
  or GNAME11462(G11462,G11464,G11463);
  and GNAME11463(G11463,G11079,G11111);
  and GNAME11464(G11464,G11466,G11465);
  not GNAME11465(G11465,G11111);
  dff DFF_11467(CK,G11466,G11462);
  and GNAME11468(G11468,G11466,G11469);
  nand GNAME11469(G11469,G80,G11471);
  buf GNAME11470(G11470,G11466);
  buf GNAME11471(G11471,G11453);
  or GNAME11484(G11484,G11486,G11485);
  and GNAME11485(G11485,G11075,G11111);
  and GNAME11486(G11486,G11488,G11487);
  not GNAME11487(G11487,G11111);
  dff DFF_11489(CK,G11488,G11484);
  and GNAME11490(G11490,G11488,G11491);
  nand GNAME11491(G11491,G80,G11493);
  buf GNAME11492(G11492,G11488);
  buf GNAME11493(G11493,G11475);
  buf GNAME11494(G11494,G11268);
  buf GNAME11495(G11495,G450);
  buf GNAME11496(G11496,G450);
  buf GNAME11497(G11497,G11118);
  buf GNAME11498(G11498,G11126);
  buf GNAME11499(G11499,G1304);
  buf GNAME11500(G11500,G1451);
  buf GNAME11501(G11501,G1430);
  buf GNAME11502(G11502,G1409);
  buf GNAME11503(G11503,G1388);
  buf GNAME11504(G11504,G1367);
  buf GNAME11505(G11505,G1346);
  buf GNAME11506(G11506,G1325);
  buf GNAME11507(G11507,G1304);
  buf GNAME11508(G11508,G1451);
  buf GNAME11509(G11509,G1430);
  buf GNAME11510(G11510,G1409);
  buf GNAME11511(G11511,G1388);
  buf GNAME11512(G11512,G1367);
  buf GNAME11513(G11513,G1346);
  buf GNAME11514(G11514,G1325);
  buf GNAME11515(G11515,G11499);
  buf GNAME11516(G11516,G11500);
  buf GNAME11517(G11517,G11501);
  buf GNAME11518(G11518,G11502);
  buf GNAME11519(G11519,G11503);
  buf GNAME11520(G11520,G11504);
  buf GNAME11521(G11521,G11505);
  buf GNAME11522(G11522,G11506);
  buf GNAME11523(G11523,G11499);
  buf GNAME11524(G11524,G11500);
  buf GNAME11525(G11525,G11501);
  buf GNAME11526(G11526,G11502);
  buf GNAME11527(G11527,G11503);
  buf GNAME11528(G11528,G11504);
  buf GNAME11529(G11529,G11505);
  buf GNAME11530(G11530,G11506);
  buf GNAME11531(G11531,G11507);
  buf GNAME11532(G11532,G11508);
  buf GNAME11533(G11533,G11509);
  buf GNAME11534(G11534,G11510);
  buf GNAME11535(G11535,G11511);
  buf GNAME11536(G11536,G11512);
  buf GNAME11537(G11537,G11513);
  buf GNAME11538(G11538,G11514);
  buf GNAME11539(G11539,G11507);
  buf GNAME11540(G11540,G11508);
  buf GNAME11541(G11541,G11509);
  buf GNAME11542(G11542,G11510);
  buf GNAME11543(G11543,G11511);
  buf GNAME11544(G11544,G11512);
  buf GNAME11545(G11545,G11513);
  buf GNAME11546(G11546,G11514);
  xor GNAME17226(G17226,G17227,G29638);
  xor GNAME17227(G17227,G28927,G28924);
  and GNAME17228(G17228,G28927,G29638);
  and GNAME17229(G17229,G28924,G29638);
  and GNAME17230(G17230,G28927,G28924);
  or GNAME17231(G17231,G17230,G17229,G17228);
  xor GNAME17241(G17241,G17242,G29641);
  xor GNAME17242(G17242,G28928,G28925);
  and GNAME17243(G17243,G28928,G29641);
  and GNAME17244(G17244,G28925,G29641);
  and GNAME17245(G17245,G28928,G28925);
  or GNAME17246(G17246,G17245,G17244,G17243);
  xor GNAME17256(G17256,G17257,G29644);
  xor GNAME17257(G17257,G28929,G28926);
  and GNAME17258(G17258,G28929,G29644);
  and GNAME17259(G17259,G28926,G29644);
  and GNAME17260(G17260,G28929,G28926);
  or GNAME17261(G17261,G17260,G17259,G17258);
  xor GNAME17271(G17271,G17272,G29647);
  xor GNAME17272(G17272,G28933,G28930);
  and GNAME17273(G17273,G28933,G29647);
  and GNAME17274(G17274,G28930,G29647);
  and GNAME17275(G17275,G28933,G28930);
  or GNAME17276(G17276,G17275,G17274,G17273);
  xor GNAME17286(G17286,G17287,G29650);
  xor GNAME17287(G17287,G28934,G28931);
  and GNAME17288(G17288,G28934,G29650);
  and GNAME17289(G17289,G28931,G29650);
  and GNAME17290(G17290,G28934,G28931);
  or GNAME17291(G17291,G17290,G17289,G17288);
  xor GNAME17301(G17301,G17302,G29653);
  xor GNAME17302(G17302,G28935,G28932);
  and GNAME17303(G17303,G28935,G29653);
  and GNAME17304(G17304,G28932,G29653);
  and GNAME17305(G17305,G28935,G28932);
  or GNAME17306(G17306,G17305,G17304,G17303);
  xor GNAME17316(G17316,G17317,G29656);
  xor GNAME17317(G17317,G28939,G28936);
  and GNAME17318(G17318,G28939,G29656);
  and GNAME17319(G17319,G28936,G29656);
  and GNAME17320(G17320,G28939,G28936);
  or GNAME17321(G17321,G17320,G17319,G17318);
  xor GNAME17331(G17331,G17332,G29659);
  xor GNAME17332(G17332,G28940,G28937);
  and GNAME17333(G17333,G28940,G29659);
  and GNAME17334(G17334,G28937,G29659);
  and GNAME17335(G17335,G28940,G28937);
  or GNAME17336(G17336,G17335,G17334,G17333);
  xor GNAME17346(G17346,G17347,G29662);
  xor GNAME17347(G17347,G28941,G28938);
  and GNAME17348(G17348,G28941,G29662);
  and GNAME17349(G17349,G28938,G29662);
  and GNAME17350(G17350,G28941,G28938);
  or GNAME17351(G17351,G17350,G17349,G17348);
  xor GNAME17361(G17361,G17362,G29665);
  xor GNAME17362(G17362,G28945,G28942);
  and GNAME17363(G17363,G28945,G29665);
  and GNAME17364(G17364,G28942,G29665);
  and GNAME17365(G17365,G28945,G28942);
  or GNAME17366(G17366,G17365,G17364,G17363);
  xor GNAME17376(G17376,G17377,G29668);
  xor GNAME17377(G17377,G28946,G28943);
  and GNAME17378(G17378,G28946,G29668);
  and GNAME17379(G17379,G28943,G29668);
  and GNAME17380(G17380,G28946,G28943);
  or GNAME17381(G17381,G17380,G17379,G17378);
  xor GNAME17391(G17391,G17392,G29671);
  xor GNAME17392(G17392,G28947,G28944);
  and GNAME17393(G17393,G28947,G29671);
  and GNAME17394(G17394,G28944,G29671);
  and GNAME17395(G17395,G28947,G28944);
  or GNAME17396(G17396,G17395,G17394,G17393);
  xor GNAME17406(G17406,G17407,G29674);
  xor GNAME17407(G17407,G28951,G28948);
  and GNAME17408(G17408,G28951,G29674);
  and GNAME17409(G17409,G28948,G29674);
  and GNAME17410(G17410,G28951,G28948);
  or GNAME17411(G17411,G17410,G17409,G17408);
  xor GNAME17421(G17421,G17422,G29677);
  xor GNAME17422(G17422,G28952,G28949);
  and GNAME17423(G17423,G28952,G29677);
  and GNAME17424(G17424,G28949,G29677);
  and GNAME17425(G17425,G28952,G28949);
  or GNAME17426(G17426,G17425,G17424,G17423);
  xor GNAME17436(G17436,G17437,G29680);
  xor GNAME17437(G17437,G28953,G28950);
  and GNAME17438(G17438,G28953,G29680);
  and GNAME17439(G17439,G28950,G29680);
  and GNAME17440(G17440,G28953,G28950);
  or GNAME17441(G17441,G17440,G17439,G17438);
  xor GNAME17451(G17451,G17452,G29683);
  xor GNAME17452(G17452,G28960,G28954);
  and GNAME17453(G17453,G28960,G29683);
  and GNAME17454(G17454,G28954,G29683);
  and GNAME17455(G17455,G28960,G28954);
  or GNAME17456(G17456,G17455,G17454,G17453);
  xor GNAME17466(G17466,G17467,G29686);
  xor GNAME17467(G17467,G28961,G28955);
  and GNAME17468(G17468,G28961,G29686);
  and GNAME17469(G17469,G28955,G29686);
  and GNAME17470(G17470,G28961,G28955);
  or GNAME17471(G17471,G17470,G17469,G17468);
  xor GNAME17481(G17481,G17482,G29689);
  xor GNAME17482(G17482,G28962,G28956);
  and GNAME17483(G17483,G28962,G29689);
  and GNAME17484(G17484,G28956,G29689);
  and GNAME17485(G17485,G28962,G28956);
  or GNAME17486(G17486,G17485,G17484,G17483);
  xor GNAME17496(G17496,G17497,G29692);
  xor GNAME17497(G17497,G28957,G31556);
  and GNAME17498(G17498,G28957,G29692);
  and GNAME17499(G17499,G31556,G29692);
  and GNAME17500(G17500,G28957,G31556);
  or GNAME17501(G17501,G17500,G17499,G17498);
  xor GNAME17511(G17511,G17512,G29695);
  xor GNAME17512(G17512,G28958,G31557);
  and GNAME17513(G17513,G28958,G29695);
  and GNAME17514(G17514,G31557,G29695);
  and GNAME17515(G17515,G28958,G31557);
  or GNAME17516(G17516,G17515,G17514,G17513);
  xor GNAME17526(G17526,G17527,G29698);
  xor GNAME17527(G17527,G28959,G31558);
  and GNAME17528(G17528,G28959,G29698);
  and GNAME17529(G17529,G31558,G29698);
  and GNAME17530(G17530,G28959,G31558);
  or GNAME17531(G17531,G17530,G17529,G17528);
  xor GNAME17541(G17541,G17542,G29701);
  xor GNAME17542(G17542,G27941,G29704);
  and GNAME17543(G17543,G27941,G29701);
  and GNAME17544(G17544,G29704,G29701);
  and GNAME17545(G17545,G27941,G29704);
  or GNAME17546(G17546,G17545,G17544,G17543);
  xor GNAME17556(G17556,G17557,G29707);
  xor GNAME17557(G17557,G27944,G29710);
  and GNAME17558(G17558,G27944,G29707);
  and GNAME17559(G17559,G29710,G29707);
  and GNAME17560(G17560,G27944,G29710);
  or GNAME17561(G17561,G17560,G17559,G17558);
  xor GNAME17571(G17571,G17572,G29713);
  xor GNAME17572(G17572,G27947,G29716);
  and GNAME17573(G17573,G27947,G29713);
  and GNAME17574(G17574,G29716,G29713);
  and GNAME17575(G17575,G27947,G29716);
  or GNAME17576(G17576,G17575,G17574,G17573);
  xor GNAME17586(G17586,G17587,G29719);
  xor GNAME17587(G17587,G27950,G29722);
  and GNAME17588(G17588,G27950,G29719);
  and GNAME17589(G17589,G29722,G29719);
  and GNAME17590(G17590,G27950,G29722);
  or GNAME17591(G17591,G17590,G17589,G17588);
  xor GNAME17601(G17601,G17602,G29725);
  xor GNAME17602(G17602,G27953,G29728);
  and GNAME17603(G17603,G27953,G29725);
  and GNAME17604(G17604,G29728,G29725);
  and GNAME17605(G17605,G27953,G29728);
  or GNAME17606(G17606,G17605,G17604,G17603);
  xor GNAME17616(G17616,G17617,G29731);
  xor GNAME17617(G17617,G27956,G29734);
  and GNAME17618(G17618,G27956,G29731);
  and GNAME17619(G17619,G29734,G29731);
  and GNAME17620(G17620,G27956,G29734);
  or GNAME17621(G17621,G17620,G17619,G17618);
  xor GNAME17631(G17631,G17632,G29773);
  xor GNAME17632(G17632,G28049,G29776);
  and GNAME17633(G17633,G28049,G29773);
  and GNAME17634(G17634,G29776,G29773);
  and GNAME17635(G17635,G28049,G29776);
  or GNAME17636(G17636,G17635,G17634,G17633);
  xor GNAME17646(G17646,G17647,G29779);
  xor GNAME17647(G17647,G28052,G29782);
  and GNAME17648(G17648,G28052,G29779);
  and GNAME17649(G17649,G29782,G29779);
  and GNAME17650(G17650,G28052,G29782);
  or GNAME17651(G17651,G17650,G17649,G17648);
  xor GNAME17661(G17661,G17662,G29785);
  xor GNAME17662(G17662,G28055,G29788);
  and GNAME17663(G17663,G28055,G29785);
  and GNAME17664(G17664,G29788,G29785);
  and GNAME17665(G17665,G28055,G29788);
  or GNAME17666(G17666,G17665,G17664,G17663);
  xor GNAME17676(G17676,G17677,G29809);
  xor GNAME17677(G17677,G28058,G29812);
  and GNAME17678(G17678,G28058,G29809);
  and GNAME17679(G17679,G29812,G29809);
  and GNAME17680(G17680,G28058,G29812);
  or GNAME17681(G17681,G17680,G17679,G17678);
  xor GNAME17691(G17691,G17692,G29815);
  xor GNAME17692(G17692,G28061,G29818);
  and GNAME17693(G17693,G28061,G29815);
  and GNAME17694(G17694,G29818,G29815);
  and GNAME17695(G17695,G28061,G29818);
  or GNAME17696(G17696,G17695,G17694,G17693);
  xor GNAME17706(G17706,G17707,G29821);
  xor GNAME17707(G17707,G28064,G29824);
  and GNAME17708(G17708,G28064,G29821);
  and GNAME17709(G17709,G29824,G29821);
  and GNAME17710(G17710,G28064,G29824);
  or GNAME17711(G17711,G17710,G17709,G17708);
  xor GNAME17721(G17721,G17722,G29845);
  xor GNAME17722(G17722,G28067,G29848);
  and GNAME17723(G17723,G28067,G29845);
  and GNAME17724(G17724,G29848,G29845);
  and GNAME17725(G17725,G28067,G29848);
  or GNAME17726(G17726,G17725,G17724,G17723);
  xor GNAME17736(G17736,G17737,G29851);
  xor GNAME17737(G17737,G28070,G29854);
  and GNAME17738(G17738,G28070,G29851);
  and GNAME17739(G17739,G29854,G29851);
  and GNAME17740(G17740,G28070,G29854);
  or GNAME17741(G17741,G17740,G17739,G17738);
  xor GNAME17751(G17751,G17752,G29857);
  xor GNAME17752(G17752,G28073,G29860);
  and GNAME17753(G17753,G28073,G29857);
  and GNAME17754(G17754,G29860,G29857);
  and GNAME17755(G17755,G28073,G29860);
  or GNAME17756(G17756,G17755,G17754,G17753);
  xor GNAME17766(G17766,G17767,G29881);
  xor GNAME17767(G17767,G28076,G29884);
  and GNAME17768(G17768,G28076,G29881);
  and GNAME17769(G17769,G29884,G29881);
  and GNAME17770(G17770,G28076,G29884);
  or GNAME17771(G17771,G17770,G17769,G17768);
  xor GNAME17781(G17781,G17782,G29887);
  xor GNAME17782(G17782,G28079,G29890);
  and GNAME17783(G17783,G28079,G29887);
  and GNAME17784(G17784,G29890,G29887);
  and GNAME17785(G17785,G28079,G29890);
  or GNAME17786(G17786,G17785,G17784,G17783);
  xor GNAME17796(G17796,G17797,G29893);
  xor GNAME17797(G17797,G28082,G29896);
  and GNAME17798(G17798,G28082,G29893);
  and GNAME17799(G17799,G29896,G29893);
  and GNAME17800(G17800,G28082,G29896);
  or GNAME17801(G17801,G17800,G17799,G17798);
  xor GNAME17811(G17811,G17812,G28216);
  xor GNAME17812(G17812,G29899,G29902);
  and GNAME17813(G17813,G29899,G28216);
  and GNAME17814(G17814,G29902,G28216);
  and GNAME17815(G17815,G29899,G29902);
  or GNAME17816(G17816,G17815,G17814,G17813);
  xor GNAME17826(G17826,G17827,G28222);
  xor GNAME17827(G17827,G29905,G29908);
  and GNAME17828(G17828,G29905,G28222);
  and GNAME17829(G17829,G29908,G28222);
  and GNAME17830(G17830,G29905,G29908);
  or GNAME17831(G17831,G17830,G17829,G17828);
  xor GNAME17841(G17841,G17842,G28228);
  xor GNAME17842(G17842,G29911,G29914);
  and GNAME17843(G17843,G29911,G28228);
  and GNAME17844(G17844,G29914,G28228);
  and GNAME17845(G17845,G29911,G29914);
  or GNAME17846(G17846,G17845,G17844,G17843);
  xor GNAME17856(G17856,G17857,G29917);
  xor GNAME17857(G17857,G28085,G29920);
  and GNAME17858(G17858,G28085,G29917);
  and GNAME17859(G17859,G29920,G29917);
  and GNAME17860(G17860,G28085,G29920);
  or GNAME17861(G17861,G17860,G17859,G17858);
  xor GNAME17871(G17871,G17872,G29923);
  xor GNAME17872(G17872,G28088,G29926);
  and GNAME17873(G17873,G28088,G29923);
  and GNAME17874(G17874,G29926,G29923);
  and GNAME17875(G17875,G28088,G29926);
  or GNAME17876(G17876,G17875,G17874,G17873);
  xor GNAME17886(G17886,G17887,G29929);
  xor GNAME17887(G17887,G28091,G29932);
  and GNAME17888(G17888,G28091,G29929);
  and GNAME17889(G17889,G29932,G29929);
  and GNAME17890(G17890,G28091,G29932);
  or GNAME17891(G17891,G17890,G17889,G17888);
  xor GNAME17901(G17901,G17902,G17231);
  xor GNAME17902(G17902,G31538,G29971);
  and GNAME17903(G17903,G31538,G17231);
  and GNAME17904(G17904,G29971,G17231);
  and GNAME17905(G17905,G31538,G29971);
  or GNAME17906(G17906,G17905,G17904,G17903);
  xor GNAME17916(G17916,G17917,G17246);
  xor GNAME17917(G17917,G31539,G29974);
  and GNAME17918(G17918,G31539,G17246);
  and GNAME17919(G17919,G29974,G17246);
  and GNAME17920(G17920,G31539,G29974);
  or GNAME17921(G17921,G17920,G17919,G17918);
  xor GNAME17931(G17931,G17932,G17261);
  xor GNAME17932(G17932,G31540,G29977);
  and GNAME17933(G17933,G31540,G17261);
  and GNAME17934(G17934,G29977,G17261);
  and GNAME17935(G17935,G31540,G29977);
  or GNAME17936(G17936,G17935,G17934,G17933);
  xor GNAME17946(G17946,G17947,G17226);
  xor GNAME17947(G17947,G29595,G18041);
  and GNAME17948(G17948,G29595,G17226);
  and GNAME17949(G17949,G18041,G17226);
  and GNAME17950(G17950,G29595,G18041);
  or GNAME17951(G17951,G17950,G17949,G17948);
  xor GNAME17961(G17961,G17962,G17241);
  xor GNAME17962(G17962,G29597,G18056);
  and GNAME17963(G17963,G29597,G17241);
  and GNAME17964(G17964,G18056,G17241);
  and GNAME17965(G17965,G29597,G18056);
  or GNAME17966(G17966,G17965,G17964,G17963);
  xor GNAME17976(G17976,G17977,G17256);
  xor GNAME17977(G17977,G29599,G18071);
  and GNAME17978(G17978,G29599,G17256);
  and GNAME17979(G17979,G18071,G17256);
  and GNAME17980(G17980,G29599,G18071);
  or GNAME17981(G17981,G17980,G17979,G17978);
  xor GNAME17991(G17991,G17992,G18086);
  xor GNAME17992(G17992,G17276,G18036);
  and GNAME17993(G17993,G17276,G18086);
  and GNAME17994(G17994,G18036,G18086);
  and GNAME17995(G17995,G17276,G18036);
  or GNAME17996(G17996,G17995,G17994,G17993);
  xor GNAME18006(G18006,G18007,G18101);
  xor GNAME18007(G18007,G17291,G18051);
  and GNAME18008(G18008,G17291,G18101);
  and GNAME18009(G18009,G18051,G18101);
  and GNAME18010(G18010,G17291,G18051);
  or GNAME18011(G18011,G18010,G18009,G18008);
  xor GNAME18021(G18021,G18022,G18116);
  xor GNAME18022(G18022,G17306,G18066);
  and GNAME18023(G18023,G17306,G18116);
  and GNAME18024(G18024,G18066,G18116);
  and GNAME18025(G18025,G17306,G18066);
  or GNAME18026(G18026,G18025,G18024,G18023);
  xor GNAME18036(G18036,G18037,G29983);
  xor GNAME18037(G18037,G31541,G29980);
  and GNAME18038(G18038,G31541,G29983);
  and GNAME18039(G18039,G29980,G29983);
  and GNAME18040(G18040,G31541,G29980);
  or GNAME18041(G18041,G18040,G18039,G18038);
  xor GNAME18051(G18051,G18052,G29989);
  xor GNAME18052(G18052,G31542,G29986);
  and GNAME18053(G18053,G31542,G29989);
  and GNAME18054(G18054,G29986,G29989);
  and GNAME18055(G18055,G31542,G29986);
  or GNAME18056(G18056,G18055,G18054,G18053);
  xor GNAME18066(G18066,G18067,G29995);
  xor GNAME18067(G18067,G31543,G29992);
  and GNAME18068(G18068,G31543,G29995);
  and GNAME18069(G18069,G29992,G29995);
  and GNAME18070(G18070,G31543,G29992);
  or GNAME18071(G18071,G18070,G18069,G18068);
  xor GNAME18081(G18081,G18082,G18221);
  xor GNAME18082(G18082,G29998,G29601);
  and GNAME18083(G18083,G29998,G18221);
  and GNAME18084(G18084,G29601,G18221);
  and GNAME18085(G18085,G29998,G29601);
  or GNAME18086(G18086,G18085,G18084,G18083);
  xor GNAME18096(G18096,G18097,G18236);
  xor GNAME18097(G18097,G30001,G29603);
  and GNAME18098(G18098,G30001,G18236);
  and GNAME18099(G18099,G29603,G18236);
  and GNAME18100(G18100,G30001,G29603);
  or GNAME18101(G18101,G18100,G18099,G18098);
  xor GNAME18111(G18111,G18112,G18251);
  xor GNAME18112(G18112,G30004,G29605);
  and GNAME18113(G18113,G30004,G18251);
  and GNAME18114(G18114,G29605,G18251);
  and GNAME18115(G18115,G30004,G29605);
  or GNAME18116(G18116,G18115,G18114,G18113);
  xor GNAME18126(G18126,G18127,G18081);
  xor GNAME18127(G18127,G17271,G18176);
  and GNAME18128(G18128,G17271,G18081);
  and GNAME18129(G18129,G18176,G18081);
  and GNAME18130(G18130,G17271,G18176);
  or GNAME18131(G18131,G18130,G18129,G18128);
  xor GNAME18141(G18141,G18142,G18096);
  xor GNAME18142(G18142,G17286,G18191);
  and GNAME18143(G18143,G17286,G18096);
  and GNAME18144(G18144,G18191,G18096);
  and GNAME18145(G18145,G17286,G18191);
  or GNAME18146(G18146,G18145,G18144,G18143);
  xor GNAME18156(G18156,G18157,G18111);
  xor GNAME18157(G18157,G17301,G18206);
  and GNAME18158(G18158,G17301,G18111);
  and GNAME18159(G18159,G18206,G18111);
  and GNAME18160(G18160,G17301,G18206);
  or GNAME18161(G18161,G18160,G18159,G18158);
  xor GNAME18171(G18171,G18172,G18266);
  xor GNAME18172(G18172,G30007,G17321);
  and GNAME18173(G18173,G30007,G18266);
  and GNAME18174(G18174,G17321,G18266);
  and GNAME18175(G18175,G30007,G17321);
  or GNAME18176(G18176,G18175,G18174,G18173);
  xor GNAME18186(G18186,G18187,G18281);
  xor GNAME18187(G18187,G30010,G17336);
  and GNAME18188(G18188,G30010,G18281);
  and GNAME18189(G18189,G17336,G18281);
  and GNAME18190(G18190,G30010,G17336);
  or GNAME18191(G18191,G18190,G18189,G18188);
  xor GNAME18201(G18201,G18202,G18296);
  xor GNAME18202(G18202,G30013,G17351);
  and GNAME18203(G18203,G30013,G18296);
  and GNAME18204(G18204,G17351,G18296);
  and GNAME18205(G18205,G30013,G17351);
  or GNAME18206(G18206,G18205,G18204,G18203);
  xor GNAME18216(G18216,G18217,G30019);
  xor GNAME18217(G18217,G31544,G30016);
  and GNAME18218(G18218,G31544,G30019);
  and GNAME18219(G18219,G30016,G30019);
  and GNAME18220(G18220,G31544,G30016);
  or GNAME18221(G18221,G18220,G18219,G18218);
  xor GNAME18231(G18231,G18232,G30025);
  xor GNAME18232(G18232,G31545,G30022);
  and GNAME18233(G18233,G31545,G30025);
  and GNAME18234(G18234,G30022,G30025);
  and GNAME18235(G18235,G31545,G30022);
  or GNAME18236(G18236,G18235,G18234,G18233);
  xor GNAME18246(G18246,G18247,G30031);
  xor GNAME18247(G18247,G31546,G30028);
  and GNAME18248(G18248,G31546,G30031);
  and GNAME18249(G18249,G30028,G30031);
  and GNAME18250(G18250,G31546,G30028);
  or GNAME18251(G18251,G18250,G18249,G18248);
  xor GNAME18261(G18261,G18262,G29607);
  xor GNAME18262(G18262,G30034,G30037);
  and GNAME18263(G18263,G30034,G29607);
  and GNAME18264(G18264,G30037,G29607);
  and GNAME18265(G18265,G30034,G30037);
  or GNAME18266(G18266,G18265,G18264,G18263);
  xor GNAME18276(G18276,G18277,G29609);
  xor GNAME18277(G18277,G30040,G30043);
  and GNAME18278(G18278,G30040,G29609);
  and GNAME18279(G18279,G30043,G29609);
  and GNAME18280(G18280,G30040,G30043);
  or GNAME18281(G18281,G18280,G18279,G18278);
  xor GNAME18291(G18291,G18292,G29611);
  xor GNAME18292(G18292,G30046,G30049);
  and GNAME18293(G18293,G30046,G29611);
  and GNAME18294(G18294,G30049,G29611);
  and GNAME18295(G18295,G30046,G30049);
  or GNAME18296(G18296,G18295,G18294,G18293);
  xor GNAME18306(G18306,G18307,G18261);
  xor GNAME18307(G18307,G18356,G17316);
  and GNAME18308(G18308,G18356,G18261);
  and GNAME18309(G18309,G17316,G18261);
  and GNAME18310(G18310,G18356,G17316);
  or GNAME18311(G18311,G18310,G18309,G18308);
  xor GNAME18321(G18321,G18322,G18276);
  xor GNAME18322(G18322,G18371,G17331);
  and GNAME18323(G18323,G18371,G18276);
  and GNAME18324(G18324,G17331,G18276);
  and GNAME18325(G18325,G18371,G17331);
  or GNAME18326(G18326,G18325,G18324,G18323);
  xor GNAME18336(G18336,G18337,G18291);
  xor GNAME18337(G18337,G18386,G17346);
  and GNAME18338(G18338,G18386,G18291);
  and GNAME18339(G18339,G17346,G18291);
  and GNAME18340(G18340,G18386,G17346);
  or GNAME18341(G18341,G18340,G18339,G18338);
  xor GNAME18351(G18351,G18352,G30055);
  xor GNAME18352(G18352,G31547,G30052);
  and GNAME18353(G18353,G31547,G30055);
  and GNAME18354(G18354,G30052,G30055);
  and GNAME18355(G18355,G31547,G30052);
  or GNAME18356(G18356,G18355,G18354,G18353);
  xor GNAME18366(G18366,G18367,G30061);
  xor GNAME18367(G18367,G31548,G30058);
  and GNAME18368(G18368,G31548,G30061);
  and GNAME18369(G18369,G30058,G30061);
  and GNAME18370(G18370,G31548,G30058);
  or GNAME18371(G18371,G18370,G18369,G18368);
  xor GNAME18381(G18381,G18382,G30067);
  xor GNAME18382(G18382,G31549,G30064);
  and GNAME18383(G18383,G31549,G30067);
  and GNAME18384(G18384,G30064,G30067);
  and GNAME18385(G18385,G31549,G30064);
  or GNAME18386(G18386,G18385,G18384,G18383);
  xor GNAME18396(G18396,G18397,G17366);
  xor GNAME18397(G18397,G30070,G30073);
  and GNAME18398(G18398,G30070,G17366);
  and GNAME18399(G18399,G30073,G17366);
  and GNAME18400(G18400,G30070,G30073);
  or GNAME18401(G18401,G18400,G18399,G18398);
  xor GNAME18411(G18411,G18412,G17381);
  xor GNAME18412(G18412,G30076,G30079);
  and GNAME18413(G18413,G30076,G17381);
  and GNAME18414(G18414,G30079,G17381);
  and GNAME18415(G18415,G30076,G30079);
  or GNAME18416(G18416,G18415,G18414,G18413);
  xor GNAME18426(G18426,G18427,G17396);
  xor GNAME18427(G18427,G30082,G30085);
  and GNAME18428(G18428,G30082,G17396);
  and GNAME18429(G18429,G30085,G17396);
  and GNAME18430(G18430,G30082,G30085);
  or GNAME18431(G18431,G18430,G18429,G18428);
  xor GNAME18441(G18441,G18442,G18536);
  xor GNAME18442(G18442,G17361,G18666);
  and GNAME18443(G18443,G17361,G18536);
  and GNAME18444(G18444,G18666,G18536);
  and GNAME18445(G18445,G17361,G18666);
  or GNAME18446(G18446,G18445,G18444,G18443);
  xor GNAME18456(G18456,G18457,G18551);
  xor GNAME18457(G18457,G17376,G18681);
  and GNAME18458(G18458,G17376,G18551);
  and GNAME18459(G18459,G18681,G18551);
  and GNAME18460(G18460,G17376,G18681);
  or GNAME18461(G18461,G18460,G18459,G18458);
  xor GNAME18471(G18471,G18472,G18566);
  xor GNAME18472(G18472,G17391,G18696);
  and GNAME18473(G18473,G17391,G18566);
  and GNAME18474(G18474,G18696,G18566);
  and GNAME18475(G18475,G17391,G18696);
  or GNAME18476(G18476,G18475,G18474,G18473);
  xor GNAME18486(G18486,G18487,G30091);
  xor GNAME18487(G18487,G31550,G30088);
  and GNAME18488(G18488,G31550,G30091);
  and GNAME18489(G18489,G30088,G30091);
  and GNAME18490(G18490,G31550,G30088);
  or GNAME18491(G18491,G18490,G18489,G18488);
  xor GNAME18501(G18501,G18502,G30097);
  xor GNAME18502(G18502,G31551,G30094);
  and GNAME18503(G18503,G31551,G30097);
  and GNAME18504(G18504,G30094,G30097);
  and GNAME18505(G18505,G31551,G30094);
  or GNAME18506(G18506,G18505,G18504,G18503);
  xor GNAME18516(G18516,G18517,G30103);
  xor GNAME18517(G18517,G31552,G30100);
  and GNAME18518(G18518,G31552,G30103);
  and GNAME18519(G18519,G30100,G30103);
  and GNAME18520(G18520,G31552,G30100);
  or GNAME18521(G18521,G18520,G18519,G18518);
  xor GNAME18531(G18531,G18532,G18486);
  xor GNAME18532(G18532,G17411,G18716);
  and GNAME18533(G18533,G17411,G18486);
  and GNAME18534(G18534,G18716,G18486);
  and GNAME18535(G18535,G17411,G18716);
  or GNAME18536(G18536,G18535,G18534,G18533);
  xor GNAME18546(G18546,G18547,G18501);
  xor GNAME18547(G18547,G17426,G18731);
  and GNAME18548(G18548,G17426,G18501);
  and GNAME18549(G18549,G18731,G18501);
  and GNAME18550(G18550,G17426,G18731);
  or GNAME18551(G18551,G18550,G18549,G18548);
  xor GNAME18561(G18561,G18562,G18516);
  xor GNAME18562(G18562,G17441,G18746);
  and GNAME18563(G18563,G17441,G18516);
  and GNAME18564(G18564,G18746,G18516);
  and GNAME18565(G18565,G17441,G18746);
  or GNAME18566(G18566,G18565,G18564,G18563);
  xor GNAME18576(G18576,G18577,G18626);
  xor GNAME18577(G18577,G30106,G18491);
  and GNAME18578(G18578,G30106,G18626);
  and GNAME18579(G18579,G18491,G18626);
  and GNAME18580(G18580,G30106,G18491);
  or GNAME18581(G18581,G18580,G18579,G18578);
  xor GNAME18591(G18591,G18592,G18641);
  xor GNAME18592(G18592,G30109,G18506);
  and GNAME18593(G18593,G30109,G18641);
  and GNAME18594(G18594,G18506,G18641);
  and GNAME18595(G18595,G30109,G18506);
  or GNAME18596(G18596,G18595,G18594,G18593);
  xor GNAME18606(G18606,G18607,G18656);
  xor GNAME18607(G18607,G30112,G18521);
  and GNAME18608(G18608,G30112,G18656);
  and GNAME18609(G18609,G18521,G18656);
  and GNAME18610(G18610,G30112,G18521);
  or GNAME18611(G18611,G18610,G18609,G18608);
  xor GNAME18621(G18621,G18622,G30121);
  xor GNAME18622(G18622,G30115,G30118);
  and GNAME18623(G18623,G30115,G30121);
  and GNAME18624(G18624,G30118,G30121);
  and GNAME18625(G18625,G30115,G30118);
  or GNAME18626(G18626,G18625,G18624,G18623);
  xor GNAME18636(G18636,G18637,G30130);
  xor GNAME18637(G18637,G30124,G30127);
  and GNAME18638(G18638,G30124,G30130);
  and GNAME18639(G18639,G30127,G30130);
  and GNAME18640(G18640,G30124,G30127);
  or GNAME18641(G18641,G18640,G18639,G18638);
  xor GNAME18651(G18651,G18652,G30139);
  xor GNAME18652(G18652,G30133,G30136);
  and GNAME18653(G18653,G30133,G30139);
  and GNAME18654(G18654,G30136,G30139);
  and GNAME18655(G18655,G30133,G30136);
  or GNAME18656(G18656,G18655,G18654,G18653);
  xor GNAME18666(G18666,G18667,G29613);
  xor GNAME18667(G18667,G30142,G30145);
  and GNAME18668(G18668,G30142,G29613);
  and GNAME18669(G18669,G30145,G29613);
  and GNAME18670(G18670,G30142,G30145);
  or GNAME18671(G18671,G18670,G18669,G18668);
  xor GNAME18681(G18681,G18682,G29615);
  xor GNAME18682(G18682,G30148,G30151);
  and GNAME18683(G18683,G30148,G29615);
  and GNAME18684(G18684,G30151,G29615);
  and GNAME18685(G18685,G30148,G30151);
  or GNAME18686(G18686,G18685,G18684,G18683);
  xor GNAME18696(G18696,G18697,G29617);
  xor GNAME18697(G18697,G30154,G30157);
  and GNAME18698(G18698,G30154,G29617);
  and GNAME18699(G18699,G30157,G29617);
  and GNAME18700(G18700,G30154,G30157);
  or GNAME18701(G18701,G18700,G18699,G18698);
  xor GNAME18711(G18711,G18712,G29619);
  xor GNAME18712(G18712,G30160,G30163);
  and GNAME18713(G18713,G30160,G29619);
  and GNAME18714(G18714,G30163,G29619);
  and GNAME18715(G18715,G30160,G30163);
  or GNAME18716(G18716,G18715,G18714,G18713);
  xor GNAME18726(G18726,G18727,G29621);
  xor GNAME18727(G18727,G30166,G30169);
  and GNAME18728(G18728,G30166,G29621);
  and GNAME18729(G18729,G30169,G29621);
  and GNAME18730(G18730,G30166,G30169);
  or GNAME18731(G18731,G18730,G18729,G18728);
  xor GNAME18741(G18741,G18742,G29623);
  xor GNAME18742(G18742,G30172,G30175);
  and GNAME18743(G18743,G30172,G29623);
  and GNAME18744(G18744,G30175,G29623);
  and GNAME18745(G18745,G30172,G30175);
  or GNAME18746(G18746,G18745,G18744,G18743);
  xor GNAME18756(G18756,G18757,G18806);
  xor GNAME18757(G18757,G30178,G30181);
  and GNAME18758(G18758,G30178,G18806);
  and GNAME18759(G18759,G30181,G18806);
  and GNAME18760(G18760,G30178,G30181);
  or GNAME18761(G18761,G18760,G18759,G18758);
  xor GNAME18771(G18771,G18772,G18821);
  xor GNAME18772(G18772,G30184,G30187);
  and GNAME18773(G18773,G30184,G18821);
  and GNAME18774(G18774,G30187,G18821);
  and GNAME18775(G18775,G30184,G30187);
  or GNAME18776(G18776,G18775,G18774,G18773);
  xor GNAME18786(G18786,G18787,G18836);
  xor GNAME18787(G18787,G30190,G30193);
  and GNAME18788(G18788,G30190,G18836);
  and GNAME18789(G18789,G30193,G18836);
  and GNAME18790(G18790,G30190,G30193);
  or GNAME18791(G18791,G18790,G18789,G18788);
  xor GNAME18801(G18801,G18802,G30199);
  xor GNAME18802(G18802,G31553,G30196);
  and GNAME18803(G18803,G31553,G30199);
  and GNAME18804(G18804,G30196,G30199);
  and GNAME18805(G18805,G31553,G30196);
  or GNAME18806(G18806,G18805,G18804,G18803);
  xor GNAME18816(G18816,G18817,G30205);
  xor GNAME18817(G18817,G31554,G30202);
  and GNAME18818(G18818,G31554,G30205);
  and GNAME18819(G18819,G30202,G30205);
  and GNAME18820(G18820,G31554,G30202);
  or GNAME18821(G18821,G18820,G18819,G18818);
  xor GNAME18831(G18831,G18832,G30211);
  xor GNAME18832(G18832,G31555,G30208);
  and GNAME18833(G18833,G31555,G30211);
  and GNAME18834(G18834,G30208,G30211);
  and GNAME18835(G18835,G31555,G30208);
  or GNAME18836(G18836,G18835,G18834,G18833);
  xor GNAME18846(G18846,G18847,G18711);
  xor GNAME18847(G18847,G18896,G17406);
  and GNAME18848(G18848,G18896,G18711);
  and GNAME18849(G18849,G17406,G18711);
  and GNAME18850(G18850,G18896,G17406);
  or GNAME18851(G18851,G18850,G18849,G18848);
  xor GNAME18861(G18861,G18862,G18726);
  xor GNAME18862(G18862,G18911,G17421);
  and GNAME18863(G18863,G18911,G18726);
  and GNAME18864(G18864,G17421,G18726);
  and GNAME18865(G18865,G18911,G17421);
  or GNAME18866(G18866,G18865,G18864,G18863);
  xor GNAME18876(G18876,G18877,G18741);
  xor GNAME18877(G18877,G18926,G17436);
  and GNAME18878(G18878,G18926,G18741);
  and GNAME18879(G18879,G17436,G18741);
  and GNAME18880(G18880,G18926,G17436);
  or GNAME18881(G18881,G18880,G18879,G18878);
  xor GNAME18891(G18891,G18892,G30220);
  xor GNAME18892(G18892,G30214,G30217);
  and GNAME18893(G18893,G30214,G30220);
  and GNAME18894(G18894,G30217,G30220);
  and GNAME18895(G18895,G30214,G30217);
  or GNAME18896(G18896,G18895,G18894,G18893);
  xor GNAME18906(G18906,G18907,G30229);
  xor GNAME18907(G18907,G30223,G30226);
  and GNAME18908(G18908,G30223,G30229);
  and GNAME18909(G18909,G30226,G30229);
  and GNAME18910(G18910,G30223,G30226);
  or GNAME18911(G18911,G18910,G18909,G18908);
  xor GNAME18921(G18921,G18922,G30238);
  xor GNAME18922(G18922,G30232,G30235);
  and GNAME18923(G18923,G30232,G30238);
  and GNAME18924(G18924,G30235,G30238);
  and GNAME18925(G18925,G30232,G30235);
  or GNAME18926(G18926,G18925,G18924,G18923);
  xor GNAME18936(G18936,G18937,G29625);
  xor GNAME18937(G18937,G30241,G30244);
  and GNAME18938(G18938,G30241,G29625);
  and GNAME18939(G18939,G30244,G29625);
  and GNAME18940(G18940,G30241,G30244);
  or GNAME18941(G18941,G18940,G18939,G18938);
  xor GNAME18951(G18951,G18952,G29627);
  xor GNAME18952(G18952,G30247,G30250);
  and GNAME18953(G18953,G30247,G29627);
  and GNAME18954(G18954,G30250,G29627);
  and GNAME18955(G18955,G30247,G30250);
  or GNAME18956(G18956,G18955,G18954,G18953);
  xor GNAME18966(G18966,G18967,G29629);
  xor GNAME18967(G18967,G30253,G30256);
  and GNAME18968(G18968,G30253,G29629);
  and GNAME18969(G18969,G30256,G29629);
  and GNAME18970(G18970,G30253,G30256);
  or GNAME18971(G18971,G18970,G18969,G18968);
  xor GNAME18981(G18981,G18982,G18941);
  xor GNAME18982(G18982,G30259,G17456);
  and GNAME18983(G18983,G30259,G18941);
  and GNAME18984(G18984,G17456,G18941);
  and GNAME18985(G18985,G30259,G17456);
  or GNAME18986(G18986,G18985,G18984,G18983);
  xor GNAME18996(G18996,G18997,G19091);
  xor GNAME18997(G18997,G17501,G19256);
  and GNAME18998(G18998,G17501,G19091);
  and GNAME18999(G18999,G19256,G19091);
  and GNAME19000(G19000,G17501,G19256);
  or GNAME19001(G19001,G19000,G18999,G18998);
  xor GNAME19011(G19011,G19012,G18956);
  xor GNAME19012(G19012,G30262,G17471);
  and GNAME19013(G19013,G30262,G18956);
  and GNAME19014(G19014,G17471,G18956);
  and GNAME19015(G19015,G30262,G17471);
  or GNAME19016(G19016,G19015,G19014,G19013);
  xor GNAME19026(G19026,G19027,G18971);
  xor GNAME19027(G19027,G30265,G17486);
  and GNAME19028(G19028,G30265,G18971);
  and GNAME19029(G19029,G17486,G18971);
  and GNAME19030(G19030,G30265,G17486);
  or GNAME19031(G19031,G19030,G19029,G19028);
  xor GNAME19041(G19041,G19042,G19136);
  xor GNAME19042(G19042,G17516,G19271);
  and GNAME19043(G19043,G17516,G19136);
  and GNAME19044(G19044,G19271,G19136);
  and GNAME19045(G19045,G17516,G19271);
  or GNAME19046(G19046,G19045,G19044,G19043);
  xor GNAME19056(G19056,G19057,G19151);
  xor GNAME19057(G19057,G17531,G19286);
  and GNAME19058(G19058,G17531,G19151);
  and GNAME19059(G19059,G19286,G19151);
  and GNAME19060(G19060,G17531,G19286);
  or GNAME19061(G19061,G19060,G19059,G19058);
  xor GNAME19071(G19071,G19072,G30274);
  xor GNAME19072(G19072,G30268,G30271);
  and GNAME19073(G19073,G30268,G30274);
  and GNAME19074(G19074,G30271,G30274);
  and GNAME19075(G19075,G30268,G30271);
  or GNAME19076(G19076,G19075,G19074,G19073);
  xor GNAME19086(G19086,G19087,G30283);
  xor GNAME19087(G19087,G30277,G30280);
  and GNAME19088(G19088,G30277,G30283);
  and GNAME19089(G19089,G30280,G30283);
  and GNAME19090(G19090,G30277,G30280);
  or GNAME19091(G19091,G19090,G19089,G19088);
  xor GNAME19101(G19101,G19102,G30292);
  xor GNAME19102(G19102,G30286,G30289);
  and GNAME19103(G19103,G30286,G30292);
  and GNAME19104(G19104,G30289,G30292);
  and GNAME19105(G19105,G30286,G30289);
  or GNAME19106(G19106,G19105,G19104,G19103);
  xor GNAME19116(G19116,G19117,G30301);
  xor GNAME19117(G19117,G30295,G30298);
  and GNAME19118(G19118,G30295,G30301);
  and GNAME19119(G19119,G30298,G30301);
  and GNAME19120(G19120,G30295,G30298);
  or GNAME19121(G19121,G19120,G19119,G19118);
  xor GNAME19131(G19131,G19132,G30310);
  xor GNAME19132(G19132,G30304,G30307);
  and GNAME19133(G19133,G30304,G30310);
  and GNAME19134(G19134,G30307,G30310);
  and GNAME19135(G19135,G30304,G30307);
  or GNAME19136(G19136,G19135,G19134,G19133);
  xor GNAME19146(G19146,G19147,G30319);
  xor GNAME19147(G19147,G30313,G30316);
  and GNAME19148(G19148,G30313,G30319);
  and GNAME19149(G19149,G30316,G30319);
  and GNAME19150(G19150,G30313,G30316);
  or GNAME19151(G19151,G19150,G19149,G19148);
  xor GNAME19161(G19161,G19162,G18936);
  xor GNAME19162(G19162,G17451,G19071);
  and GNAME19163(G19163,G17451,G18936);
  and GNAME19164(G19164,G19071,G18936);
  and GNAME19165(G19165,G17451,G19071);
  or GNAME19166(G19166,G19165,G19164,G19163);
  xor GNAME19176(G19176,G19177,G19251);
  xor GNAME19177(G19177,G17496,G19086);
  and GNAME19178(G19178,G17496,G19251);
  and GNAME19179(G19179,G19086,G19251);
  and GNAME19180(G19180,G17496,G19086);
  or GNAME19181(G19181,G19180,G19179,G19178);
  xor GNAME19191(G19191,G19192,G18951);
  xor GNAME19192(G19192,G17466,G19101);
  and GNAME19193(G19193,G17466,G18951);
  and GNAME19194(G19194,G19101,G18951);
  and GNAME19195(G19195,G17466,G19101);
  or GNAME19196(G19196,G19195,G19194,G19193);
  xor GNAME19206(G19206,G19207,G19266);
  xor GNAME19207(G19207,G17511,G19131);
  and GNAME19208(G19208,G17511,G19266);
  and GNAME19209(G19209,G19131,G19266);
  and GNAME19210(G19210,G17511,G19131);
  or GNAME19211(G19211,G19210,G19209,G19208);
  xor GNAME19221(G19221,G19222,G18966);
  xor GNAME19222(G19222,G17481,G19116);
  and GNAME19223(G19223,G17481,G18966);
  and GNAME19224(G19224,G19116,G18966);
  and GNAME19225(G19225,G17481,G19116);
  or GNAME19226(G19226,G19225,G19224,G19223);
  xor GNAME19236(G19236,G19237,G19281);
  xor GNAME19237(G19237,G17526,G19146);
  and GNAME19238(G19238,G17526,G19281);
  and GNAME19239(G19239,G19146,G19281);
  and GNAME19240(G19240,G17526,G19146);
  or GNAME19241(G19241,G19240,G19239,G19238);
  xor GNAME19251(G19251,G19252,G30328);
  xor GNAME19252(G19252,G30322,G30325);
  and GNAME19253(G19253,G30322,G30328);
  and GNAME19254(G19254,G30325,G30328);
  and GNAME19255(G19255,G30322,G30325);
  or GNAME19256(G19256,G19255,G19254,G19253);
  xor GNAME19266(G19266,G19267,G30337);
  xor GNAME19267(G19267,G30331,G30334);
  and GNAME19268(G19268,G30331,G30337);
  and GNAME19269(G19269,G30334,G30337);
  and GNAME19270(G19270,G30331,G30334);
  or GNAME19271(G19271,G19270,G19269,G19268);
  xor GNAME19281(G19281,G19282,G30346);
  xor GNAME19282(G19282,G30340,G30343);
  and GNAME19283(G19283,G30340,G30346);
  and GNAME19284(G19284,G30343,G30346);
  and GNAME19285(G19285,G30340,G30343);
  or GNAME19286(G19286,G19285,G19284,G19283);
  xor GNAME19296(G19296,G19297,G29631);
  xor GNAME19297(G19297,G30349,G30352);
  and GNAME19298(G19298,G30349,G29631);
  and GNAME19299(G19299,G30352,G29631);
  and GNAME19300(G19300,G30349,G30352);
  or GNAME19301(G19301,G19300,G19299,G19298);
  xor GNAME19311(G19311,G19312,G29633);
  xor GNAME19312(G19312,G30355,G30358);
  and GNAME19313(G19313,G30355,G29633);
  and GNAME19314(G19314,G30358,G29633);
  and GNAME19315(G19315,G30355,G30358);
  or GNAME19316(G19316,G19315,G19314,G19313);
  xor GNAME19326(G19326,G19327,G29635);
  xor GNAME19327(G19327,G30361,G30364);
  and GNAME19328(G19328,G30361,G29635);
  and GNAME19329(G19329,G30364,G29635);
  and GNAME19330(G19330,G30361,G30364);
  or GNAME19331(G19331,G19330,G19329,G19328);
  xor GNAME19341(G19341,G19342,G30373);
  xor GNAME19342(G19342,G30367,G30370);
  and GNAME19343(G19343,G30367,G30373);
  and GNAME19344(G19344,G30370,G30373);
  and GNAME19345(G19345,G30367,G30370);
  or GNAME19346(G19346,G19345,G19344,G19343);
  xor GNAME19356(G19356,G19357,G30382);
  xor GNAME19357(G19357,G30376,G30379);
  and GNAME19358(G19358,G30376,G30382);
  and GNAME19359(G19359,G30379,G30382);
  and GNAME19360(G19360,G30376,G30379);
  or GNAME19361(G19361,G19360,G19359,G19358);
  xor GNAME19371(G19371,G19372,G30391);
  xor GNAME19372(G19372,G30385,G30388);
  and GNAME19373(G19373,G30385,G30391);
  and GNAME19374(G19374,G30388,G30391);
  and GNAME19375(G19375,G30385,G30388);
  or GNAME19376(G19376,G19375,G19374,G19373);
  xor GNAME19386(G19386,G19387,G30394);
  xor GNAME19387(G19387,G28963,G30397);
  and GNAME19388(G19388,G28963,G30394);
  and GNAME19389(G19389,G30397,G30394);
  and GNAME19390(G19390,G28963,G30397);
  or GNAME19391(G19391,G19390,G19389,G19388);
  xor GNAME19401(G19401,G19402,G30400);
  xor GNAME19402(G19402,G28964,G30403);
  and GNAME19403(G19403,G28964,G30400);
  and GNAME19404(G19404,G30403,G30400);
  and GNAME19405(G19405,G28964,G30403);
  or GNAME19406(G19406,G19405,G19404,G19403);
  xor GNAME19416(G19416,G19417,G30406);
  xor GNAME19417(G19417,G28965,G30409);
  and GNAME19418(G19418,G28965,G30406);
  and GNAME19419(G19419,G30409,G30406);
  and GNAME19420(G19420,G28965,G30409);
  or GNAME19421(G19421,G19420,G19419,G19418);
  xor GNAME19431(G19431,G19432,G30415);
  xor GNAME19432(G19432,G31556,G30412);
  and GNAME19433(G19433,G31556,G30415);
  and GNAME19434(G19434,G30412,G30415);
  and GNAME19435(G19435,G31556,G30412);
  or GNAME19436(G19436,G19435,G19434,G19433);
  xor GNAME19446(G19446,G19447,G30421);
  xor GNAME19447(G19447,G31557,G30418);
  and GNAME19448(G19448,G31557,G30421);
  and GNAME19449(G19449,G30418,G30421);
  and GNAME19450(G19450,G31557,G30418);
  or GNAME19451(G19451,G19450,G19449,G19448);
  xor GNAME19461(G19461,G19462,G30427);
  xor GNAME19462(G19462,G31558,G30424);
  and GNAME19463(G19463,G31558,G30427);
  and GNAME19464(G19464,G30424,G30427);
  and GNAME19465(G19465,G31558,G30424);
  or GNAME19466(G19466,G19465,G19464,G19463);
  xor GNAME19476(G19476,G19477,G30436);
  xor GNAME19477(G19477,G30430,G30433);
  and GNAME19478(G19478,G30430,G30436);
  and GNAME19479(G19479,G30433,G30436);
  and GNAME19480(G19480,G30430,G30433);
  or GNAME19481(G19481,G19480,G19479,G19478);
  xor GNAME19491(G19491,G19492,G30445);
  xor GNAME19492(G19492,G30439,G30442);
  and GNAME19493(G19493,G30439,G30445);
  and GNAME19494(G19494,G30442,G30445);
  and GNAME19495(G19495,G30439,G30442);
  or GNAME19496(G19496,G19495,G19494,G19493);
  xor GNAME19506(G19506,G19507,G30454);
  xor GNAME19507(G19507,G30448,G30451);
  and GNAME19508(G19508,G30448,G30454);
  and GNAME19509(G19509,G30451,G30454);
  and GNAME19510(G19510,G30448,G30451);
  or GNAME19511(G19511,G19510,G19509,G19508);
  xor GNAME19521(G19521,G19522,G30463);
  xor GNAME19522(G19522,G30457,G30460);
  and GNAME19523(G19523,G30457,G30463);
  and GNAME19524(G19524,G30460,G30463);
  and GNAME19525(G19525,G30457,G30460);
  or GNAME19526(G19526,G19525,G19524,G19523);
  xor GNAME19536(G19536,G19537,G30472);
  xor GNAME19537(G19537,G30466,G30469);
  and GNAME19538(G19538,G30466,G30472);
  and GNAME19539(G19539,G30469,G30472);
  and GNAME19540(G19540,G30466,G30469);
  or GNAME19541(G19541,G19540,G19539,G19538);
  xor GNAME19551(G19551,G19552,G30481);
  xor GNAME19552(G19552,G30475,G30478);
  and GNAME19553(G19553,G30475,G30481);
  and GNAME19554(G19554,G30478,G30481);
  and GNAME19555(G19555,G30475,G30478);
  or GNAME19556(G19556,G19555,G19554,G19553);
  xor GNAME19566(G19566,G19567,G30490);
  xor GNAME19567(G19567,G30484,G30487);
  and GNAME19568(G19568,G30484,G30490);
  and GNAME19569(G19569,G30487,G30490);
  and GNAME19570(G19570,G30484,G30487);
  or GNAME19571(G19571,G19570,G19569,G19568);
  xor GNAME19581(G19581,G19582,G30499);
  xor GNAME19582(G19582,G30493,G30496);
  and GNAME19583(G19583,G30493,G30499);
  and GNAME19584(G19584,G30496,G30499);
  and GNAME19585(G19585,G30493,G30496);
  or GNAME19586(G19586,G19585,G19584,G19583);
  xor GNAME19596(G19596,G19597,G30508);
  xor GNAME19597(G19597,G30502,G30505);
  and GNAME19598(G19598,G30502,G30508);
  and GNAME19599(G19599,G30505,G30508);
  and GNAME19600(G19600,G30502,G30505);
  or GNAME19601(G19601,G19600,G19599,G19598);
  xor GNAME19611(G19611,G19612,G30517);
  xor GNAME19612(G19612,G30511,G30514);
  and GNAME19613(G19613,G30511,G30517);
  and GNAME19614(G19614,G30514,G30517);
  and GNAME19615(G19615,G30511,G30514);
  or GNAME19616(G19616,G19615,G19614,G19613);
  xor GNAME19626(G19626,G19627,G30526);
  xor GNAME19627(G19627,G30520,G30523);
  and GNAME19628(G19628,G30520,G30526);
  and GNAME19629(G19629,G30523,G30526);
  and GNAME19630(G19630,G30520,G30523);
  or GNAME19631(G19631,G19630,G19629,G19628);
  xor GNAME19641(G19641,G19642,G30535);
  xor GNAME19642(G19642,G30529,G30532);
  and GNAME19643(G19643,G30529,G30535);
  and GNAME19644(G19644,G30532,G30535);
  and GNAME19645(G19645,G30529,G30532);
  or GNAME19646(G19646,G19645,G19644,G19643);
  xor GNAME19656(G19656,G19657,G30538);
  xor GNAME19657(G19657,G28966,G30541);
  and GNAME19658(G19658,G28966,G30538);
  and GNAME19659(G19659,G30541,G30538);
  and GNAME19660(G19660,G28966,G30541);
  or GNAME19661(G19661,G19660,G19659,G19658);
  xor GNAME19671(G19671,G19672,G30544);
  xor GNAME19672(G19672,G28967,G30547);
  and GNAME19673(G19673,G28967,G30544);
  and GNAME19674(G19674,G30547,G30544);
  and GNAME19675(G19675,G28967,G30547);
  or GNAME19676(G19676,G19675,G19674,G19673);
  xor GNAME19686(G19686,G19687,G30550);
  xor GNAME19687(G19687,G28968,G30553);
  and GNAME19688(G19688,G28968,G30550);
  and GNAME19689(G19689,G30553,G30550);
  and GNAME19690(G19690,G28968,G30553);
  or GNAME19691(G19691,G19690,G19689,G19688);
  xor GNAME19701(G19701,G19702,G30556);
  xor GNAME19702(G19702,G28969,G30559);
  and GNAME19703(G19703,G28969,G30556);
  and GNAME19704(G19704,G30559,G30556);
  and GNAME19705(G19705,G28969,G30559);
  or GNAME19706(G19706,G19705,G19704,G19703);
  xor GNAME19716(G19716,G19717,G30562);
  xor GNAME19717(G19717,G28970,G30565);
  and GNAME19718(G19718,G28970,G30562);
  and GNAME19719(G19719,G30565,G30562);
  and GNAME19720(G19720,G28970,G30565);
  or GNAME19721(G19721,G19720,G19719,G19718);
  xor GNAME19731(G19731,G19732,G30568);
  xor GNAME19732(G19732,G28971,G30571);
  and GNAME19733(G19733,G28971,G30568);
  and GNAME19734(G19734,G30571,G30568);
  and GNAME19735(G19735,G28971,G30571);
  or GNAME19736(G19736,G19735,G19734,G19733);
  xor GNAME19746(G19746,G19747,G30580);
  xor GNAME19747(G19747,G30574,G30577);
  and GNAME19748(G19748,G30574,G30580);
  and GNAME19749(G19749,G30577,G30580);
  and GNAME19750(G19750,G30574,G30577);
  or GNAME19751(G19751,G19750,G19749,G19748);
  xor GNAME19761(G19761,G19762,G30589);
  xor GNAME19762(G19762,G30583,G30586);
  and GNAME19763(G19763,G30583,G30589);
  and GNAME19764(G19764,G30586,G30589);
  and GNAME19765(G19765,G30583,G30586);
  or GNAME19766(G19766,G19765,G19764,G19763);
  xor GNAME19776(G19776,G19777,G30598);
  xor GNAME19777(G19777,G30592,G30595);
  and GNAME19778(G19778,G30592,G30598);
  and GNAME19779(G19779,G30595,G30598);
  and GNAME19780(G19780,G30592,G30595);
  or GNAME19781(G19781,G19780,G19779,G19778);
  xor GNAME19791(G19791,G19792,G30607);
  xor GNAME19792(G19792,G30601,G30604);
  and GNAME19793(G19793,G30601,G30607);
  and GNAME19794(G19794,G30604,G30607);
  and GNAME19795(G19795,G30601,G30604);
  or GNAME19796(G19796,G19795,G19794,G19793);
  xor GNAME19806(G19806,G19807,G30616);
  xor GNAME19807(G19807,G30610,G30613);
  and GNAME19808(G19808,G30610,G30616);
  and GNAME19809(G19809,G30613,G30616);
  and GNAME19810(G19810,G30610,G30613);
  or GNAME19811(G19811,G19810,G19809,G19808);
  xor GNAME19821(G19821,G19822,G30625);
  xor GNAME19822(G19822,G30619,G30622);
  and GNAME19823(G19823,G30619,G30625);
  and GNAME19824(G19824,G30622,G30625);
  and GNAME19825(G19825,G30619,G30622);
  or GNAME19826(G19826,G19825,G19824,G19823);
  xor GNAME19836(G19836,G19837,G30634);
  xor GNAME19837(G19837,G30628,G30631);
  and GNAME19838(G19838,G30628,G30634);
  and GNAME19839(G19839,G30631,G30634);
  and GNAME19840(G19840,G30628,G30631);
  or GNAME19841(G19841,G19840,G19839,G19838);
  xor GNAME19851(G19851,G19852,G30643);
  xor GNAME19852(G19852,G30637,G30640);
  and GNAME19853(G19853,G30637,G30643);
  and GNAME19854(G19854,G30640,G30643);
  and GNAME19855(G19855,G30637,G30640);
  or GNAME19856(G19856,G19855,G19854,G19853);
  xor GNAME19866(G19866,G19867,G30652);
  xor GNAME19867(G19867,G30646,G30649);
  and GNAME19868(G19868,G30646,G30652);
  and GNAME19869(G19869,G30649,G30652);
  and GNAME19870(G19870,G30646,G30649);
  or GNAME19871(G19871,G19870,G19869,G19868);
  xor GNAME19881(G19881,G19882,G30661);
  xor GNAME19882(G19882,G30655,G30658);
  and GNAME19883(G19883,G30655,G30661);
  and GNAME19884(G19884,G30658,G30661);
  and GNAME19885(G19885,G30655,G30658);
  or GNAME19886(G19886,G19885,G19884,G19883);
  xor GNAME19896(G19896,G19897,G30670);
  xor GNAME19897(G19897,G30664,G30667);
  and GNAME19898(G19898,G30664,G30670);
  and GNAME19899(G19899,G30667,G30670);
  and GNAME19900(G19900,G30664,G30667);
  or GNAME19901(G19901,G19900,G19899,G19898);
  xor GNAME19911(G19911,G19912,G30679);
  xor GNAME19912(G19912,G30673,G30676);
  and GNAME19913(G19913,G30673,G30679);
  and GNAME19914(G19914,G30676,G30679);
  and GNAME19915(G19915,G30673,G30676);
  or GNAME19916(G19916,G19915,G19914,G19913);
  xor GNAME19926(G19926,G19927,G30682);
  xor GNAME19927(G19927,G28972,G30685);
  and GNAME19928(G19928,G28972,G30682);
  and GNAME19929(G19929,G30685,G30682);
  and GNAME19930(G19930,G28972,G30685);
  or GNAME19931(G19931,G19930,G19929,G19928);
  xor GNAME19941(G19941,G19942,G30688);
  xor GNAME19942(G19942,G28973,G30691);
  and GNAME19943(G19943,G28973,G30688);
  and GNAME19944(G19944,G30691,G30688);
  and GNAME19945(G19945,G28973,G30691);
  or GNAME19946(G19946,G19945,G19944,G19943);
  xor GNAME19956(G19956,G19957,G30694);
  xor GNAME19957(G19957,G28974,G30697);
  and GNAME19958(G19958,G28974,G30694);
  and GNAME19959(G19959,G30697,G30694);
  and GNAME19960(G19960,G28974,G30697);
  or GNAME19961(G19961,G19960,G19959,G19958);
  xor GNAME19971(G19971,G19972,G30700);
  xor GNAME19972(G19972,G28975,G30703);
  and GNAME19973(G19973,G28975,G30700);
  and GNAME19974(G19974,G30703,G30700);
  and GNAME19975(G19975,G28975,G30703);
  or GNAME19976(G19976,G19975,G19974,G19973);
  xor GNAME19986(G19986,G19987,G30706);
  xor GNAME19987(G19987,G28976,G30709);
  and GNAME19988(G19988,G28976,G30706);
  and GNAME19989(G19989,G30709,G30706);
  and GNAME19990(G19990,G28976,G30709);
  or GNAME19991(G19991,G19990,G19989,G19988);
  xor GNAME20001(G20001,G20002,G30712);
  xor GNAME20002(G20002,G28977,G30715);
  and GNAME20003(G20003,G28977,G30712);
  and GNAME20004(G20004,G30715,G30712);
  and GNAME20005(G20005,G28977,G30715);
  or GNAME20006(G20006,G20005,G20004,G20003);
  xor GNAME20016(G20016,G20017,G30724);
  xor GNAME20017(G20017,G30718,G30721);
  and GNAME20018(G20018,G30718,G30724);
  and GNAME20019(G20019,G30721,G30724);
  and GNAME20020(G20020,G30718,G30721);
  or GNAME20021(G20021,G20020,G20019,G20018);
  xor GNAME20031(G20031,G20032,G30733);
  xor GNAME20032(G20032,G30727,G30730);
  and GNAME20033(G20033,G30727,G30733);
  and GNAME20034(G20034,G30730,G30733);
  and GNAME20035(G20035,G30727,G30730);
  or GNAME20036(G20036,G20035,G20034,G20033);
  xor GNAME20046(G20046,G20047,G30742);
  xor GNAME20047(G20047,G30736,G30739);
  and GNAME20048(G20048,G30736,G30742);
  and GNAME20049(G20049,G30739,G30742);
  and GNAME20050(G20050,G30736,G30739);
  or GNAME20051(G20051,G20050,G20049,G20048);
  xor GNAME20061(G20061,G20062,G30751);
  xor GNAME20062(G20062,G30745,G30748);
  and GNAME20063(G20063,G30745,G30751);
  and GNAME20064(G20064,G30748,G30751);
  and GNAME20065(G20065,G30745,G30748);
  or GNAME20066(G20066,G20065,G20064,G20063);
  xor GNAME20076(G20076,G20077,G30760);
  xor GNAME20077(G20077,G30754,G30757);
  and GNAME20078(G20078,G30754,G30760);
  and GNAME20079(G20079,G30757,G30760);
  and GNAME20080(G20080,G30754,G30757);
  or GNAME20081(G20081,G20080,G20079,G20078);
  xor GNAME20091(G20091,G20092,G30769);
  xor GNAME20092(G20092,G30763,G30766);
  and GNAME20093(G20093,G30763,G30769);
  and GNAME20094(G20094,G30766,G30769);
  and GNAME20095(G20095,G30763,G30766);
  or GNAME20096(G20096,G20095,G20094,G20093);
  xor GNAME20106(G20106,G20107,G30778);
  xor GNAME20107(G20107,G30772,G30775);
  and GNAME20108(G20108,G30772,G30778);
  and GNAME20109(G20109,G30775,G30778);
  and GNAME20110(G20110,G30772,G30775);
  or GNAME20111(G20111,G20110,G20109,G20108);
  xor GNAME20121(G20121,G20122,G30787);
  xor GNAME20122(G20122,G30781,G30784);
  and GNAME20123(G20123,G30781,G30787);
  and GNAME20124(G20124,G30784,G30787);
  and GNAME20125(G20125,G30781,G30784);
  or GNAME20126(G20126,G20125,G20124,G20123);
  xor GNAME20136(G20136,G20137,G30796);
  xor GNAME20137(G20137,G30790,G30793);
  and GNAME20138(G20138,G30790,G30796);
  and GNAME20139(G20139,G30793,G30796);
  and GNAME20140(G20140,G30790,G30793);
  or GNAME20141(G20141,G20140,G20139,G20138);
  xor GNAME20151(G20151,G20152,G30805);
  xor GNAME20152(G20152,G30799,G30802);
  and GNAME20153(G20153,G30799,G30805);
  and GNAME20154(G20154,G30802,G30805);
  and GNAME20155(G20155,G30799,G30802);
  or GNAME20156(G20156,G20155,G20154,G20153);
  xor GNAME20166(G20166,G20167,G30814);
  xor GNAME20167(G20167,G30808,G30811);
  and GNAME20168(G20168,G30808,G30814);
  and GNAME20169(G20169,G30811,G30814);
  and GNAME20170(G20170,G30808,G30811);
  or GNAME20171(G20171,G20170,G20169,G20168);
  xor GNAME20181(G20181,G20182,G30823);
  xor GNAME20182(G20182,G30817,G30820);
  and GNAME20183(G20183,G30817,G30823);
  and GNAME20184(G20184,G30820,G30823);
  and GNAME20185(G20185,G30817,G30820);
  or GNAME20186(G20186,G20185,G20184,G20183);
  xor GNAME20196(G20196,G20197,G30826);
  xor GNAME20197(G20197,G28978,G30829);
  and GNAME20198(G20198,G28978,G30826);
  and GNAME20199(G20199,G30829,G30826);
  and GNAME20200(G20200,G28978,G30829);
  or GNAME20201(G20201,G20200,G20199,G20198);
  xor GNAME20211(G20211,G20212,G30832);
  xor GNAME20212(G20212,G28979,G30835);
  and GNAME20213(G20213,G28979,G30832);
  and GNAME20214(G20214,G30835,G30832);
  and GNAME20215(G20215,G28979,G30835);
  or GNAME20216(G20216,G20215,G20214,G20213);
  xor GNAME20226(G20226,G20227,G30838);
  xor GNAME20227(G20227,G28980,G30841);
  and GNAME20228(G20228,G28980,G30838);
  and GNAME20229(G20229,G30841,G30838);
  and GNAME20230(G20230,G28980,G30841);
  or GNAME20231(G20231,G20230,G20229,G20228);
  xor GNAME20241(G20241,G20242,G30844);
  xor GNAME20242(G20242,G28981,G30847);
  and GNAME20243(G20243,G28981,G30844);
  and GNAME20244(G20244,G30847,G30844);
  and GNAME20245(G20245,G28981,G30847);
  or GNAME20246(G20246,G20245,G20244,G20243);
  xor GNAME20256(G20256,G20257,G30850);
  xor GNAME20257(G20257,G28982,G30853);
  and GNAME20258(G20258,G28982,G30850);
  and GNAME20259(G20259,G30853,G30850);
  and GNAME20260(G20260,G28982,G30853);
  or GNAME20261(G20261,G20260,G20259,G20258);
  xor GNAME20271(G20271,G20272,G30856);
  xor GNAME20272(G20272,G28983,G30859);
  and GNAME20273(G20273,G28983,G30856);
  and GNAME20274(G20274,G30859,G30856);
  and GNAME20275(G20275,G28983,G30859);
  or GNAME20276(G20276,G20275,G20274,G20273);
  xor GNAME20286(G20286,G20287,G30868);
  xor GNAME20287(G20287,G30862,G30865);
  and GNAME20288(G20288,G30862,G30868);
  and GNAME20289(G20289,G30865,G30868);
  and GNAME20290(G20290,G30862,G30865);
  or GNAME20291(G20291,G20290,G20289,G20288);
  xor GNAME20301(G20301,G20302,G30877);
  xor GNAME20302(G20302,G30871,G30874);
  and GNAME20303(G20303,G30871,G30877);
  and GNAME20304(G20304,G30874,G30877);
  and GNAME20305(G20305,G30871,G30874);
  or GNAME20306(G20306,G20305,G20304,G20303);
  xor GNAME20316(G20316,G20317,G30886);
  xor GNAME20317(G20317,G30880,G30883);
  and GNAME20318(G20318,G30880,G30886);
  and GNAME20319(G20319,G30883,G30886);
  and GNAME20320(G20320,G30880,G30883);
  or GNAME20321(G20321,G20320,G20319,G20318);
  xor GNAME20331(G20331,G20332,G30895);
  xor GNAME20332(G20332,G30889,G30892);
  and GNAME20333(G20333,G30889,G30895);
  and GNAME20334(G20334,G30892,G30895);
  and GNAME20335(G20335,G30889,G30892);
  or GNAME20336(G20336,G20335,G20334,G20333);
  xor GNAME20346(G20346,G20347,G30904);
  xor GNAME20347(G20347,G30898,G30901);
  and GNAME20348(G20348,G30898,G30904);
  and GNAME20349(G20349,G30901,G30904);
  and GNAME20350(G20350,G30898,G30901);
  or GNAME20351(G20351,G20350,G20349,G20348);
  xor GNAME20361(G20361,G20362,G30913);
  xor GNAME20362(G20362,G30907,G30910);
  and GNAME20363(G20363,G30907,G30913);
  and GNAME20364(G20364,G30910,G30913);
  and GNAME20365(G20365,G30907,G30910);
  or GNAME20366(G20366,G20365,G20364,G20363);
  xor GNAME20376(G20376,G20377,G20441);
  xor GNAME20377(G20377,G17546,G20621);
  and GNAME20378(G20378,G17546,G20441);
  and GNAME20379(G20379,G20621,G20441);
  and GNAME20380(G20380,G17546,G20621);
  or GNAME20381(G20381,G20380,G20379,G20378);
  xor GNAME20391(G20391,G20392,G20486);
  xor GNAME20392(G20392,G17561,G20666);
  and GNAME20393(G20393,G17561,G20486);
  and GNAME20394(G20394,G20666,G20486);
  and GNAME20395(G20395,G17561,G20666);
  or GNAME20396(G20396,G20395,G20394,G20393);
  xor GNAME20406(G20406,G20407,G20501);
  xor GNAME20407(G20407,G17576,G20681);
  and GNAME20408(G20408,G17576,G20501);
  and GNAME20409(G20409,G20681,G20501);
  and GNAME20410(G20410,G17576,G20681);
  or GNAME20411(G20411,G20410,G20409,G20408);
  xor GNAME20421(G20421,G20422,G30922);
  xor GNAME20422(G20422,G30916,G30919);
  and GNAME20423(G20423,G30916,G30922);
  and GNAME20424(G20424,G30919,G30922);
  and GNAME20425(G20425,G30916,G30919);
  or GNAME20426(G20426,G20425,G20424,G20423);
  xor GNAME20436(G20436,G20437,G30931);
  xor GNAME20437(G20437,G30925,G30928);
  and GNAME20438(G20438,G30925,G30931);
  and GNAME20439(G20439,G30928,G30931);
  and GNAME20440(G20440,G30925,G30928);
  or GNAME20441(G20441,G20440,G20439,G20438);
  xor GNAME20451(G20451,G20452,G30940);
  xor GNAME20452(G20452,G30934,G30937);
  and GNAME20453(G20453,G30934,G30940);
  and GNAME20454(G20454,G30937,G30940);
  and GNAME20455(G20455,G30934,G30937);
  or GNAME20456(G20456,G20455,G20454,G20453);
  xor GNAME20466(G20466,G20467,G30949);
  xor GNAME20467(G20467,G30943,G30946);
  and GNAME20468(G20468,G30943,G30949);
  and GNAME20469(G20469,G30946,G30949);
  and GNAME20470(G20470,G30943,G30946);
  or GNAME20471(G20471,G20470,G20469,G20468);
  xor GNAME20481(G20481,G20482,G30958);
  xor GNAME20482(G20482,G30952,G30955);
  and GNAME20483(G20483,G30952,G30958);
  and GNAME20484(G20484,G30955,G30958);
  and GNAME20485(G20485,G30952,G30955);
  or GNAME20486(G20486,G20485,G20484,G20483);
  xor GNAME20496(G20496,G20497,G30967);
  xor GNAME20497(G20497,G30961,G30964);
  and GNAME20498(G20498,G30961,G30967);
  and GNAME20499(G20499,G30964,G30967);
  and GNAME20500(G20500,G30961,G30964);
  or GNAME20501(G20501,G20500,G20499,G20498);
  xor GNAME20511(G20511,G20512,G20616);
  xor GNAME20512(G20512,G17541,G20436);
  and GNAME20513(G20513,G17541,G20616);
  and GNAME20514(G20514,G20436,G20616);
  and GNAME20515(G20515,G17541,G20436);
  or GNAME20516(G20516,G20515,G20514,G20513);
  xor GNAME20526(G20526,G20527,G20661);
  xor GNAME20527(G20527,G17556,G20481);
  and GNAME20528(G20528,G17556,G20661);
  and GNAME20529(G20529,G20481,G20661);
  and GNAME20530(G20530,G17556,G20481);
  or GNAME20531(G20531,G20530,G20529,G20528);
  xor GNAME20541(G20541,G20542,G20676);
  xor GNAME20542(G20542,G17571,G20496);
  and GNAME20543(G20543,G17571,G20676);
  and GNAME20544(G20544,G20496,G20676);
  and GNAME20545(G20545,G17571,G20496);
  or GNAME20546(G20546,G20545,G20544,G20543);
  xor GNAME20556(G20556,G20557,G30970);
  xor GNAME20557(G20557,G28984,G30973);
  and GNAME20558(G20558,G28984,G30970);
  and GNAME20559(G20559,G30973,G30970);
  and GNAME20560(G20560,G28984,G30973);
  or GNAME20561(G20561,G20560,G20559,G20558);
  xor GNAME20571(G20571,G20572,G30976);
  xor GNAME20572(G20572,G28985,G30979);
  and GNAME20573(G20573,G28985,G30976);
  and GNAME20574(G20574,G30979,G30976);
  and GNAME20575(G20575,G28985,G30979);
  or GNAME20576(G20576,G20575,G20574,G20573);
  xor GNAME20586(G20586,G20587,G30982);
  xor GNAME20587(G20587,G28986,G30985);
  and GNAME20588(G20588,G28986,G30982);
  and GNAME20589(G20589,G30985,G30982);
  and GNAME20590(G20590,G28986,G30985);
  or GNAME20591(G20591,G20590,G20589,G20588);
  xor GNAME20601(G20601,G20602,G30994);
  xor GNAME20602(G20602,G30988,G30991);
  and GNAME20603(G20603,G30988,G30994);
  and GNAME20604(G20604,G30991,G30994);
  and GNAME20605(G20605,G30988,G30991);
  or GNAME20606(G20606,G20605,G20604,G20603);
  xor GNAME20616(G20616,G20617,G31003);
  xor GNAME20617(G20617,G30997,G31000);
  and GNAME20618(G20618,G30997,G31003);
  and GNAME20619(G20619,G31000,G31003);
  and GNAME20620(G20620,G30997,G31000);
  or GNAME20621(G20621,G20620,G20619,G20618);
  xor GNAME20631(G20631,G20632,G31012);
  xor GNAME20632(G20632,G31006,G31009);
  and GNAME20633(G20633,G31006,G31012);
  and GNAME20634(G20634,G31009,G31012);
  and GNAME20635(G20635,G31006,G31009);
  or GNAME20636(G20636,G20635,G20634,G20633);
  xor GNAME20646(G20646,G20647,G31021);
  xor GNAME20647(G20647,G31015,G31018);
  and GNAME20648(G20648,G31015,G31021);
  and GNAME20649(G20649,G31018,G31021);
  and GNAME20650(G20650,G31015,G31018);
  or GNAME20651(G20651,G20650,G20649,G20648);
  xor GNAME20661(G20661,G20662,G31030);
  xor GNAME20662(G20662,G31024,G31027);
  and GNAME20663(G20663,G31024,G31030);
  and GNAME20664(G20664,G31027,G31030);
  and GNAME20665(G20665,G31024,G31027);
  or GNAME20666(G20666,G20665,G20664,G20663);
  xor GNAME20676(G20676,G20677,G31039);
  xor GNAME20677(G20677,G31033,G31036);
  and GNAME20678(G20678,G31033,G31039);
  and GNAME20679(G20679,G31036,G31039);
  and GNAME20680(G20680,G31033,G31036);
  or GNAME20681(G20681,G20680,G20679,G20678);
  xor GNAME20691(G20691,G20692,G31048);
  xor GNAME20692(G20692,G31042,G31045);
  and GNAME20693(G20693,G31042,G31048);
  and GNAME20694(G20694,G31045,G31048);
  and GNAME20695(G20695,G31042,G31045);
  or GNAME20696(G20696,G20695,G20694,G20693);
  xor GNAME20706(G20706,G20707,G31057);
  xor GNAME20707(G20707,G31051,G31054);
  and GNAME20708(G20708,G31051,G31057);
  and GNAME20709(G20709,G31054,G31057);
  and GNAME20710(G20710,G31051,G31054);
  or GNAME20711(G20711,G20710,G20709,G20708);
  xor GNAME20721(G20721,G20722,G31066);
  xor GNAME20722(G20722,G31060,G31063);
  and GNAME20723(G20723,G31060,G31066);
  and GNAME20724(G20724,G31063,G31066);
  and GNAME20725(G20725,G31060,G31063);
  or GNAME20726(G20726,G20725,G20724,G20723);
  xor GNAME20736(G20736,G20737,G20696);
  xor GNAME20737(G20737,G28127,G20921);
  and GNAME20738(G20738,G28127,G20696);
  and GNAME20739(G20739,G20921,G20696);
  and GNAME20740(G20740,G28127,G20921);
  or GNAME20741(G20741,G20740,G20739,G20738);
  xor GNAME20751(G20751,G20752,G20711);
  xor GNAME20752(G20752,G28133,G20951);
  and GNAME20753(G20753,G28133,G20711);
  and GNAME20754(G20754,G20951,G20711);
  and GNAME20755(G20755,G28133,G20951);
  or GNAME20756(G20756,G20755,G20754,G20753);
  xor GNAME20766(G20766,G20767,G20726);
  xor GNAME20767(G20767,G28139,G20966);
  and GNAME20768(G20768,G28139,G20726);
  and GNAME20769(G20769,G20966,G20726);
  and GNAME20770(G20770,G28139,G20966);
  or GNAME20771(G20771,G20770,G20769,G20768);
  xor GNAME20781(G20781,G20782,G28109);
  xor GNAME20782(G20782,G31069,G31072);
  and GNAME20783(G20783,G31069,G28109);
  and GNAME20784(G20784,G31072,G28109);
  and GNAME20785(G20785,G31069,G31072);
  or GNAME20786(G20786,G20785,G20784,G20783);
  xor GNAME20796(G20796,G20797,G28115);
  xor GNAME20797(G20797,G31075,G31078);
  and GNAME20798(G20798,G31075,G28115);
  and GNAME20799(G20799,G31078,G28115);
  and GNAME20800(G20800,G31075,G31078);
  or GNAME20801(G20801,G20800,G20799,G20798);
  xor GNAME20811(G20811,G20812,G28121);
  xor GNAME20812(G20812,G31081,G31084);
  and GNAME20813(G20813,G31081,G28121);
  and GNAME20814(G20814,G31084,G28121);
  and GNAME20815(G20815,G31081,G31084);
  or GNAME20816(G20816,G20815,G20814,G20813);
  xor GNAME20826(G20826,G20827,G17591);
  xor GNAME20827(G20827,G31087,G28126);
  and GNAME20828(G20828,G31087,G17591);
  and GNAME20829(G20829,G28126,G17591);
  and GNAME20830(G20830,G31087,G28126);
  or GNAME20831(G20831,G20830,G20829,G20828);
  xor GNAME20841(G20841,G20842,G17606);
  xor GNAME20842(G20842,G31090,G28132);
  and GNAME20843(G20843,G31090,G17606);
  and GNAME20844(G20844,G28132,G17606);
  and GNAME20845(G20845,G31090,G28132);
  or GNAME20846(G20846,G20845,G20844,G20843);
  xor GNAME20856(G20856,G20857,G17621);
  xor GNAME20857(G20857,G31093,G28138);
  and GNAME20858(G20858,G31093,G17621);
  and GNAME20859(G20859,G28138,G17621);
  and GNAME20860(G20860,G31093,G28138);
  or GNAME20861(G20861,G20860,G20859,G20858);
  xor GNAME20871(G20871,G20872,G17586);
  xor GNAME20872(G20872,G21056,G21281);
  and GNAME20873(G20873,G21056,G17586);
  and GNAME20874(G20874,G21281,G17586);
  and GNAME20875(G20875,G21056,G21281);
  or GNAME20876(G20876,G20875,G20874,G20873);
  xor GNAME20886(G20886,G20887,G17601);
  xor GNAME20887(G20887,G21086,G21296);
  and GNAME20888(G20888,G21086,G17601);
  and GNAME20889(G20889,G21296,G17601);
  and GNAME20890(G20890,G21086,G21296);
  or GNAME20891(G20891,G20890,G20889,G20888);
  xor GNAME20901(G20901,G20902,G17616);
  xor GNAME20902(G20902,G21101,G21311);
  and GNAME20903(G20903,G21101,G17616);
  and GNAME20904(G20904,G21311,G17616);
  and GNAME20905(G20905,G21101,G21311);
  or GNAME20906(G20906,G20905,G20904,G20903);
  xor GNAME20916(G20916,G20917,G31099);
  xor GNAME20917(G20917,G31096,G31102);
  and GNAME20918(G20918,G31096,G31099);
  and GNAME20919(G20919,G31102,G31099);
  and GNAME20920(G20920,G31096,G31102);
  or GNAME20921(G20921,G20920,G20919,G20918);
  xor GNAME20931(G20931,G20932,G31111);
  xor GNAME20932(G20932,G31105,G31108);
  and GNAME20933(G20933,G31105,G31111);
  and GNAME20934(G20934,G31108,G31111);
  and GNAME20935(G20935,G31105,G31108);
  or GNAME20936(G20936,G20935,G20934,G20933);
  xor GNAME20946(G20946,G20947,G31117);
  xor GNAME20947(G20947,G31114,G31120);
  and GNAME20948(G20948,G31114,G31117);
  and GNAME20949(G20949,G31120,G31117);
  and GNAME20950(G20950,G31114,G31120);
  or GNAME20951(G20951,G20950,G20949,G20948);
  xor GNAME20961(G20961,G20962,G31126);
  xor GNAME20962(G20962,G31123,G31129);
  and GNAME20963(G20963,G31123,G31126);
  and GNAME20964(G20964,G31129,G31126);
  and GNAME20965(G20965,G31123,G31129);
  or GNAME20966(G20966,G20965,G20964,G20963);
  xor GNAME20976(G20976,G20977,G31138);
  xor GNAME20977(G20977,G31132,G31135);
  and GNAME20978(G20978,G31132,G31138);
  and GNAME20979(G20979,G31135,G31138);
  and GNAME20980(G20980,G31132,G31135);
  or GNAME20981(G20981,G20980,G20979,G20978);
  xor GNAME20991(G20991,G20992,G31147);
  xor GNAME20992(G20992,G31141,G31144);
  and GNAME20993(G20993,G31141,G31147);
  and GNAME20994(G20994,G31144,G31147);
  and GNAME20995(G20995,G31141,G31144);
  or GNAME20996(G20996,G20995,G20994,G20993);
  xor GNAME21006(G21006,G21007,G21206);
  xor GNAME21007(G21007,G17631,G21066);
  and GNAME21008(G21008,G17631,G21206);
  and GNAME21009(G21009,G21066,G21206);
  and GNAME21010(G21010,G17631,G21066);
  or GNAME21011(G21011,G21010,G21009,G21008);
  xor GNAME21021(G21021,G21022,G21251);
  xor GNAME21022(G21022,G17646,G21111);
  and GNAME21023(G21023,G17646,G21251);
  and GNAME21024(G21024,G21111,G21251);
  and GNAME21025(G21025,G17646,G21111);
  or GNAME21026(G21026,G21025,G21024,G21023);
  xor GNAME21036(G21036,G21037,G21266);
  xor GNAME21037(G21037,G17661,G21126);
  and GNAME21038(G21038,G17661,G21266);
  and GNAME21039(G21039,G21126,G21266);
  and GNAME21040(G21040,G17661,G21126);
  or GNAME21041(G21041,G21040,G21039,G21038);
  xor GNAME21051(G21051,G21052,G31156);
  xor GNAME21052(G21052,G31150,G31153);
  and GNAME21053(G21053,G31150,G31156);
  and GNAME21054(G21054,G31153,G31156);
  and GNAME21055(G21055,G31150,G31153);
  or GNAME21056(G21056,G21055,G21054,G21053);
  xor GNAME21066(G21066,G21067,G31165);
  xor GNAME21067(G21067,G31159,G31162);
  and GNAME21068(G21068,G31159,G31165);
  and GNAME21069(G21069,G31162,G31165);
  and GNAME21070(G21070,G31159,G31162);
  or GNAME21071(G21071,G21070,G21069,G21068);
  xor GNAME21081(G21081,G21082,G31174);
  xor GNAME21082(G21082,G31168,G31171);
  and GNAME21083(G21083,G31168,G31174);
  and GNAME21084(G21084,G31171,G31174);
  and GNAME21085(G21085,G31168,G31171);
  or GNAME21086(G21086,G21085,G21084,G21083);
  xor GNAME21096(G21096,G21097,G31183);
  xor GNAME21097(G21097,G31177,G31180);
  and GNAME21098(G21098,G31177,G31183);
  and GNAME21099(G21099,G31180,G31183);
  and GNAME21100(G21100,G31177,G31180);
  or GNAME21101(G21101,G21100,G21099,G21098);
  xor GNAME21111(G21111,G21112,G31192);
  xor GNAME21112(G21112,G31186,G31189);
  and GNAME21113(G21113,G31186,G31192);
  and GNAME21114(G21114,G31189,G31192);
  and GNAME21115(G21115,G31186,G31189);
  or GNAME21116(G21116,G21115,G21114,G21113);
  xor GNAME21126(G21126,G21127,G31201);
  xor GNAME21127(G21127,G31195,G31198);
  and GNAME21128(G21128,G31195,G31201);
  and GNAME21129(G21129,G31198,G31201);
  and GNAME21130(G21130,G31195,G31198);
  or GNAME21131(G21131,G21130,G21129,G21128);
  xor GNAME21141(G21141,G21142,G21071);
  xor GNAME21142(G21142,G28108,G17636);
  and GNAME21143(G21143,G28108,G21071);
  and GNAME21144(G21144,G17636,G21071);
  and GNAME21145(G21145,G28108,G17636);
  or GNAME21146(G21146,G21145,G21144,G21143);
  xor GNAME21156(G21156,G21157,G21116);
  xor GNAME21157(G21157,G28114,G17651);
  and GNAME21158(G21158,G28114,G21116);
  and GNAME21159(G21159,G17651,G21116);
  and GNAME21160(G21160,G28114,G17651);
  or GNAME21161(G21161,G21160,G21159,G21158);
  xor GNAME21171(G21171,G21172,G21131);
  xor GNAME21172(G21172,G28120,G17666);
  and GNAME21173(G21173,G28120,G21131);
  and GNAME21174(G21174,G17666,G21131);
  and GNAME21175(G21175,G28120,G17666);
  or GNAME21176(G21176,G21175,G21174,G21173);
  xor GNAME21186(G21186,G21187,G21326);
  xor GNAME21187(G21187,G31204,G28145);
  and GNAME21188(G21188,G31204,G21326);
  and GNAME21189(G21189,G28145,G21326);
  and GNAME21190(G21190,G31204,G28145);
  or GNAME21191(G21191,G21190,G21189,G21188);
  xor GNAME21201(G21201,G21202,G28144);
  xor GNAME21202(G21202,G31207,G31210);
  and GNAME21203(G21203,G31207,G28144);
  and GNAME21204(G21204,G31210,G28144);
  and GNAME21205(G21205,G31207,G31210);
  or GNAME21206(G21206,G21205,G21204,G21203);
  xor GNAME21216(G21216,G21217,G21341);
  xor GNAME21217(G21217,G31213,G28151);
  and GNAME21218(G21218,G31213,G21341);
  and GNAME21219(G21219,G28151,G21341);
  and GNAME21220(G21220,G31213,G28151);
  or GNAME21221(G21221,G21220,G21219,G21218);
  xor GNAME21231(G21231,G21232,G21356);
  xor GNAME21232(G21232,G31216,G28157);
  and GNAME21233(G21233,G31216,G21356);
  and GNAME21234(G21234,G28157,G21356);
  and GNAME21235(G21235,G31216,G28157);
  or GNAME21236(G21236,G21235,G21234,G21233);
  xor GNAME21246(G21246,G21247,G28150);
  xor GNAME21247(G21247,G31219,G31222);
  and GNAME21248(G21248,G31219,G28150);
  and GNAME21249(G21249,G31222,G28150);
  and GNAME21250(G21250,G31219,G31222);
  or GNAME21251(G21251,G21250,G21249,G21248);
  xor GNAME21261(G21261,G21262,G28156);
  xor GNAME21262(G21262,G31225,G31228);
  and GNAME21263(G21263,G31225,G28156);
  and GNAME21264(G21264,G31228,G28156);
  and GNAME21265(G21265,G31225,G31228);
  or GNAME21266(G21266,G21265,G21264,G21263);
  xor GNAME21276(G21276,G21277,G31234);
  xor GNAME21277(G21277,G31231,G31237);
  and GNAME21278(G21278,G31231,G31234);
  and GNAME21279(G21279,G31237,G31234);
  and GNAME21280(G21280,G31231,G31237);
  or GNAME21281(G21281,G21280,G21279,G21278);
  xor GNAME21291(G21291,G21292,G31243);
  xor GNAME21292(G21292,G31240,G31246);
  and GNAME21293(G21293,G31240,G31243);
  and GNAME21294(G21294,G31246,G31243);
  and GNAME21295(G21295,G31240,G31246);
  or GNAME21296(G21296,G21295,G21294,G21293);
  xor GNAME21306(G21306,G21307,G31252);
  xor GNAME21307(G21307,G31249,G31255);
  and GNAME21308(G21308,G31249,G31252);
  and GNAME21309(G21309,G31255,G31252);
  and GNAME21310(G21310,G31249,G31255);
  or GNAME21311(G21311,G21310,G21309,G21308);
  xor GNAME21321(G21321,G21322,G31261);
  xor GNAME21322(G21322,G31258,G31264);
  and GNAME21323(G21323,G31258,G31261);
  and GNAME21324(G21324,G31264,G31261);
  and GNAME21325(G21325,G31258,G31264);
  or GNAME21326(G21326,G21325,G21324,G21323);
  xor GNAME21336(G21336,G21337,G31270);
  xor GNAME21337(G21337,G31267,G31273);
  and GNAME21338(G21338,G31267,G31270);
  and GNAME21339(G21339,G31273,G31270);
  and GNAME21340(G21340,G31267,G31273);
  or GNAME21341(G21341,G21340,G21339,G21338);
  xor GNAME21351(G21351,G21352,G31279);
  xor GNAME21352(G21352,G31276,G31282);
  and GNAME21353(G21353,G31276,G31279);
  and GNAME21354(G21354,G31282,G31279);
  and GNAME21355(G21355,G31276,G31282);
  or GNAME21356(G21356,G21355,G21354,G21353);
  xor GNAME21366(G21366,G21367,G21321);
  xor GNAME21367(G21367,G17681,G21506);
  and GNAME21368(G21368,G17681,G21321);
  and GNAME21369(G21369,G21506,G21321);
  and GNAME21370(G21370,G17681,G21506);
  or GNAME21371(G21371,G21370,G21369,G21368);
  xor GNAME21381(G21381,G21382,G17676);
  xor GNAME21382(G21382,G28163,G21461);
  and GNAME21383(G21383,G28163,G17676);
  and GNAME21384(G21384,G21461,G17676);
  and GNAME21385(G21385,G28163,G21461);
  or GNAME21386(G21386,G21385,G21384,G21383);
  xor GNAME21396(G21396,G21397,G21336);
  xor GNAME21397(G21397,G17696,G21521);
  and GNAME21398(G21398,G17696,G21336);
  and GNAME21399(G21399,G21521,G21336);
  and GNAME21400(G21400,G17696,G21521);
  or GNAME21401(G21401,G21400,G21399,G21398);
  xor GNAME21411(G21411,G21412,G21351);
  xor GNAME21412(G21412,G17711,G21536);
  and GNAME21413(G21413,G17711,G21351);
  and GNAME21414(G21414,G21536,G21351);
  and GNAME21415(G21415,G17711,G21536);
  or GNAME21416(G21416,G21415,G21414,G21413);
  xor GNAME21426(G21426,G21427,G17691);
  xor GNAME21427(G21427,G28169,G21476);
  and GNAME21428(G21428,G28169,G17691);
  and GNAME21429(G21429,G21476,G17691);
  and GNAME21430(G21430,G28169,G21476);
  or GNAME21431(G21431,G21430,G21429,G21428);
  xor GNAME21441(G21441,G21442,G17706);
  xor GNAME21442(G21442,G28175,G21491);
  and GNAME21443(G21443,G28175,G17706);
  and GNAME21444(G21444,G21491,G17706);
  and GNAME21445(G21445,G28175,G21491);
  or GNAME21446(G21446,G21445,G21444,G21443);
  xor GNAME21456(G21456,G21457,G31288);
  xor GNAME21457(G21457,G31285,G31291);
  and GNAME21458(G21458,G31285,G31288);
  and GNAME21459(G21459,G31291,G31288);
  and GNAME21460(G21460,G31285,G31291);
  or GNAME21461(G21461,G21460,G21459,G21458);
  xor GNAME21471(G21471,G21472,G31297);
  xor GNAME21472(G21472,G31294,G31300);
  and GNAME21473(G21473,G31294,G31297);
  and GNAME21474(G21474,G31300,G31297);
  and GNAME21475(G21475,G31294,G31300);
  or GNAME21476(G21476,G21475,G21474,G21473);
  xor GNAME21486(G21486,G21487,G31306);
  xor GNAME21487(G21487,G31303,G31309);
  and GNAME21488(G21488,G31303,G31306);
  and GNAME21489(G21489,G31309,G31306);
  and GNAME21490(G21490,G31303,G31309);
  or GNAME21491(G21491,G21490,G21489,G21488);
  xor GNAME21501(G21501,G21502,G31318);
  xor GNAME21502(G21502,G31312,G31315);
  and GNAME21503(G21503,G31312,G31318);
  and GNAME21504(G21504,G31315,G31318);
  and GNAME21505(G21505,G31312,G31315);
  or GNAME21506(G21506,G21505,G21504,G21503);
  xor GNAME21516(G21516,G21517,G31327);
  xor GNAME21517(G21517,G31321,G31324);
  and GNAME21518(G21518,G31321,G31327);
  and GNAME21519(G21519,G31324,G31327);
  and GNAME21520(G21520,G31321,G31324);
  or GNAME21521(G21521,G21520,G21519,G21518);
  xor GNAME21531(G21531,G21532,G31336);
  xor GNAME21532(G21532,G31330,G31333);
  and GNAME21533(G21533,G31330,G31336);
  and GNAME21534(G21534,G31333,G31336);
  and GNAME21535(G21535,G31330,G31333);
  or GNAME21536(G21536,G21535,G21534,G21533);
  xor GNAME21546(G21546,G21547,G31342);
  xor GNAME21547(G21547,G31339,G31345);
  and GNAME21548(G21548,G31339,G31342);
  and GNAME21549(G21549,G31345,G31342);
  and GNAME21550(G21550,G31339,G31345);
  or GNAME21551(G21551,G21550,G21549,G21548);
  xor GNAME21561(G21561,G21562,G31351);
  xor GNAME21562(G21562,G31348,G31354);
  and GNAME21563(G21563,G31348,G31351);
  and GNAME21564(G21564,G31354,G31351);
  and GNAME21565(G21565,G31348,G31354);
  or GNAME21566(G21566,G21565,G21564,G21563);
  xor GNAME21576(G21576,G21577,G31360);
  xor GNAME21577(G21577,G31357,G31363);
  and GNAME21578(G21578,G31357,G31360);
  and GNAME21579(G21579,G31363,G31360);
  and GNAME21580(G21580,G31357,G31363);
  or GNAME21581(G21581,G21580,G21579,G21578);
  xor GNAME21591(G21591,G21592,G28181);
  xor GNAME21592(G21592,G31366,G31369);
  and GNAME21593(G21593,G31366,G28181);
  and GNAME21594(G21594,G31369,G28181);
  and GNAME21595(G21595,G31366,G31369);
  or GNAME21596(G21596,G21595,G21594,G21593);
  xor GNAME21606(G21606,G21607,G28187);
  xor GNAME21607(G21607,G31372,G31375);
  and GNAME21608(G21608,G31372,G28187);
  and GNAME21609(G21609,G31375,G28187);
  and GNAME21610(G21610,G31372,G31375);
  or GNAME21611(G21611,G21610,G21609,G21608);
  xor GNAME21621(G21621,G21622,G28193);
  xor GNAME21622(G21622,G31378,G31381);
  and GNAME21623(G21623,G31378,G28193);
  and GNAME21624(G21624,G31381,G28193);
  and GNAME21625(G21625,G31378,G31381);
  or GNAME21626(G21626,G21625,G21624,G21623);
  xor GNAME21636(G21636,G21637,G17726);
  xor GNAME21637(G21637,G31384,G28162);
  and GNAME21638(G21638,G31384,G17726);
  and GNAME21639(G21639,G28162,G17726);
  and GNAME21640(G21640,G31384,G28162);
  or GNAME21641(G21641,G21640,G21639,G21638);
  xor GNAME21651(G21651,G21652,G17741);
  xor GNAME21652(G21652,G31387,G28168);
  and GNAME21653(G21653,G31387,G17741);
  and GNAME21654(G21654,G28168,G17741);
  and GNAME21655(G21655,G31387,G28168);
  or GNAME21656(G21656,G21655,G21654,G21653);
  xor GNAME21666(G21666,G21667,G17756);
  xor GNAME21667(G21667,G31390,G28174);
  and GNAME21668(G21668,G31390,G17756);
  and GNAME21669(G21669,G28174,G17756);
  and GNAME21670(G21670,G31390,G28174);
  or GNAME21671(G21671,G21670,G21669,G21668);
  xor GNAME21681(G21681,G21682,G21546);
  xor GNAME21682(G21682,G28180,G17771);
  and GNAME21683(G21683,G28180,G21546);
  and GNAME21684(G21684,G17771,G21546);
  and GNAME21685(G21685,G28180,G17771);
  or GNAME21686(G21686,G21685,G21684,G21683);
  xor GNAME21696(G21696,G21697,G21591);
  xor GNAME21697(G21697,G21551,G17721);
  and GNAME21698(G21698,G21551,G21591);
  and GNAME21699(G21699,G17721,G21591);
  and GNAME21700(G21700,G21551,G17721);
  or GNAME21701(G21701,G21700,G21699,G21698);
  xor GNAME21711(G21711,G21712,G21606);
  xor GNAME21712(G21712,G21566,G17736);
  and GNAME21713(G21713,G21566,G21606);
  and GNAME21714(G21714,G17736,G21606);
  and GNAME21715(G21715,G21566,G17736);
  or GNAME21716(G21716,G21715,G21714,G21713);
  xor GNAME21726(G21726,G21727,G21621);
  xor GNAME21727(G21727,G21581,G17751);
  and GNAME21728(G21728,G21581,G21621);
  and GNAME21729(G21729,G17751,G21621);
  and GNAME21730(G21730,G21581,G17751);
  or GNAME21731(G21731,G21730,G21729,G21728);
  xor GNAME21741(G21741,G21742,G21561);
  xor GNAME21742(G21742,G28186,G17786);
  and GNAME21743(G21743,G28186,G21561);
  and GNAME21744(G21744,G17786,G21561);
  and GNAME21745(G21745,G28186,G17786);
  or GNAME21746(G21746,G21745,G21744,G21743);
  xor GNAME21756(G21756,G21757,G21576);
  xor GNAME21757(G21757,G28192,G17801);
  and GNAME21758(G21758,G28192,G21576);
  and GNAME21759(G21759,G17801,G21576);
  and GNAME21760(G21760,G28192,G17801);
  or GNAME21761(G21761,G21760,G21759,G21758);
  xor GNAME21771(G21771,G21772,G17766);
  xor GNAME21772(G21772,G31393,G28217);
  and GNAME21773(G21773,G31393,G17766);
  and GNAME21774(G21774,G28217,G17766);
  and GNAME21775(G21775,G31393,G28217);
  or GNAME21776(G21776,G21775,G21774,G21773);
  xor GNAME21786(G21786,G21787,G28879);
  xor GNAME21787(G21787,G21776,G21681);
  and GNAME21788(G21788,G21776,G28879);
  and GNAME21789(G21789,G21681,G28879);
  and GNAME21790(G21790,G21776,G21681);
  or GNAME21791(G21791,G21790,G21789,G21788);
  xor GNAME21801(G21801,G21802,G17781);
  xor GNAME21802(G21802,G31396,G28223);
  and GNAME21803(G21803,G31396,G17781);
  and GNAME21804(G21804,G28223,G17781);
  and GNAME21805(G21805,G31396,G28223);
  or GNAME21806(G21806,G21805,G21804,G21803);
  xor GNAME21816(G21816,G21817,G28899);
  xor GNAME21817(G21817,G21806,G21741);
  and GNAME21818(G21818,G21806,G28899);
  and GNAME21819(G21819,G21741,G28899);
  and GNAME21820(G21820,G21806,G21741);
  or GNAME21821(G21821,G21820,G21819,G21818);
  xor GNAME21831(G21831,G21832,G17796);
  xor GNAME21832(G21832,G31399,G28229);
  and GNAME21833(G21833,G31399,G17796);
  and GNAME21834(G21834,G28229,G17796);
  and GNAME21835(G21835,G31399,G28229);
  or GNAME21836(G21836,G21835,G21834,G21833);
  xor GNAME21846(G21846,G21847,G28919);
  xor GNAME21847(G21847,G21836,G21756);
  and GNAME21848(G21848,G21836,G28919);
  and GNAME21849(G21849,G21756,G28919);
  and GNAME21850(G21850,G21836,G21756);
  or GNAME21851(G21851,G21850,G21849,G21848);
  xor GNAME21861(G21861,G21862,G18311);
  xor GNAME21862(G21862,G18216,G18171);
  and GNAME21863(G21863,G18216,G18311);
  and GNAME21864(G21864,G18171,G18311);
  and GNAME21865(G21865,G18216,G18171);
  or GNAME21866(G21866,G21865,G21864,G21863);
  xor GNAME21876(G21876,G21877,G18326);
  xor GNAME21877(G21877,G18231,G18186);
  and GNAME21878(G21878,G18231,G18326);
  and GNAME21879(G21879,G18186,G18326);
  and GNAME21880(G21880,G18231,G18186);
  or GNAME21881(G21881,G21880,G21879,G21878);
  xor GNAME21891(G21891,G21892,G18341);
  xor GNAME21892(G21892,G18246,G18201);
  and GNAME21893(G21893,G18246,G18341);
  and GNAME21894(G21894,G18201,G18341);
  and GNAME21895(G21895,G18246,G18201);
  or GNAME21896(G21896,G21895,G21894,G21893);
  xor GNAME21906(G21906,G21907,G21956);
  xor GNAME21907(G21907,G18401,G18306);
  and GNAME21908(G21908,G18401,G21956);
  and GNAME21909(G21909,G18306,G21956);
  and GNAME21910(G21910,G18401,G18306);
  or GNAME21911(G21911,G21910,G21909,G21908);
  xor GNAME21921(G21921,G21922,G21971);
  xor GNAME21922(G21922,G18416,G18321);
  and GNAME21923(G21923,G18416,G21971);
  and GNAME21924(G21924,G18321,G21971);
  and GNAME21925(G21925,G18416,G18321);
  or GNAME21926(G21926,G21925,G21924,G21923);
  xor GNAME21936(G21936,G21937,G21986);
  xor GNAME21937(G21937,G18431,G18336);
  and GNAME21938(G21938,G18431,G21986);
  and GNAME21939(G21939,G18336,G21986);
  and GNAME21940(G21940,G18431,G18336);
  or GNAME21941(G21941,G21940,G21939,G21938);
  xor GNAME21951(G21951,G21952,G18581);
  xor GNAME21952(G21952,G18671,G18351);
  and GNAME21953(G21953,G18671,G18581);
  and GNAME21954(G21954,G18351,G18581);
  and GNAME21955(G21955,G18671,G18351);
  or GNAME21956(G21956,G21955,G21954,G21953);
  xor GNAME21966(G21966,G21967,G18596);
  xor GNAME21967(G21967,G18686,G18366);
  and GNAME21968(G21968,G18686,G18596);
  and GNAME21969(G21969,G18366,G18596);
  and GNAME21970(G21970,G18686,G18366);
  or GNAME21971(G21971,G21970,G21969,G21968);
  xor GNAME21981(G21981,G21982,G18611);
  xor GNAME21982(G21982,G18701,G18381);
  and GNAME21983(G21983,G18701,G18611);
  and GNAME21984(G21984,G18381,G18611);
  and GNAME21985(G21985,G18701,G18381);
  or GNAME21986(G21986,G21985,G21984,G21983);
  xor GNAME21996(G21996,G21997,G21951);
  xor GNAME21997(G21997,G18396,G18446);
  and GNAME21998(G21998,G18396,G21951);
  and GNAME21999(G21999,G18446,G21951);
  and GNAME22000(G22000,G18396,G18446);
  or GNAME22001(G22001,G22000,G21999,G21998);
  xor GNAME22011(G22011,G22012,G18441);
  xor GNAME22012(G22012,G18576,G22091);
  and GNAME22013(G22013,G18576,G18441);
  and GNAME22014(G22014,G22091,G18441);
  and GNAME22015(G22015,G18576,G22091);
  or GNAME22016(G22016,G22015,G22014,G22013);
  xor GNAME22026(G22026,G22027,G21966);
  xor GNAME22027(G22027,G18411,G18461);
  and GNAME22028(G22028,G18411,G21966);
  and GNAME22029(G22029,G18461,G21966);
  and GNAME22030(G22030,G18411,G18461);
  or GNAME22031(G22031,G22030,G22029,G22028);
  xor GNAME22041(G22041,G22042,G21981);
  xor GNAME22042(G22042,G18426,G18476);
  and GNAME22043(G22043,G18426,G21981);
  and GNAME22044(G22044,G18476,G21981);
  and GNAME22045(G22045,G18426,G18476);
  or GNAME22046(G22046,G22045,G22044,G22043);
  xor GNAME22056(G22056,G22057,G18456);
  xor GNAME22057(G22057,G18591,G22121);
  and GNAME22058(G22058,G18591,G18456);
  and GNAME22059(G22059,G22121,G18456);
  and GNAME22060(G22060,G18591,G22121);
  or GNAME22061(G22061,G22060,G22059,G22058);
  xor GNAME22071(G22071,G22072,G18471);
  xor GNAME22072(G22072,G18606,G22151);
  and GNAME22073(G22073,G18606,G18471);
  and GNAME22074(G22074,G22151,G18471);
  and GNAME22075(G22075,G18606,G22151);
  or GNAME22076(G22076,G22075,G22074,G22073);
  xor GNAME22086(G22086,G22087,G18851);
  xor GNAME22087(G22087,G18621,G18761);
  and GNAME22088(G22088,G18621,G18851);
  and GNAME22089(G22089,G18761,G18851);
  and GNAME22090(G22090,G18621,G18761);
  or GNAME22091(G22091,G22090,G22089,G22088);
  xor GNAME22101(G22101,G22102,G22271);
  xor GNAME22102(G22102,G18986,G18756);
  and GNAME22103(G22103,G18986,G22271);
  and GNAME22104(G22104,G18756,G22271);
  and GNAME22105(G22105,G18986,G18756);
  or GNAME22106(G22106,G22105,G22104,G22103);
  xor GNAME22116(G22116,G22117,G18866);
  xor GNAME22117(G22117,G18636,G18776);
  and GNAME22118(G22118,G18636,G18866);
  and GNAME22119(G22119,G18776,G18866);
  and GNAME22120(G22120,G18636,G18776);
  or GNAME22121(G22121,G22120,G22119,G22118);
  xor GNAME22131(G22131,G22132,G22286);
  xor GNAME22132(G22132,G19016,G18771);
  and GNAME22133(G22133,G19016,G22286);
  and GNAME22134(G22134,G18771,G22286);
  and GNAME22135(G22135,G19016,G18771);
  or GNAME22136(G22136,G22135,G22134,G22133);
  xor GNAME22146(G22146,G22147,G18881);
  xor GNAME22147(G22147,G18651,G18791);
  and GNAME22148(G22148,G18651,G18881);
  and GNAME22149(G22149,G18791,G18881);
  and GNAME22150(G22150,G18651,G18791);
  or GNAME22151(G22151,G22150,G22149,G22148);
  xor GNAME22161(G22161,G22162,G22301);
  xor GNAME22162(G22162,G19031,G18786);
  and GNAME22163(G22163,G19031,G22301);
  and GNAME22164(G22164,G18786,G22301);
  and GNAME22165(G22165,G19031,G18786);
  or GNAME22166(G22166,G22165,G22164,G22163);
  xor GNAME22176(G22176,G22177,G22086);
  xor GNAME22177(G22177,G18531,G22106);
  and GNAME22178(G22178,G18531,G22086);
  and GNAME22179(G22179,G22106,G22086);
  and GNAME22180(G22180,G18531,G22106);
  or GNAME22181(G22181,G22180,G22179,G22178);
  xor GNAME22191(G22191,G22192,G22101);
  xor GNAME22192(G22192,G18846,G22316);
  and GNAME22193(G22193,G18846,G22101);
  and GNAME22194(G22194,G22316,G22101);
  and GNAME22195(G22195,G18846,G22316);
  or GNAME22196(G22196,G22195,G22194,G22193);
  xor GNAME22206(G22206,G22207,G22116);
  xor GNAME22207(G22207,G18546,G22136);
  and GNAME22208(G22208,G18546,G22116);
  and GNAME22209(G22209,G22136,G22116);
  and GNAME22210(G22210,G18546,G22136);
  or GNAME22211(G22211,G22210,G22209,G22208);
  xor GNAME22221(G22221,G22222,G22146);
  xor GNAME22222(G22222,G18561,G22166);
  and GNAME22223(G22223,G18561,G22146);
  and GNAME22224(G22224,G22166,G22146);
  and GNAME22225(G22225,G18561,G22166);
  or GNAME22226(G22226,G22225,G22224,G22223);
  xor GNAME22236(G22236,G22237,G22131);
  xor GNAME22237(G22237,G18861,G22346);
  and GNAME22238(G22238,G18861,G22131);
  and GNAME22239(G22239,G22346,G22131);
  and GNAME22240(G22240,G18861,G22346);
  or GNAME22241(G22241,G22240,G22239,G22238);
  xor GNAME22251(G22251,G22252,G22161);
  xor GNAME22252(G22252,G18876,G22376);
  and GNAME22253(G22253,G18876,G22161);
  and GNAME22254(G22254,G22376,G22161);
  and GNAME22255(G22255,G18876,G22376);
  or GNAME22256(G22256,G22255,G22254,G22253);
  xor GNAME22266(G22266,G22267,G18891);
  xor GNAME22267(G22267,G19076,G18801);
  and GNAME22268(G22268,G19076,G18891);
  and GNAME22269(G22269,G18801,G18891);
  and GNAME22270(G22270,G19076,G18801);
  or GNAME22271(G22271,G22270,G22269,G22268);
  xor GNAME22281(G22281,G22282,G18906);
  xor GNAME22282(G22282,G19106,G18816);
  and GNAME22283(G22283,G19106,G18906);
  and GNAME22284(G22284,G18816,G18906);
  and GNAME22285(G22285,G19106,G18816);
  or GNAME22286(G22286,G22285,G22284,G22283);
  xor GNAME22296(G22296,G22297,G18921);
  xor GNAME22297(G22297,G19121,G18831);
  and GNAME22298(G22298,G19121,G18921);
  and GNAME22299(G22299,G18831,G18921);
  and GNAME22300(G22300,G19121,G18831);
  or GNAME22301(G22301,G22300,G22299,G22298);
  xor GNAME22311(G22311,G22312,G19166);
  xor GNAME22312(G22312,G19001,G18981);
  and GNAME22313(G22313,G19001,G19166);
  and GNAME22314(G22314,G18981,G19166);
  and GNAME22315(G22315,G19001,G18981);
  or GNAME22316(G22316,G22315,G22314,G22313);
  xor GNAME22326(G22326,G22327,G19181);
  xor GNAME22327(G22327,G22451,G18996);
  and GNAME22328(G22328,G22451,G19181);
  and GNAME22329(G22329,G18996,G19181);
  and GNAME22330(G22330,G22451,G18996);
  or GNAME22331(G22331,G22330,G22329,G22328);
  xor GNAME22341(G22341,G22342,G19196);
  xor GNAME22342(G22342,G19046,G19011);
  and GNAME22343(G22343,G19046,G19196);
  and GNAME22344(G22344,G19011,G19196);
  and GNAME22345(G22345,G19046,G19011);
  or GNAME22346(G22346,G22345,G22344,G22343);
  xor GNAME22356(G22356,G22357,G19211);
  xor GNAME22357(G22357,G22466,G19041);
  and GNAME22358(G22358,G22466,G19211);
  and GNAME22359(G22359,G19041,G19211);
  and GNAME22360(G22360,G22466,G19041);
  or GNAME22361(G22361,G22360,G22359,G22358);
  xor GNAME22371(G22371,G22372,G19226);
  xor GNAME22372(G22372,G19061,G19026);
  and GNAME22373(G22373,G19061,G19226);
  and GNAME22374(G22374,G19026,G19226);
  and GNAME22375(G22375,G19061,G19026);
  or GNAME22376(G22376,G22375,G22374,G22373);
  xor GNAME22386(G22386,G22387,G19241);
  xor GNAME22387(G22387,G22481,G19056);
  and GNAME22388(G22388,G22481,G19241);
  and GNAME22389(G22389,G19056,G19241);
  and GNAME22390(G22390,G22481,G19056);
  or GNAME22391(G22391,G22390,G22389,G22388);
  xor GNAME22401(G22401,G22402,G22326);
  xor GNAME22402(G22402,G19161,G24251);
  and GNAME22403(G22403,G19161,G22326);
  and GNAME22404(G22404,G24251,G22326);
  and GNAME22405(G22405,G19161,G24251);
  or GNAME22406(G22406,G22405,G22404,G22403);
  xor GNAME22416(G22416,G22417,G22356);
  xor GNAME22417(G22417,G19191,G24281);
  and GNAME22418(G22418,G19191,G22356);
  and GNAME22419(G22419,G24281,G22356);
  and GNAME22420(G22420,G19191,G24281);
  or GNAME22421(G22421,G22420,G22419,G22418);
  xor GNAME22431(G22431,G22432,G22386);
  xor GNAME22432(G22432,G19221,G24311);
  and GNAME22433(G22433,G19221,G22386);
  and GNAME22434(G22434,G24311,G22386);
  and GNAME22435(G22435,G19221,G24311);
  or GNAME22436(G22436,G22435,G22434,G22433);
  xor GNAME22446(G22446,G22447,G19301);
  xor GNAME22447(G22447,G19436,G19481);
  and GNAME22448(G22448,G19436,G19301);
  and GNAME22449(G22449,G19481,G19301);
  and GNAME22450(G22450,G19436,G19481);
  or GNAME22451(G22451,G22450,G22449,G22448);
  xor GNAME22461(G22461,G22462,G19316);
  xor GNAME22462(G22462,G19451,G19511);
  and GNAME22463(G22463,G19451,G19316);
  and GNAME22464(G22464,G19511,G19316);
  and GNAME22465(G22465,G19451,G19511);
  or GNAME22466(G22466,G22465,G22464,G22463);
  xor GNAME22476(G22476,G22477,G19331);
  xor GNAME22477(G22477,G19466,G19526);
  and GNAME22478(G22478,G19466,G19331);
  and GNAME22479(G22479,G19526,G19331);
  and GNAME22480(G22480,G19466,G19526);
  or GNAME22481(G22481,G22480,G22479,G22478);
  xor GNAME22491(G22491,G22492,G24246);
  xor GNAME22492(G22492,G19176,G24266);
  and GNAME22493(G22493,G19176,G24246);
  and GNAME22494(G22494,G24266,G24246);
  and GNAME22495(G22495,G19176,G24266);
  or GNAME22496(G22496,G22495,G22494,G22493);
  xor GNAME22506(G22506,G22507,G24276);
  xor GNAME22507(G22507,G19206,G24296);
  and GNAME22508(G22508,G19206,G24276);
  and GNAME22509(G22509,G24296,G24276);
  and GNAME22510(G22510,G19206,G24296);
  or GNAME22511(G22511,G22510,G22509,G22508);
  xor GNAME22521(G22521,G22522,G24306);
  xor GNAME22522(G22522,G19236,G24326);
  and GNAME22523(G22523,G19236,G24306);
  and GNAME22524(G22524,G24326,G24306);
  and GNAME22525(G22525,G19236,G24326);
  or GNAME22526(G22526,G22525,G22524,G22523);
  xor GNAME22536(G22536,G22537,G19346);
  xor GNAME22537(G22537,G19391,G19496);
  and GNAME22538(G22538,G19391,G19346);
  and GNAME22539(G22539,G19496,G19346);
  and GNAME22540(G22540,G19391,G19496);
  or GNAME22541(G22541,G22540,G22539,G22538);
  xor GNAME22551(G22551,G22552,G19361);
  xor GNAME22552(G22552,G19406,G19541);
  and GNAME22553(G22553,G19406,G19361);
  and GNAME22554(G22554,G19541,G19361);
  and GNAME22555(G22555,G19406,G19541);
  or GNAME22556(G22556,G22555,G22554,G22553);
  xor GNAME22566(G22566,G22567,G19376);
  xor GNAME22567(G22567,G19421,G19556);
  and GNAME22568(G22568,G19421,G19376);
  and GNAME22569(G22569,G19556,G19376);
  and GNAME22570(G22570,G19421,G19556);
  or GNAME22571(G22571,G22570,G22569,G22568);
  xor GNAME22581(G22581,G22582,G19476);
  xor GNAME22582(G22582,G19431,G19296);
  and GNAME22583(G22583,G19431,G19476);
  and GNAME22584(G22584,G19296,G19476);
  and GNAME22585(G22585,G19431,G19296);
  or GNAME22586(G22586,G22585,G22584,G22583);
  xor GNAME22596(G22596,G22597,G19491);
  xor GNAME22597(G22597,G19386,G19341);
  and GNAME22598(G22598,G19386,G19491);
  and GNAME22599(G22599,G19341,G19491);
  and GNAME22600(G22600,G19386,G19341);
  or GNAME22601(G22601,G22600,G22599,G22598);
  xor GNAME22611(G22611,G22612,G19506);
  xor GNAME22612(G22612,G19446,G19311);
  and GNAME22613(G22613,G19446,G19506);
  and GNAME22614(G22614,G19311,G19506);
  and GNAME22615(G22615,G19446,G19311);
  or GNAME22616(G22616,G22615,G22614,G22613);
  xor GNAME22626(G22626,G22627,G19536);
  xor GNAME22627(G22627,G19401,G19356);
  and GNAME22628(G22628,G19401,G19536);
  and GNAME22629(G22629,G19356,G19536);
  and GNAME22630(G22630,G19401,G19356);
  or GNAME22631(G22631,G22630,G22629,G22628);
  xor GNAME22641(G22641,G22642,G19521);
  xor GNAME22642(G22642,G19461,G19326);
  and GNAME22643(G22643,G19461,G19521);
  and GNAME22644(G22644,G19326,G19521);
  and GNAME22645(G22645,G19461,G19326);
  or GNAME22646(G22646,G22645,G22644,G22643);
  xor GNAME22656(G22656,G22657,G19551);
  xor GNAME22657(G22657,G19416,G19371);
  and GNAME22658(G22658,G19416,G19551);
  and GNAME22659(G22659,G19371,G19551);
  and GNAME22660(G22660,G19416,G19371);
  or GNAME22661(G22661,G22660,G22659,G22658);
  xor GNAME22671(G22671,G22672,G19571);
  xor GNAME22672(G22672,G19661,G19751);
  and GNAME22673(G22673,G19661,G19571);
  and GNAME22674(G22674,G19751,G19571);
  and GNAME22675(G22675,G19661,G19751);
  or GNAME22676(G22676,G22675,G22674,G22673);
  xor GNAME22686(G22686,G22687,G19586);
  xor GNAME22687(G22687,G19676,G19766);
  and GNAME22688(G22688,G19676,G19586);
  and GNAME22689(G22689,G19766,G19586);
  and GNAME22690(G22690,G19676,G19766);
  or GNAME22691(G22691,G22690,G22689,G22688);
  xor GNAME22701(G22701,G22702,G19601);
  xor GNAME22702(G22702,G19691,G19781);
  and GNAME22703(G22703,G19691,G19601);
  and GNAME22704(G22704,G19781,G19601);
  and GNAME22705(G22705,G19691,G19781);
  or GNAME22706(G22706,G22705,G22704,G22703);
  xor GNAME22716(G22716,G22717,G19616);
  xor GNAME22717(G22717,G19706,G19796);
  and GNAME22718(G22718,G19706,G19616);
  and GNAME22719(G22719,G19796,G19616);
  and GNAME22720(G22720,G19706,G19796);
  or GNAME22721(G22721,G22720,G22719,G22718);
  xor GNAME22731(G22731,G22732,G19631);
  xor GNAME22732(G22732,G19721,G19811);
  and GNAME22733(G22733,G19721,G19631);
  and GNAME22734(G22734,G19811,G19631);
  and GNAME22735(G22735,G19721,G19811);
  or GNAME22736(G22736,G22735,G22734,G22733);
  xor GNAME22746(G22746,G22747,G19646);
  xor GNAME22747(G22747,G19736,G19826);
  and GNAME22748(G22748,G19736,G19646);
  and GNAME22749(G22749,G19826,G19646);
  and GNAME22750(G22750,G19736,G19826);
  or GNAME22751(G22751,G22750,G22749,G22748);
  xor GNAME22761(G22761,G22762,G19746);
  xor GNAME22762(G22762,G19656,G19566);
  and GNAME22763(G22763,G19656,G19746);
  and GNAME22764(G22764,G19566,G19746);
  and GNAME22765(G22765,G19656,G19566);
  or GNAME22766(G22766,G22765,G22764,G22763);
  xor GNAME22776(G22776,G22777,G19761);
  xor GNAME22777(G22777,G19671,G19581);
  and GNAME22778(G22778,G19671,G19761);
  and GNAME22779(G22779,G19581,G19761);
  and GNAME22780(G22780,G19671,G19581);
  or GNAME22781(G22781,G22780,G22779,G22778);
  xor GNAME22791(G22791,G22792,G19776);
  xor GNAME22792(G22792,G19686,G19596);
  and GNAME22793(G22793,G19686,G19776);
  and GNAME22794(G22794,G19596,G19776);
  and GNAME22795(G22795,G19686,G19596);
  or GNAME22796(G22796,G22795,G22794,G22793);
  xor GNAME22806(G22806,G22807,G19806);
  xor GNAME22807(G22807,G19716,G19626);
  and GNAME22808(G22808,G19716,G19806);
  and GNAME22809(G22809,G19626,G19806);
  and GNAME22810(G22810,G19716,G19626);
  or GNAME22811(G22811,G22810,G22809,G22808);
  xor GNAME22821(G22821,G22822,G19791);
  xor GNAME22822(G22822,G19701,G19611);
  and GNAME22823(G22823,G19701,G19791);
  and GNAME22824(G22824,G19611,G19791);
  and GNAME22825(G22825,G19701,G19611);
  or GNAME22826(G22826,G22825,G22824,G22823);
  xor GNAME22836(G22836,G22837,G19821);
  xor GNAME22837(G22837,G19731,G19641);
  and GNAME22838(G22838,G19731,G19821);
  and GNAME22839(G22839,G19641,G19821);
  and GNAME22840(G22840,G19731,G19641);
  or GNAME22841(G22841,G22840,G22839,G22838);
  xor GNAME22851(G22851,G22852,G19841);
  xor GNAME22852(G22852,G19931,G20021);
  and GNAME22853(G22853,G19931,G19841);
  and GNAME22854(G22854,G20021,G19841);
  and GNAME22855(G22855,G19931,G20021);
  or GNAME22856(G22856,G22855,G22854,G22853);
  xor GNAME22866(G22866,G22867,G19856);
  xor GNAME22867(G22867,G19946,G20036);
  and GNAME22868(G22868,G19946,G19856);
  and GNAME22869(G22869,G20036,G19856);
  and GNAME22870(G22870,G19946,G20036);
  or GNAME22871(G22871,G22870,G22869,G22868);
  xor GNAME22881(G22881,G22882,G19871);
  xor GNAME22882(G22882,G19961,G20051);
  and GNAME22883(G22883,G19961,G19871);
  and GNAME22884(G22884,G20051,G19871);
  and GNAME22885(G22885,G19961,G20051);
  or GNAME22886(G22886,G22885,G22884,G22883);
  xor GNAME22896(G22896,G22897,G19886);
  xor GNAME22897(G22897,G19976,G20066);
  and GNAME22898(G22898,G19976,G19886);
  and GNAME22899(G22899,G20066,G19886);
  and GNAME22900(G22900,G19976,G20066);
  or GNAME22901(G22901,G22900,G22899,G22898);
  xor GNAME22911(G22911,G22912,G19901);
  xor GNAME22912(G22912,G19991,G20081);
  and GNAME22913(G22913,G19991,G19901);
  and GNAME22914(G22914,G20081,G19901);
  and GNAME22915(G22915,G19991,G20081);
  or GNAME22916(G22916,G22915,G22914,G22913);
  xor GNAME22926(G22926,G22927,G19916);
  xor GNAME22927(G22927,G20006,G20096);
  and GNAME22928(G22928,G20006,G19916);
  and GNAME22929(G22929,G20096,G19916);
  and GNAME22930(G22930,G20006,G20096);
  or GNAME22931(G22931,G22930,G22929,G22928);
  xor GNAME22941(G22941,G22942,G20016);
  xor GNAME22942(G22942,G19926,G19836);
  and GNAME22943(G22943,G19926,G20016);
  and GNAME22944(G22944,G19836,G20016);
  and GNAME22945(G22945,G19926,G19836);
  or GNAME22946(G22946,G22945,G22944,G22943);
  xor GNAME22956(G22956,G22957,G20031);
  xor GNAME22957(G22957,G19941,G19851);
  and GNAME22958(G22958,G19941,G20031);
  and GNAME22959(G22959,G19851,G20031);
  and GNAME22960(G22960,G19941,G19851);
  or GNAME22961(G22961,G22960,G22959,G22958);
  xor GNAME22971(G22971,G22972,G20046);
  xor GNAME22972(G22972,G19956,G19866);
  and GNAME22973(G22973,G19956,G20046);
  and GNAME22974(G22974,G19866,G20046);
  and GNAME22975(G22975,G19956,G19866);
  or GNAME22976(G22976,G22975,G22974,G22973);
  xor GNAME22986(G22986,G22987,G20076);
  xor GNAME22987(G22987,G19986,G19896);
  and GNAME22988(G22988,G19986,G20076);
  and GNAME22989(G22989,G19896,G20076);
  and GNAME22990(G22990,G19986,G19896);
  or GNAME22991(G22991,G22990,G22989,G22988);
  xor GNAME23001(G23001,G23002,G20061);
  xor GNAME23002(G23002,G19971,G19881);
  and GNAME23003(G23003,G19971,G20061);
  and GNAME23004(G23004,G19881,G20061);
  and GNAME23005(G23005,G19971,G19881);
  or GNAME23006(G23006,G23005,G23004,G23003);
  xor GNAME23016(G23016,G23017,G20091);
  xor GNAME23017(G23017,G20001,G19911);
  and GNAME23018(G23018,G20001,G20091);
  and GNAME23019(G23019,G19911,G20091);
  and GNAME23020(G23020,G20001,G19911);
  or GNAME23021(G23021,G23020,G23019,G23018);
  xor GNAME23031(G23031,G23032,G20111);
  xor GNAME23032(G23032,G20201,G20291);
  and GNAME23033(G23033,G20201,G20111);
  and GNAME23034(G23034,G20291,G20111);
  and GNAME23035(G23035,G20201,G20291);
  or GNAME23036(G23036,G23035,G23034,G23033);
  xor GNAME23046(G23046,G23047,G20126);
  xor GNAME23047(G23047,G20216,G20306);
  and GNAME23048(G23048,G20216,G20126);
  and GNAME23049(G23049,G20306,G20126);
  and GNAME23050(G23050,G20216,G20306);
  or GNAME23051(G23051,G23050,G23049,G23048);
  xor GNAME23061(G23061,G23062,G20141);
  xor GNAME23062(G23062,G20231,G20321);
  and GNAME23063(G23063,G20231,G20141);
  and GNAME23064(G23064,G20321,G20141);
  and GNAME23065(G23065,G20231,G20321);
  or GNAME23066(G23066,G23065,G23064,G23063);
  xor GNAME23076(G23076,G23077,G20156);
  xor GNAME23077(G23077,G20246,G20336);
  and GNAME23078(G23078,G20246,G20156);
  and GNAME23079(G23079,G20336,G20156);
  and GNAME23080(G23080,G20246,G20336);
  or GNAME23081(G23081,G23080,G23079,G23078);
  xor GNAME23091(G23091,G23092,G20171);
  xor GNAME23092(G23092,G20261,G20351);
  and GNAME23093(G23093,G20261,G20171);
  and GNAME23094(G23094,G20351,G20171);
  and GNAME23095(G23095,G20261,G20351);
  or GNAME23096(G23096,G23095,G23094,G23093);
  xor GNAME23106(G23106,G23107,G20186);
  xor GNAME23107(G23107,G20276,G20366);
  and GNAME23108(G23108,G20276,G20186);
  and GNAME23109(G23109,G20366,G20186);
  and GNAME23110(G23110,G20276,G20366);
  or GNAME23111(G23111,G23110,G23109,G23108);
  xor GNAME23121(G23121,G23122,G20286);
  xor GNAME23122(G23122,G20196,G20106);
  and GNAME23123(G23123,G20196,G20286);
  and GNAME23124(G23124,G20106,G20286);
  and GNAME23125(G23125,G20196,G20106);
  or GNAME23126(G23126,G23125,G23124,G23123);
  xor GNAME23136(G23136,G23137,G20301);
  xor GNAME23137(G23137,G20211,G20121);
  and GNAME23138(G23138,G20211,G20301);
  and GNAME23139(G23139,G20121,G20301);
  and GNAME23140(G23140,G20211,G20121);
  or GNAME23141(G23141,G23140,G23139,G23138);
  xor GNAME23151(G23151,G23152,G20316);
  xor GNAME23152(G23152,G20226,G20136);
  and GNAME23153(G23153,G20226,G20316);
  and GNAME23154(G23154,G20136,G20316);
  and GNAME23155(G23155,G20226,G20136);
  or GNAME23156(G23156,G23155,G23154,G23153);
  xor GNAME23166(G23166,G23167,G20346);
  xor GNAME23167(G23167,G20256,G20166);
  and GNAME23168(G23168,G20256,G20346);
  and GNAME23169(G23169,G20166,G20346);
  and GNAME23170(G23170,G20256,G20166);
  or GNAME23171(G23171,G23170,G23169,G23168);
  xor GNAME23181(G23181,G23182,G20331);
  xor GNAME23182(G23182,G20241,G20151);
  and GNAME23183(G23183,G20241,G20331);
  and GNAME23184(G23184,G20151,G20331);
  and GNAME23185(G23185,G20241,G20151);
  or GNAME23186(G23186,G23185,G23184,G23183);
  xor GNAME23196(G23196,G23197,G20361);
  xor GNAME23197(G23197,G20271,G20181);
  and GNAME23198(G23198,G20271,G20361);
  and GNAME23199(G23199,G20181,G20361);
  and GNAME23200(G23200,G20271,G20181);
  or GNAME23201(G23201,G23200,G23199,G23198);
  xor GNAME23211(G23211,G23212,G23351);
  xor GNAME23212(G23212,G20381,G23301);
  and GNAME23213(G23213,G20381,G23351);
  and GNAME23214(G23214,G23301,G23351);
  and GNAME23215(G23215,G20381,G23301);
  or GNAME23216(G23216,G23215,G23214,G23213);
  xor GNAME23226(G23226,G23227,G20516);
  xor GNAME23227(G23227,G20741,G20376);
  and GNAME23228(G23228,G20741,G20516);
  and GNAME23229(G23229,G20376,G20516);
  and GNAME23230(G23230,G20741,G20376);
  or GNAME23231(G23231,G23230,G23229,G23228);
  xor GNAME23241(G23241,G23242,G23366);
  xor GNAME23242(G23242,G20396,G23316);
  and GNAME23243(G23243,G20396,G23366);
  and GNAME23244(G23244,G23316,G23366);
  and GNAME23245(G23245,G20396,G23316);
  or GNAME23246(G23246,G23245,G23244,G23243);
  xor GNAME23256(G23256,G23257,G20531);
  xor GNAME23257(G23257,G20756,G20391);
  and GNAME23258(G23258,G20756,G20531);
  and GNAME23259(G23259,G20391,G20531);
  and GNAME23260(G23260,G20756,G20391);
  or GNAME23261(G23261,G23260,G23259,G23258);
  xor GNAME23271(G23271,G23272,G23381);
  xor GNAME23272(G23272,G20411,G23331);
  and GNAME23273(G23273,G20411,G23381);
  and GNAME23274(G23274,G23331,G23381);
  and GNAME23275(G23275,G20411,G23331);
  or GNAME23276(G23276,G23275,G23274,G23273);
  xor GNAME23286(G23286,G23287,G20546);
  xor GNAME23287(G23287,G20771,G20406);
  and GNAME23288(G23288,G20771,G20546);
  and GNAME23289(G23289,G20406,G20546);
  and GNAME23290(G23290,G20771,G20406);
  or GNAME23291(G23291,G23290,G23289,G23288);
  xor GNAME23301(G23301,G23302,G20426);
  xor GNAME23302(G23302,G20561,G20606);
  and GNAME23303(G23303,G20561,G20426);
  and GNAME23304(G23304,G20606,G20426);
  and GNAME23305(G23305,G20561,G20606);
  or GNAME23306(G23306,G23305,G23304,G23303);
  xor GNAME23316(G23316,G23317,G20456);
  xor GNAME23317(G23317,G20576,G20636);
  and GNAME23318(G23318,G20576,G20456);
  and GNAME23319(G23319,G20636,G20456);
  and GNAME23320(G23320,G20576,G20636);
  or GNAME23321(G23321,G23320,G23319,G23318);
  xor GNAME23331(G23331,G23332,G20471);
  xor GNAME23332(G23332,G20591,G20651);
  and GNAME23333(G23333,G20591,G20471);
  and GNAME23334(G23334,G20651,G20471);
  and GNAME23335(G23335,G20591,G20651);
  or GNAME23336(G23336,G23335,G23334,G23333);
  xor GNAME23346(G23346,G23347,G20601);
  xor GNAME23347(G23347,G20556,G20421);
  and GNAME23348(G23348,G20556,G20601);
  and GNAME23349(G23349,G20421,G20601);
  and GNAME23350(G23350,G20556,G20421);
  or GNAME23351(G23351,G23350,G23349,G23348);
  xor GNAME23361(G23361,G23362,G20631);
  xor GNAME23362(G23362,G20571,G20451);
  and GNAME23363(G23363,G20571,G20631);
  and GNAME23364(G23364,G20451,G20631);
  and GNAME23365(G23365,G20571,G20451);
  or GNAME23366(G23366,G23365,G23364,G23363);
  xor GNAME23376(G23376,G23377,G20646);
  xor GNAME23377(G23377,G20586,G20466);
  and GNAME23378(G23378,G20586,G20646);
  and GNAME23379(G23379,G20466,G20646);
  and GNAME23380(G23380,G20586,G20466);
  or GNAME23381(G23381,G23380,G23379,G23378);
  xor GNAME23391(G23391,G23392,G20736);
  xor GNAME23392(G23392,G20831,G23531);
  and GNAME23393(G23393,G20831,G20736);
  and GNAME23394(G23394,G23531,G20736);
  and GNAME23395(G23395,G20831,G23531);
  or GNAME23396(G23396,G23395,G23394,G23393);
  xor GNAME23406(G23406,G23407,G20876);
  xor GNAME23407(G23407,G20916,G20826);
  and GNAME23408(G23408,G20916,G20876);
  and GNAME23409(G23409,G20826,G20876);
  and GNAME23410(G23410,G20916,G20826);
  or GNAME23411(G23411,G23410,G23409,G23408);
  xor GNAME23421(G23421,G23422,G20751);
  xor GNAME23422(G23422,G20846,G23546);
  and GNAME23423(G23423,G20846,G20751);
  and GNAME23424(G23424,G23546,G20751);
  and GNAME23425(G23425,G20846,G23546);
  or GNAME23426(G23426,G23425,G23424,G23423);
  xor GNAME23436(G23436,G23437,G20891);
  xor GNAME23437(G23437,G20946,G20841);
  and GNAME23438(G23438,G20946,G20891);
  and GNAME23439(G23439,G20841,G20891);
  and GNAME23440(G23440,G20946,G20841);
  or GNAME23441(G23441,G23440,G23439,G23438);
  xor GNAME23451(G23451,G23452,G20766);
  xor GNAME23452(G23452,G20861,G23561);
  and GNAME23453(G23453,G20861,G20766);
  and GNAME23454(G23454,G23561,G20766);
  and GNAME23455(G23455,G20861,G23561);
  or GNAME23456(G23456,G23455,G23454,G23453);
  xor GNAME23466(G23466,G23467,G20906);
  xor GNAME23467(G23467,G20961,G20856);
  and GNAME23468(G23468,G20961,G20906);
  and GNAME23469(G23469,G20856,G20906);
  and GNAME23470(G23470,G20961,G20856);
  or GNAME23471(G23471,G23470,G23469,G23468);
  xor GNAME23481(G23481,G23482,G23391);
  xor GNAME23482(G23482,G20511,G23411);
  and GNAME23483(G23483,G20511,G23391);
  and GNAME23484(G23484,G23411,G23391);
  and GNAME23485(G23485,G20511,G23411);
  or GNAME23486(G23486,G23485,G23484,G23483);
  xor GNAME23496(G23496,G23497,G23421);
  xor GNAME23497(G23497,G20526,G23441);
  and GNAME23498(G23498,G20526,G23421);
  and GNAME23499(G23499,G23441,G23421);
  and GNAME23500(G23500,G20526,G23441);
  or GNAME23501(G23501,G23500,G23499,G23498);
  xor GNAME23511(G23511,G23512,G23451);
  xor GNAME23512(G23512,G20541,G23471);
  and GNAME23513(G23513,G20541,G23451);
  and GNAME23514(G23514,G23471,G23451);
  and GNAME23515(G23515,G20541,G23471);
  or GNAME23516(G23516,G23515,G23514,G23513);
  xor GNAME23526(G23526,G23527,G20691);
  xor GNAME23527(G23527,G20936,G20786);
  and GNAME23528(G23528,G20936,G20691);
  and GNAME23529(G23529,G20786,G20691);
  and GNAME23530(G23530,G20936,G20786);
  or GNAME23531(G23531,G23530,G23529,G23528);
  xor GNAME23541(G23541,G23542,G20706);
  xor GNAME23542(G23542,G20981,G20801);
  and GNAME23543(G23543,G20981,G20706);
  and GNAME23544(G23544,G20801,G20706);
  and GNAME23545(G23545,G20981,G20801);
  or GNAME23546(G23546,G23545,G23544,G23543);
  xor GNAME23556(G23556,G23557,G20721);
  xor GNAME23557(G23557,G20996,G20816);
  and GNAME23558(G23558,G20996,G20721);
  and GNAME23559(G23559,G20816,G20721);
  and GNAME23560(G23560,G20996,G20816);
  or GNAME23561(G23561,G23560,G23559,G23558);
  xor GNAME23571(G23571,G23572,G21146);
  xor GNAME23572(G23572,G20931,G20781);
  and GNAME23573(G23573,G20931,G21146);
  and GNAME23574(G23574,G20781,G21146);
  and GNAME23575(G23575,G20931,G20781);
  or GNAME23576(G23576,G23575,G23574,G23573);
  xor GNAME23586(G23586,G23587,G21191);
  xor GNAME23587(G23587,G21276,G21051);
  and GNAME23588(G23588,G21276,G21191);
  and GNAME23589(G23589,G21051,G21191);
  and GNAME23590(G23590,G21276,G21051);
  or GNAME23591(G23591,G23590,G23589,G23588);
  xor GNAME23601(G23601,G23602,G21161);
  xor GNAME23602(G23602,G20976,G20796);
  and GNAME23603(G23603,G20976,G21161);
  and GNAME23604(G23604,G20796,G21161);
  and GNAME23605(G23605,G20976,G20796);
  or GNAME23606(G23606,G23605,G23604,G23603);
  xor GNAME23616(G23616,G23617,G21221);
  xor GNAME23617(G23617,G21291,G21081);
  and GNAME23618(G23618,G21291,G21221);
  and GNAME23619(G23619,G21081,G21221);
  and GNAME23620(G23620,G21291,G21081);
  or GNAME23621(G23621,G23620,G23619,G23618);
  xor GNAME23631(G23631,G23632,G21176);
  xor GNAME23632(G23632,G20991,G20811);
  and GNAME23633(G23633,G20991,G21176);
  and GNAME23634(G23634,G20811,G21176);
  and GNAME23635(G23635,G20991,G20811);
  or GNAME23636(G23636,G23635,G23634,G23633);
  xor GNAME23646(G23646,G23647,G21236);
  xor GNAME23647(G23647,G21306,G21096);
  and GNAME23648(G23648,G21306,G21236);
  and GNAME23649(G23649,G21096,G21236);
  and GNAME23650(G23650,G21306,G21096);
  or GNAME23651(G23651,G23650,G23649,G23648);
  xor GNAME23661(G23661,G23662,G23571);
  xor GNAME23662(G23662,G20871,G23591);
  and GNAME23663(G23663,G20871,G23571);
  and GNAME23664(G23664,G23591,G23571);
  and GNAME23665(G23665,G20871,G23591);
  or GNAME23666(G23666,G23665,G23664,G23663);
  xor GNAME23676(G23676,G23677,G23586);
  xor GNAME23677(G23677,G21141,G21011);
  and GNAME23678(G23678,G21141,G23586);
  and GNAME23679(G23679,G21011,G23586);
  and GNAME23680(G23680,G21141,G21011);
  or GNAME23681(G23681,G23680,G23679,G23678);
  xor GNAME23691(G23691,G23692,G21006);
  xor GNAME23692(G23692,G21186,G21371);
  and GNAME23693(G23693,G21186,G21006);
  and GNAME23694(G23694,G21371,G21006);
  and GNAME23695(G23695,G21186,G21371);
  or GNAME23696(G23696,G23695,G23694,G23693);
  xor GNAME23706(G23706,G23707,G23601);
  xor GNAME23707(G23707,G20886,G23621);
  and GNAME23708(G23708,G20886,G23601);
  and GNAME23709(G23709,G23621,G23601);
  and GNAME23710(G23710,G20886,G23621);
  or GNAME23711(G23711,G23710,G23709,G23708);
  xor GNAME23721(G23721,G23722,G23631);
  xor GNAME23722(G23722,G20901,G23651);
  and GNAME23723(G23723,G20901,G23631);
  and GNAME23724(G23724,G23651,G23631);
  and GNAME23725(G23725,G20901,G23651);
  or GNAME23726(G23726,G23725,G23724,G23723);
  xor GNAME23736(G23736,G23737,G23616);
  xor GNAME23737(G23737,G21156,G21026);
  and GNAME23738(G23738,G21156,G23616);
  and GNAME23739(G23739,G21026,G23616);
  and GNAME23740(G23740,G21156,G21026);
  or GNAME23741(G23741,G23740,G23739,G23738);
  xor GNAME23751(G23751,G23752,G21021);
  xor GNAME23752(G23752,G21216,G21401);
  and GNAME23753(G23753,G21216,G21021);
  and GNAME23754(G23754,G21401,G21021);
  and GNAME23755(G23755,G21216,G21401);
  or GNAME23756(G23756,G23755,G23754,G23753);
  xor GNAME23766(G23766,G23767,G23646);
  xor GNAME23767(G23767,G21171,G21041);
  and GNAME23768(G23768,G21171,G23646);
  and GNAME23769(G23769,G21041,G23646);
  and GNAME23770(G23770,G21171,G21041);
  or GNAME23771(G23771,G23770,G23769,G23768);
  xor GNAME23781(G23781,G23782,G21036);
  xor GNAME23782(G23782,G21231,G21416);
  and GNAME23783(G23783,G21231,G21036);
  and GNAME23784(G23784,G21416,G21036);
  and GNAME23785(G23785,G21231,G21416);
  or GNAME23786(G23786,G23785,G23784,G23783);
  xor GNAME23796(G23796,G23797,G21366);
  xor GNAME23797(G23797,G21201,G21386);
  and GNAME23798(G23798,G21201,G21366);
  and GNAME23799(G23799,G21386,G21366);
  and GNAME23800(G23800,G21201,G21386);
  or GNAME23801(G23801,G23800,G23799,G23798);
  xor GNAME23811(G23811,G23812,G21381);
  xor GNAME23812(G23812,G21501,G21641);
  and GNAME23813(G23813,G21501,G21381);
  and GNAME23814(G23814,G21641,G21381);
  and GNAME23815(G23815,G21501,G21641);
  or GNAME23816(G23816,G23815,G23814,G23813);
  xor GNAME23826(G23826,G23827,G21396);
  xor GNAME23827(G23827,G21246,G21431);
  and GNAME23828(G23828,G21246,G21396);
  and GNAME23829(G23829,G21431,G21396);
  and GNAME23830(G23830,G21246,G21431);
  or GNAME23831(G23831,G23830,G23829,G23828);
  xor GNAME23841(G23841,G23842,G21426);
  xor GNAME23842(G23842,G21516,G21656);
  and GNAME23843(G23843,G21516,G21426);
  and GNAME23844(G23844,G21656,G21426);
  and GNAME23845(G23845,G21516,G21656);
  or GNAME23846(G23846,G23845,G23844,G23843);
  xor GNAME23856(G23856,G23857,G21411);
  xor GNAME23857(G23857,G21261,G21446);
  and GNAME23858(G23858,G21261,G21411);
  and GNAME23859(G23859,G21446,G21411);
  and GNAME23860(G23860,G21261,G21446);
  or GNAME23861(G23861,G23860,G23859,G23858);
  xor GNAME23871(G23871,G23872,G21441);
  xor GNAME23872(G23872,G21531,G21671);
  and GNAME23873(G23873,G21531,G21441);
  and GNAME23874(G23874,G21671,G21441);
  and GNAME23875(G23875,G21531,G21671);
  or GNAME23876(G23876,G23875,G23874,G23873);
  xor GNAME23886(G23886,G23887,G21636);
  xor GNAME23887(G23887,G21596,G21456);
  and GNAME23888(G23888,G21596,G21636);
  and GNAME23889(G23889,G21456,G21636);
  and GNAME23890(G23890,G21596,G21456);
  or GNAME23891(G23891,G23890,G23889,G23888);
  xor GNAME23901(G23901,G23902,G21651);
  xor GNAME23902(G23902,G21611,G21471);
  and GNAME23903(G23903,G21611,G21651);
  and GNAME23904(G23904,G21471,G21651);
  and GNAME23905(G23905,G21611,G21471);
  or GNAME23906(G23906,G23905,G23904,G23903);
  xor GNAME23916(G23916,G23917,G21666);
  xor GNAME23917(G23917,G21626,G21486);
  and GNAME23918(G23918,G21626,G21666);
  and GNAME23919(G23919,G21486,G21666);
  and GNAME23920(G23920,G21626,G21486);
  or GNAME23921(G23921,G23920,G23919,G23918);
  xor GNAME23931(G23931,G23932,G23951);
  xor GNAME23932(G23932,G17946,G17996);
  and GNAME23933(G23933,G17946,G23951);
  and GNAME23934(G23934,G17996,G23951);
  and GNAME23935(G23935,G17946,G17996);
  or GNAME23936(G23936,G23935,G23934,G23933);
  xor GNAME23946(G23946,G23947,G23966);
  xor GNAME23947(G23947,G18131,G17991);
  and GNAME23948(G23948,G18131,G23966);
  and GNAME23949(G23949,G17991,G23966);
  and GNAME23950(G23950,G18131,G17991);
  or GNAME23951(G23951,G23950,G23949,G23948);
  xor GNAME23961(G23961,G23962,G25061);
  xor GNAME23962(G23962,G21866,G18126);
  and GNAME23963(G23963,G21866,G25061);
  and GNAME23964(G23964,G18126,G25061);
  and GNAME23965(G23965,G21866,G18126);
  or GNAME23966(G23966,G23965,G23964,G23963);
  xor GNAME23976(G23976,G23977,G24011);
  xor GNAME23977(G23977,G17961,G18011);
  and GNAME23978(G23978,G17961,G24011);
  and GNAME23979(G23979,G18011,G24011);
  and GNAME23980(G23980,G17961,G18011);
  or GNAME23981(G23981,G23980,G23979,G23978);
  xor GNAME23991(G23991,G23992,G24041);
  xor GNAME23992(G23992,G17976,G18026);
  and GNAME23993(G23993,G17976,G24041);
  and GNAME23994(G23994,G18026,G24041);
  and GNAME23995(G23995,G17976,G18026);
  or GNAME23996(G23996,G23995,G23994,G23993);
  xor GNAME24006(G24006,G24007,G24026);
  xor GNAME24007(G24007,G18146,G18006);
  and GNAME24008(G24008,G18146,G24026);
  and GNAME24009(G24009,G18006,G24026);
  and GNAME24010(G24010,G18146,G18006);
  or GNAME24011(G24011,G24010,G24009,G24008);
  xor GNAME24021(G24021,G24022,G25196);
  xor GNAME24022(G24022,G21881,G18141);
  and GNAME24023(G24023,G21881,G25196);
  and GNAME24024(G24024,G18141,G25196);
  and GNAME24025(G24025,G21881,G18141);
  or GNAME24026(G24026,G24025,G24024,G24023);
  xor GNAME24036(G24036,G24037,G24056);
  xor GNAME24037(G24037,G18161,G18021);
  and GNAME24038(G24038,G18161,G24056);
  and GNAME24039(G24039,G18021,G24056);
  and GNAME24040(G24040,G18161,G18021);
  or GNAME24041(G24041,G24040,G24039,G24038);
  xor GNAME24051(G24051,G24052,G25226);
  xor GNAME24052(G24052,G21896,G18156);
  and GNAME24053(G24053,G21896,G25226);
  and GNAME24054(G24054,G18156,G25226);
  and GNAME24055(G24055,G21896,G18156);
  or GNAME24056(G24056,G24055,G24054,G24053);
  xor GNAME24066(G24066,G24067,G24086);
  xor GNAME24067(G24067,G21701,G23886);
  and GNAME24068(G24068,G21701,G24086);
  and GNAME24069(G24069,G23886,G24086);
  and GNAME24070(G24070,G21701,G23886);
  or GNAME24071(G24071,G24070,G24069,G24068);
  xor GNAME24081(G24081,G24082,G21791);
  xor GNAME24082(G24082,G21686,G21696);
  and GNAME24083(G24083,G21686,G21791);
  and GNAME24084(G24084,G21696,G21791);
  and GNAME24085(G24085,G21686,G21696);
  or GNAME24086(G24086,G24085,G24084,G24083);
  xor GNAME24096(G24096,G24097,G24131);
  xor GNAME24097(G24097,G21716,G23901);
  and GNAME24098(G24098,G21716,G24131);
  and GNAME24099(G24099,G23901,G24131);
  and GNAME24100(G24100,G21716,G23901);
  or GNAME24101(G24101,G24100,G24099,G24098);
  xor GNAME24111(G24111,G24112,G24146);
  xor GNAME24112(G24112,G21731,G23916);
  and GNAME24113(G24113,G21731,G24146);
  and GNAME24114(G24114,G23916,G24146);
  and GNAME24115(G24115,G21731,G23916);
  or GNAME24116(G24116,G24115,G24114,G24113);
  xor GNAME24126(G24126,G24127,G21821);
  xor GNAME24127(G24127,G21746,G21711);
  and GNAME24128(G24128,G21746,G21821);
  and GNAME24129(G24129,G21711,G21821);
  and GNAME24130(G24130,G21746,G21711);
  or GNAME24131(G24131,G24130,G24129,G24128);
  xor GNAME24141(G24141,G24142,G21851);
  xor GNAME24142(G24142,G21761,G21726);
  and GNAME24143(G24143,G21761,G21851);
  and GNAME24144(G24144,G21726,G21851);
  and GNAME24145(G24145,G21761,G21726);
  or GNAME24146(G24146,G24145,G24144,G24143);
  xor GNAME24156(G24156,G24157,G23936);
  xor GNAME24157(G24157,G17951,G17901);
  and GNAME24158(G24158,G17951,G23936);
  and GNAME24159(G24159,G17901,G23936);
  and GNAME24160(G24160,G17951,G17901);
  or GNAME24161(G24161,G24160,G24159,G24158);
  xor GNAME24171(G24171,G24172,G23981);
  xor GNAME24172(G24172,G17966,G17916);
  and GNAME24173(G24173,G17966,G23981);
  and GNAME24174(G24174,G17916,G23981);
  and GNAME24175(G24175,G17966,G17916);
  or GNAME24176(G24176,G24175,G24174,G24173);
  xor GNAME24186(G24186,G24187,G23996);
  xor GNAME24187(G24187,G17981,G17931);
  and GNAME24188(G24188,G17981,G23996);
  and GNAME24189(G24189,G17931,G23996);
  and GNAME24190(G24190,G17981,G17931);
  or GNAME24191(G24191,G24190,G24189,G24188);
  xor GNAME24201(G24201,G24202,G22311);
  xor GNAME24202(G24202,G22266,G22331);
  and GNAME24203(G24203,G22266,G22311);
  and GNAME24204(G24204,G22331,G22311);
  and GNAME24205(G24205,G22266,G22331);
  or GNAME24206(G24206,G24205,G24204,G24203);
  xor GNAME24216(G24216,G24217,G22341);
  xor GNAME24217(G24217,G22281,G22361);
  and GNAME24218(G24218,G22281,G22341);
  and GNAME24219(G24219,G22361,G22341);
  and GNAME24220(G24220,G22281,G22361);
  or GNAME24221(G24221,G24220,G24219,G24218);
  xor GNAME24231(G24231,G24232,G22371);
  xor GNAME24232(G24232,G22296,G22391);
  and GNAME24233(G24233,G22296,G22371);
  and GNAME24234(G24234,G22391,G22371);
  and GNAME24235(G24235,G22296,G22391);
  or GNAME24236(G24236,G24235,G24234,G24233);
  xor GNAME24246(G24246,G24247,G22446);
  xor GNAME24247(G24247,G22541,G22586);
  and GNAME24248(G24248,G22541,G22446);
  and GNAME24249(G24249,G22586,G22446);
  and GNAME24250(G24250,G22541,G22586);
  or GNAME24251(G24251,G24250,G24249,G24248);
  xor GNAME24261(G24261,G24262,G22601);
  xor GNAME24262(G24262,G22676,G22536);
  and GNAME24263(G24263,G22676,G22601);
  and GNAME24264(G24264,G22536,G22601);
  and GNAME24265(G24265,G22676,G22536);
  or GNAME24266(G24266,G24265,G24264,G24263);
  xor GNAME24276(G24276,G24277,G22461);
  xor GNAME24277(G24277,G22556,G22616);
  and GNAME24278(G24278,G22556,G22461);
  and GNAME24279(G24279,G22616,G22461);
  and GNAME24280(G24280,G22556,G22616);
  or GNAME24281(G24281,G24280,G24279,G24278);
  xor GNAME24291(G24291,G24292,G22631);
  xor GNAME24292(G24292,G22706,G22551);
  and GNAME24293(G24293,G22706,G22631);
  and GNAME24294(G24294,G22551,G22631);
  and GNAME24295(G24295,G22706,G22551);
  or GNAME24296(G24296,G24295,G24294,G24293);
  xor GNAME24306(G24306,G24307,G22476);
  xor GNAME24307(G24307,G22571,G22646);
  and GNAME24308(G24308,G22571,G22476);
  and GNAME24309(G24309,G22646,G22476);
  and GNAME24310(G24310,G22571,G22646);
  or GNAME24311(G24311,G24310,G24309,G24308);
  xor GNAME24321(G24321,G24322,G22661);
  xor GNAME24322(G24322,G22721,G22566);
  and GNAME24323(G24323,G22721,G22661);
  and GNAME24324(G24324,G22566,G22661);
  and GNAME24325(G24325,G22721,G22566);
  or GNAME24326(G24326,G24325,G24324,G24323);
  xor GNAME24336(G24336,G24337,G24261);
  xor GNAME24337(G24337,G22581,G24386);
  and GNAME24338(G24338,G22581,G24261);
  and GNAME24339(G24339,G24386,G24261);
  and GNAME24340(G24340,G22581,G24386);
  or GNAME24341(G24341,G24340,G24339,G24338);
  xor GNAME24351(G24351,G24352,G24291);
  xor GNAME24352(G24352,G22611,G24416);
  and GNAME24353(G24353,G22611,G24291);
  and GNAME24354(G24354,G24416,G24291);
  and GNAME24355(G24355,G22611,G24416);
  or GNAME24356(G24356,G24355,G24354,G24353);
  xor GNAME24366(G24366,G24367,G24321);
  xor GNAME24367(G24367,G22641,G24446);
  and GNAME24368(G24368,G22641,G24321);
  and GNAME24369(G24369,G24446,G24321);
  and GNAME24370(G24370,G22641,G24446);
  or GNAME24371(G24371,G24370,G24369,G24368);
  xor GNAME24381(G24381,G24382,G22766);
  xor GNAME24382(G24382,G22691,G22671);
  and GNAME24383(G24383,G22691,G22766);
  and GNAME24384(G24384,G22671,G22766);
  and GNAME24385(G24385,G22691,G22671);
  or GNAME24386(G24386,G24385,G24384,G24383);
  xor GNAME24396(G24396,G24397,G22781);
  xor GNAME24397(G24397,G22856,G22686);
  and GNAME24398(G24398,G22856,G22781);
  and GNAME24399(G24399,G22686,G22781);
  and GNAME24400(G24400,G22856,G22686);
  or GNAME24401(G24401,G24400,G24399,G24398);
  xor GNAME24411(G24411,G24412,G22796);
  xor GNAME24412(G24412,G22736,G22701);
  and GNAME24413(G24413,G22736,G22796);
  and GNAME24414(G24414,G22701,G22796);
  and GNAME24415(G24415,G22736,G22701);
  or GNAME24416(G24416,G24415,G24414,G24413);
  xor GNAME24426(G24426,G24427,G22811);
  xor GNAME24427(G24427,G22886,G22731);
  and GNAME24428(G24428,G22886,G22811);
  and GNAME24429(G24429,G22731,G22811);
  and GNAME24430(G24430,G22886,G22731);
  or GNAME24431(G24431,G24430,G24429,G24428);
  xor GNAME24441(G24441,G24442,G22826);
  xor GNAME24442(G24442,G22751,G22716);
  and GNAME24443(G24443,G22751,G22826);
  and GNAME24444(G24444,G22716,G22826);
  and GNAME24445(G24445,G22751,G22716);
  or GNAME24446(G24446,G24445,G24444,G24443);
  xor GNAME24456(G24456,G24457,G22841);
  xor GNAME24457(G24457,G22901,G22746);
  and GNAME24458(G24458,G22901,G22841);
  and GNAME24459(G24459,G22746,G22841);
  and GNAME24460(G24460,G22901,G22746);
  or GNAME24461(G24461,G24460,G24459,G24458);
  xor GNAME24471(G24471,G24472,G24381);
  xor GNAME24472(G24472,G22596,G24401);
  and GNAME24473(G24473,G22596,G24381);
  and GNAME24474(G24474,G24401,G24381);
  and GNAME24475(G24475,G22596,G24401);
  or GNAME24476(G24476,G24475,G24474,G24473);
  xor GNAME24486(G24486,G24487,G24396);
  xor GNAME24487(G24487,G22761,G24566);
  and GNAME24488(G24488,G22761,G24396);
  and GNAME24489(G24489,G24566,G24396);
  and GNAME24490(G24490,G22761,G24566);
  or GNAME24491(G24491,G24490,G24489,G24488);
  xor GNAME24501(G24501,G24502,G24411);
  xor GNAME24502(G24502,G22626,G24431);
  and GNAME24503(G24503,G22626,G24411);
  and GNAME24504(G24504,G24431,G24411);
  and GNAME24505(G24505,G22626,G24431);
  or GNAME24506(G24506,G24505,G24504,G24503);
  xor GNAME24516(G24516,G24517,G24441);
  xor GNAME24517(G24517,G22656,G24461);
  and GNAME24518(G24518,G22656,G24441);
  and GNAME24519(G24519,G24461,G24441);
  and GNAME24520(G24520,G22656,G24461);
  or GNAME24521(G24521,G24520,G24519,G24518);
  xor GNAME24531(G24531,G24532,G24426);
  xor GNAME24532(G24532,G22791,G24596);
  and GNAME24533(G24533,G22791,G24426);
  and GNAME24534(G24534,G24596,G24426);
  and GNAME24535(G24535,G22791,G24596);
  or GNAME24536(G24536,G24535,G24534,G24533);
  xor GNAME24546(G24546,G24547,G24456);
  xor GNAME24547(G24547,G22821,G24626);
  and GNAME24548(G24548,G22821,G24456);
  and GNAME24549(G24549,G24626,G24456);
  and GNAME24550(G24550,G22821,G24626);
  or GNAME24551(G24551,G24550,G24549,G24548);
  xor GNAME24561(G24561,G24562,G22946);
  xor GNAME24562(G24562,G22871,G22851);
  and GNAME24563(G24563,G22871,G22946);
  and GNAME24564(G24564,G22851,G22946);
  and GNAME24565(G24565,G22871,G22851);
  or GNAME24566(G24566,G24565,G24564,G24563);
  xor GNAME24576(G24576,G24577,G22961);
  xor GNAME24577(G24577,G23036,G22866);
  and GNAME24578(G24578,G23036,G22961);
  and GNAME24579(G24579,G22866,G22961);
  and GNAME24580(G24580,G23036,G22866);
  or GNAME24581(G24581,G24580,G24579,G24578);
  xor GNAME24591(G24591,G24592,G22976);
  xor GNAME24592(G24592,G22916,G22881);
  and GNAME24593(G24593,G22916,G22976);
  and GNAME24594(G24594,G22881,G22976);
  and GNAME24595(G24595,G22916,G22881);
  or GNAME24596(G24596,G24595,G24594,G24593);
  xor GNAME24606(G24606,G24607,G22991);
  xor GNAME24607(G24607,G23066,G22911);
  and GNAME24608(G24608,G23066,G22991);
  and GNAME24609(G24609,G22911,G22991);
  and GNAME24610(G24610,G23066,G22911);
  or GNAME24611(G24611,G24610,G24609,G24608);
  xor GNAME24621(G24621,G24622,G23006);
  xor GNAME24622(G24622,G22931,G22896);
  and GNAME24623(G24623,G22931,G23006);
  and GNAME24624(G24624,G22896,G23006);
  and GNAME24625(G24625,G22931,G22896);
  or GNAME24626(G24626,G24625,G24624,G24623);
  xor GNAME24636(G24636,G24637,G23021);
  xor GNAME24637(G24637,G23081,G22926);
  and GNAME24638(G24638,G23081,G23021);
  and GNAME24639(G24639,G22926,G23021);
  and GNAME24640(G24640,G23081,G22926);
  or GNAME24641(G24641,G24640,G24639,G24638);
  xor GNAME24651(G24651,G24652,G24561);
  xor GNAME24652(G24652,G22776,G24581);
  and GNAME24653(G24653,G22776,G24561);
  and GNAME24654(G24654,G24581,G24561);
  and GNAME24655(G24655,G22776,G24581);
  or GNAME24656(G24656,G24655,G24654,G24653);
  xor GNAME24666(G24666,G24667,G24576);
  xor GNAME24667(G24667,G22941,G24746);
  and GNAME24668(G24668,G22941,G24576);
  and GNAME24669(G24669,G24746,G24576);
  and GNAME24670(G24670,G22941,G24746);
  or GNAME24671(G24671,G24670,G24669,G24668);
  xor GNAME24681(G24681,G24682,G24591);
  xor GNAME24682(G24682,G22806,G24611);
  and GNAME24683(G24683,G22806,G24591);
  and GNAME24684(G24684,G24611,G24591);
  and GNAME24685(G24685,G22806,G24611);
  or GNAME24686(G24686,G24685,G24684,G24683);
  xor GNAME24696(G24696,G24697,G24621);
  xor GNAME24697(G24697,G22836,G24641);
  and GNAME24698(G24698,G22836,G24621);
  and GNAME24699(G24699,G24641,G24621);
  and GNAME24700(G24700,G22836,G24641);
  or GNAME24701(G24701,G24700,G24699,G24698);
  xor GNAME24711(G24711,G24712,G24606);
  xor GNAME24712(G24712,G22971,G24776);
  and GNAME24713(G24713,G22971,G24606);
  and GNAME24714(G24714,G24776,G24606);
  and GNAME24715(G24715,G22971,G24776);
  or GNAME24716(G24716,G24715,G24714,G24713);
  xor GNAME24726(G24726,G24727,G24636);
  xor GNAME24727(G24727,G23001,G24806);
  and GNAME24728(G24728,G23001,G24636);
  and GNAME24729(G24729,G24806,G24636);
  and GNAME24730(G24730,G23001,G24806);
  or GNAME24731(G24731,G24730,G24729,G24728);
  xor GNAME24741(G24741,G24742,G23126);
  xor GNAME24742(G24742,G23051,G23031);
  and GNAME24743(G24743,G23051,G23126);
  and GNAME24744(G24744,G23031,G23126);
  and GNAME24745(G24745,G23051,G23031);
  or GNAME24746(G24746,G24745,G24744,G24743);
  xor GNAME24756(G24756,G24757,G23141);
  xor GNAME24757(G24757,G23306,G23046);
  and GNAME24758(G24758,G23306,G23141);
  and GNAME24759(G24759,G23046,G23141);
  and GNAME24760(G24760,G23306,G23046);
  or GNAME24761(G24761,G24760,G24759,G24758);
  xor GNAME24771(G24771,G24772,G23156);
  xor GNAME24772(G24772,G23096,G23061);
  and GNAME24773(G24773,G23096,G23156);
  and GNAME24774(G24774,G23061,G23156);
  and GNAME24775(G24775,G23096,G23061);
  or GNAME24776(G24776,G24775,G24774,G24773);
  xor GNAME24786(G24786,G24787,G23171);
  xor GNAME24787(G24787,G23321,G23091);
  and GNAME24788(G24788,G23321,G23171);
  and GNAME24789(G24789,G23091,G23171);
  and GNAME24790(G24790,G23321,G23091);
  or GNAME24791(G24791,G24790,G24789,G24788);
  xor GNAME24801(G24801,G24802,G23186);
  xor GNAME24802(G24802,G23111,G23076);
  and GNAME24803(G24803,G23111,G23186);
  and GNAME24804(G24804,G23076,G23186);
  and GNAME24805(G24805,G23111,G23076);
  or GNAME24806(G24806,G24805,G24804,G24803);
  xor GNAME24816(G24816,G24817,G23201);
  xor GNAME24817(G24817,G23336,G23106);
  and GNAME24818(G24818,G23336,G23201);
  and GNAME24819(G24819,G23106,G23201);
  and GNAME24820(G24820,G23336,G23106);
  or GNAME24821(G24821,G24820,G24819,G24818);
  xor GNAME24831(G24831,G24832,G24741);
  xor GNAME24832(G24832,G22956,G24761);
  and GNAME24833(G24833,G22956,G24741);
  and GNAME24834(G24834,G24761,G24741);
  and GNAME24835(G24835,G22956,G24761);
  or GNAME24836(G24836,G24835,G24834,G24833);
  xor GNAME24846(G24846,G24847,G24756);
  xor GNAME24847(G24847,G23121,G23216);
  and GNAME24848(G24848,G23121,G24756);
  and GNAME24849(G24849,G23216,G24756);
  and GNAME24850(G24850,G23121,G23216);
  or GNAME24851(G24851,G24850,G24849,G24848);
  xor GNAME24861(G24861,G24862,G24771);
  xor GNAME24862(G24862,G22986,G24791);
  and GNAME24863(G24863,G22986,G24771);
  and GNAME24864(G24864,G24791,G24771);
  and GNAME24865(G24865,G22986,G24791);
  or GNAME24866(G24866,G24865,G24864,G24863);
  xor GNAME24876(G24876,G24877,G24801);
  xor GNAME24877(G24877,G23016,G24821);
  and GNAME24878(G24878,G23016,G24801);
  and GNAME24879(G24879,G24821,G24801);
  and GNAME24880(G24880,G23016,G24821);
  or GNAME24881(G24881,G24880,G24879,G24878);
  xor GNAME24891(G24891,G24892,G24786);
  xor GNAME24892(G24892,G23151,G23246);
  and GNAME24893(G24893,G23151,G24786);
  and GNAME24894(G24894,G23246,G24786);
  and GNAME24895(G24895,G23151,G23246);
  or GNAME24896(G24896,G24895,G24894,G24893);
  xor GNAME24906(G24906,G24907,G24816);
  xor GNAME24907(G24907,G23181,G23276);
  and GNAME24908(G24908,G23181,G24816);
  and GNAME24909(G24909,G23276,G24816);
  and GNAME24910(G24910,G23181,G23276);
  or GNAME24911(G24911,G24910,G24909,G24908);
  xor GNAME24921(G24921,G24922,G23211);
  xor GNAME24922(G24922,G23136,G23231);
  and GNAME24923(G24923,G23136,G23211);
  and GNAME24924(G24924,G23231,G23211);
  and GNAME24925(G24925,G23136,G23231);
  or GNAME24926(G24926,G24925,G24924,G24923);
  xor GNAME24936(G24936,G24937,G23226);
  xor GNAME24937(G24937,G23346,G23396);
  and GNAME24938(G24938,G23346,G23226);
  and GNAME24939(G24939,G23396,G23226);
  and GNAME24940(G24940,G23346,G23396);
  or GNAME24941(G24941,G24940,G24939,G24938);
  xor GNAME24951(G24951,G24952,G23241);
  xor GNAME24952(G24952,G23166,G23261);
  and GNAME24953(G24953,G23166,G23241);
  and GNAME24954(G24954,G23261,G23241);
  and GNAME24955(G24955,G23166,G23261);
  or GNAME24956(G24956,G24955,G24954,G24953);
  xor GNAME24966(G24966,G24967,G23271);
  xor GNAME24967(G24967,G23196,G23291);
  and GNAME24968(G24968,G23196,G23271);
  and GNAME24969(G24969,G23291,G23271);
  and GNAME24970(G24970,G23196,G23291);
  or GNAME24971(G24971,G24970,G24969,G24968);
  xor GNAME24981(G24981,G24982,G23256);
  xor GNAME24982(G24982,G23361,G23426);
  and GNAME24983(G24983,G23361,G23256);
  and GNAME24984(G24984,G23426,G23256);
  and GNAME24985(G24985,G23361,G23426);
  or GNAME24986(G24986,G24985,G24984,G24983);
  xor GNAME24996(G24996,G24997,G23286);
  xor GNAME24997(G24997,G23376,G23456);
  and GNAME24998(G24998,G23376,G23286);
  and GNAME24999(G24999,G23456,G23286);
  and GNAME25000(G25000,G23376,G23456);
  or GNAME25001(G25001,G25000,G24999,G24998);
  xor GNAME25011(G25011,G25012,G23406);
  xor GNAME25012(G25012,G23526,G23576);
  and GNAME25013(G25013,G23526,G23406);
  and GNAME25014(G25014,G23576,G23406);
  and GNAME25015(G25015,G23526,G23576);
  or GNAME25016(G25016,G25015,G25014,G25013);
  xor GNAME25026(G25026,G25027,G23436);
  xor GNAME25027(G25027,G23541,G23606);
  and GNAME25028(G25028,G23541,G23436);
  and GNAME25029(G25029,G23606,G23436);
  and GNAME25030(G25030,G23541,G23606);
  or GNAME25031(G25031,G25030,G25029,G25028);
  xor GNAME25041(G25041,G25042,G23466);
  xor GNAME25042(G25042,G23556,G23636);
  and GNAME25043(G25043,G23556,G23466);
  and GNAME25044(G25044,G23636,G23466);
  and GNAME25045(G25045,G23556,G23636);
  or GNAME25046(G25046,G25045,G25044,G25043);
  xor GNAME25056(G25056,G25057,G25076);
  xor GNAME25057(G25057,G21861,G21911);
  and GNAME25058(G25058,G21861,G25076);
  and GNAME25059(G25059,G21911,G25076);
  and GNAME25060(G25060,G21861,G21911);
  or GNAME25061(G25061,G25060,G25059,G25058);
  xor GNAME25071(G25071,G25072,G25091);
  xor GNAME25072(G25072,G21906,G22001);
  and GNAME25073(G25073,G21906,G25091);
  and GNAME25074(G25074,G22001,G25091);
  and GNAME25075(G25075,G21906,G22001);
  or GNAME25076(G25076,G25075,G25074,G25073);
  xor GNAME25086(G25086,G25087,G25106);
  xor GNAME25087(G25087,G22016,G21996);
  and GNAME25088(G25088,G22016,G25106);
  and GNAME25089(G25089,G21996,G25106);
  and GNAME25090(G25090,G22016,G21996);
  or GNAME25091(G25091,G25090,G25089,G25088);
  xor GNAME25101(G25101,G25102,G25121);
  xor GNAME25102(G25102,G22181,G22011);
  and GNAME25103(G25103,G22181,G25121);
  and GNAME25104(G25104,G22011,G25121);
  and GNAME25105(G25105,G22181,G22011);
  or GNAME25106(G25106,G25105,G25104,G25103);
  xor GNAME25116(G25116,G25117,G25136);
  xor GNAME25117(G25117,G22196,G22176);
  and GNAME25118(G25118,G22196,G25136);
  and GNAME25119(G25119,G22176,G25136);
  and GNAME25120(G25120,G22196,G22176);
  or GNAME25121(G25121,G25120,G25119,G25118);
  xor GNAME25131(G25131,G25132,G25151);
  xor GNAME25132(G25132,G24206,G22191);
  and GNAME25133(G25133,G24206,G25151);
  and GNAME25134(G25134,G22191,G25151);
  and GNAME25135(G25135,G24206,G22191);
  or GNAME25136(G25136,G25135,G25134,G25133);
  xor GNAME25146(G25146,G25147,G25166);
  xor GNAME25147(G25147,G22406,G24201);
  and GNAME25148(G25148,G22406,G25166);
  and GNAME25149(G25149,G24201,G25166);
  and GNAME25150(G25150,G22406,G24201);
  or GNAME25151(G25151,G25150,G25149,G25148);
  xor GNAME25161(G25161,G25162,G25181);
  xor GNAME25162(G25162,G22496,G22401);
  and GNAME25163(G25163,G22496,G25181);
  and GNAME25164(G25164,G22401,G25181);
  and GNAME25165(G25165,G22496,G22401);
  or GNAME25166(G25166,G25165,G25164,G25163);
  xor GNAME25176(G25176,G25177,G25826);
  xor GNAME25177(G25177,G24341,G22491);
  and GNAME25178(G25178,G24341,G25826);
  and GNAME25179(G25179,G22491,G25826);
  and GNAME25180(G25180,G24341,G22491);
  or GNAME25181(G25181,G25180,G25179,G25178);
  xor GNAME25191(G25191,G25192,G25211);
  xor GNAME25192(G25192,G21876,G21926);
  and GNAME25193(G25193,G21876,G25211);
  and GNAME25194(G25194,G21926,G25211);
  and GNAME25195(G25195,G21876,G21926);
  or GNAME25196(G25196,G25195,G25194,G25193);
  xor GNAME25206(G25206,G25207,G25256);
  xor GNAME25207(G25207,G21921,G22031);
  and GNAME25208(G25208,G21921,G25256);
  and GNAME25209(G25209,G22031,G25256);
  and GNAME25210(G25210,G21921,G22031);
  or GNAME25211(G25211,G25210,G25209,G25208);
  xor GNAME25221(G25221,G25222,G25241);
  xor GNAME25222(G25222,G21891,G21941);
  and GNAME25223(G25223,G21891,G25241);
  and GNAME25224(G25224,G21941,G25241);
  and GNAME25225(G25225,G21891,G21941);
  or GNAME25226(G25226,G25225,G25224,G25223);
  xor GNAME25236(G25236,G25237,G25301);
  xor GNAME25237(G25237,G21936,G22046);
  and GNAME25238(G25238,G21936,G25301);
  and GNAME25239(G25239,G22046,G25301);
  and GNAME25240(G25240,G21936,G22046);
  or GNAME25241(G25241,G25240,G25239,G25238);
  xor GNAME25251(G25251,G25252,G25271);
  xor GNAME25252(G25252,G22061,G22026);
  and GNAME25253(G25253,G22061,G25271);
  and GNAME25254(G25254,G22026,G25271);
  and GNAME25255(G25255,G22061,G22026);
  or GNAME25256(G25256,G25255,G25254,G25253);
  xor GNAME25266(G25266,G25267,G25331);
  xor GNAME25267(G25267,G22211,G22056);
  and GNAME25268(G25268,G22211,G25331);
  and GNAME25269(G25269,G22056,G25331);
  and GNAME25270(G25270,G22211,G22056);
  or GNAME25271(G25271,G25270,G25269,G25268);
  xor GNAME25281(G25281,G25282,G25361);
  xor GNAME25282(G25282,G23486,G24936);
  and GNAME25283(G25283,G23486,G25361);
  and GNAME25284(G25284,G24936,G25361);
  and GNAME25285(G25285,G23486,G24936);
  or GNAME25286(G25286,G25285,G25284,G25283);
  xor GNAME25296(G25296,G25297,G25316);
  xor GNAME25297(G25297,G22076,G22041);
  and GNAME25298(G25298,G22076,G25316);
  and GNAME25299(G25299,G22041,G25316);
  and GNAME25300(G25300,G22076,G22041);
  or GNAME25301(G25301,G25300,G25299,G25298);
  xor GNAME25311(G25311,G25312,G25421);
  xor GNAME25312(G25312,G22226,G22071);
  and GNAME25313(G25313,G22226,G25421);
  and GNAME25314(G25314,G22071,G25421);
  and GNAME25315(G25315,G22226,G22071);
  or GNAME25316(G25316,G25315,G25314,G25313);
  xor GNAME25326(G25326,G25327,G25346);
  xor GNAME25327(G25327,G22241,G22206);
  and GNAME25328(G25328,G22241,G25346);
  and GNAME25329(G25329,G22206,G25346);
  and GNAME25330(G25330,G22241,G22206);
  or GNAME25331(G25331,G25330,G25329,G25328);
  xor GNAME25341(G25341,G25342,G25451);
  xor GNAME25342(G25342,G24221,G22236);
  and GNAME25343(G25343,G24221,G25451);
  and GNAME25344(G25344,G22236,G25451);
  and GNAME25345(G25345,G24221,G22236);
  or GNAME25346(G25346,G25345,G25344,G25343);
  xor GNAME25356(G25356,G25357,G25376);
  xor GNAME25357(G25357,G25016,G23481);
  and GNAME25358(G25358,G25016,G25376);
  and GNAME25359(G25359,G23481,G25376);
  and GNAME25360(G25360,G25016,G23481);
  or GNAME25361(G25361,G25360,G25359,G25358);
  xor GNAME25371(G25371,G25372,G25391);
  xor GNAME25372(G25372,G23666,G25011);
  and GNAME25373(G25373,G23666,G25391);
  and GNAME25374(G25374,G25011,G25391);
  and GNAME25375(G25375,G23666,G25011);
  or GNAME25376(G25376,G25375,G25374,G25373);
  xor GNAME25386(G25386,G25387,G25406);
  xor GNAME25387(G25387,G23681,G23661);
  and GNAME25388(G25388,G23681,G25406);
  and GNAME25389(G25389,G23661,G25406);
  and GNAME25390(G25390,G23681,G23661);
  or GNAME25391(G25391,G25390,G25389,G25388);
  xor GNAME25401(G25401,G25402,G25481);
  xor GNAME25402(G25402,G23696,G23676);
  and GNAME25403(G25403,G23696,G25481);
  and GNAME25404(G25404,G23676,G25481);
  and GNAME25405(G25405,G23696,G23676);
  or GNAME25406(G25406,G25405,G25404,G25403);
  xor GNAME25416(G25416,G25417,G25436);
  xor GNAME25417(G25417,G22256,G22221);
  and GNAME25418(G25418,G22256,G25436);
  and GNAME25419(G25419,G22221,G25436);
  and GNAME25420(G25420,G22256,G22221);
  or GNAME25421(G25421,G25420,G25419,G25418);
  xor GNAME25431(G25431,G25432,G25526);
  xor GNAME25432(G25432,G24236,G22251);
  and GNAME25433(G25433,G24236,G25526);
  and GNAME25434(G25434,G22251,G25526);
  and GNAME25435(G25435,G24236,G22251);
  or GNAME25436(G25436,G25435,G25434,G25433);
  xor GNAME25446(G25446,G25447,G25466);
  xor GNAME25447(G25447,G22421,G24216);
  and GNAME25448(G25448,G22421,G25466);
  and GNAME25449(G25449,G24216,G25466);
  and GNAME25450(G25450,G22421,G24216);
  or GNAME25451(G25451,G25450,G25449,G25448);
  xor GNAME25461(G25461,G25462,G25556);
  xor GNAME25462(G25462,G22511,G22416);
  and GNAME25463(G25463,G22511,G25556);
  and GNAME25464(G25464,G22416,G25556);
  and GNAME25465(G25465,G22511,G22416);
  or GNAME25466(G25466,G25465,G25464,G25463);
  xor GNAME25476(G25476,G25477,G25496);
  xor GNAME25477(G25477,G23801,G23691);
  and GNAME25478(G25478,G23801,G25496);
  and GNAME25479(G25479,G23691,G25496);
  and GNAME25480(G25480,G23801,G23691);
  or GNAME25481(G25481,G25480,G25479,G25478);
  xor GNAME25491(G25491,G25492,G25511);
  xor GNAME25492(G25492,G23816,G23796);
  and GNAME25493(G25493,G23816,G25511);
  and GNAME25494(G25494,G23796,G25511);
  and GNAME25495(G25495,G23816,G23796);
  or GNAME25496(G25496,G25495,G25494,G25493);
  xor GNAME25506(G25506,G25507,G24071);
  xor GNAME25507(G25507,G23891,G23811);
  and GNAME25508(G25508,G23891,G24071);
  and GNAME25509(G25509,G23811,G24071);
  and GNAME25510(G25510,G23891,G23811);
  or GNAME25511(G25511,G25510,G25509,G25508);
  xor GNAME25521(G25521,G25522,G25541);
  xor GNAME25522(G25522,G22436,G24231);
  and GNAME25523(G25523,G22436,G25541);
  and GNAME25524(G25524,G24231,G25541);
  and GNAME25525(G25525,G22436,G24231);
  or GNAME25526(G25526,G25525,G25524,G25523);
  xor GNAME25536(G25536,G25537,G25571);
  xor GNAME25537(G25537,G22526,G22431);
  and GNAME25538(G25538,G22526,G25571);
  and GNAME25539(G25539,G22431,G25571);
  and GNAME25540(G25540,G22526,G22431);
  or GNAME25541(G25541,G25540,G25539,G25538);
  xor GNAME25551(G25551,G25552,G25946);
  xor GNAME25552(G25552,G24356,G22506);
  and GNAME25553(G25553,G24356,G25946);
  and GNAME25554(G25554,G22506,G25946);
  and GNAME25555(G25555,G24356,G22506);
  or GNAME25556(G25556,G25555,G25554,G25553);
  xor GNAME25566(G25566,G25567,G25961);
  xor GNAME25567(G25567,G24371,G22521);
  and GNAME25568(G25568,G24371,G25961);
  and GNAME25569(G25569,G22521,G25961);
  and GNAME25570(G25570,G24371,G22521);
  or GNAME25571(G25571,G25570,G25569,G25568);
  xor GNAME25581(G25581,G25582,G25616);
  xor GNAME25582(G25582,G23501,G24981);
  and GNAME25583(G25583,G23501,G25616);
  and GNAME25584(G25584,G24981,G25616);
  and GNAME25585(G25585,G23501,G24981);
  or GNAME25586(G25586,G25585,G25584,G25583);
  xor GNAME25596(G25596,G25597,G25646);
  xor GNAME25597(G25597,G23516,G24996);
  and GNAME25598(G25598,G23516,G25646);
  and GNAME25599(G25599,G24996,G25646);
  and GNAME25600(G25600,G23516,G24996);
  or GNAME25601(G25601,G25600,G25599,G25598);
  xor GNAME25611(G25611,G25612,G25631);
  xor GNAME25612(G25612,G25031,G23496);
  and GNAME25613(G25613,G25031,G25631);
  and GNAME25614(G25614,G23496,G25631);
  and GNAME25615(G25615,G25031,G23496);
  or GNAME25616(G25616,G25615,G25614,G25613);
  xor GNAME25626(G25626,G25627,G25676);
  xor GNAME25627(G25627,G23711,G25026);
  and GNAME25628(G25628,G23711,G25676);
  and GNAME25629(G25629,G25026,G25676);
  and GNAME25630(G25630,G23711,G25026);
  or GNAME25631(G25631,G25630,G25629,G25628);
  xor GNAME25641(G25641,G25642,G25661);
  xor GNAME25642(G25642,G25046,G23511);
  and GNAME25643(G25643,G25046,G25661);
  and GNAME25644(G25644,G23511,G25661);
  and GNAME25645(G25645,G25046,G23511);
  or GNAME25646(G25646,G25645,G25644,G25643);
  xor GNAME25656(G25656,G25657,G25706);
  xor GNAME25657(G25657,G23726,G25041);
  and GNAME25658(G25658,G23726,G25706);
  and GNAME25659(G25659,G25041,G25706);
  and GNAME25660(G25660,G23726,G25041);
  or GNAME25661(G25661,G25660,G25659,G25658);
  xor GNAME25671(G25671,G25672,G25691);
  xor GNAME25672(G25672,G23741,G23706);
  and GNAME25673(G25673,G23741,G25691);
  and GNAME25674(G25674,G23706,G25691);
  and GNAME25675(G25675,G23741,G23706);
  or GNAME25676(G25676,G25675,G25674,G25673);
  xor GNAME25686(G25686,G25687,G25736);
  xor GNAME25687(G25687,G23756,G23736);
  and GNAME25688(G25688,G23756,G25736);
  and GNAME25689(G25689,G23736,G25736);
  and GNAME25690(G25690,G23756,G23736);
  or GNAME25691(G25691,G25690,G25689,G25688);
  xor GNAME25701(G25701,G25702,G25721);
  xor GNAME25702(G25702,G23771,G23721);
  and GNAME25703(G25703,G23771,G25721);
  and GNAME25704(G25704,G23721,G25721);
  and GNAME25705(G25705,G23771,G23721);
  or GNAME25706(G25706,G25705,G25704,G25703);
  xor GNAME25716(G25716,G25717,G25766);
  xor GNAME25717(G25717,G23786,G23766);
  and GNAME25718(G25718,G23786,G25766);
  and GNAME25719(G25719,G23766,G25766);
  and GNAME25720(G25720,G23786,G23766);
  or GNAME25721(G25721,G25720,G25719,G25718);
  xor GNAME25731(G25731,G25732,G25751);
  xor GNAME25732(G25732,G23831,G23751);
  and GNAME25733(G25733,G23831,G25751);
  and GNAME25734(G25734,G23751,G25751);
  and GNAME25735(G25735,G23831,G23751);
  or GNAME25736(G25736,G25735,G25734,G25733);
  xor GNAME25746(G25746,G25747,G25796);
  xor GNAME25747(G25747,G23846,G23826);
  and GNAME25748(G25748,G23846,G25796);
  and GNAME25749(G25749,G23826,G25796);
  and GNAME25750(G25750,G23846,G23826);
  or GNAME25751(G25751,G25750,G25749,G25748);
  xor GNAME25761(G25761,G25762,G25781);
  xor GNAME25762(G25762,G23861,G23781);
  and GNAME25763(G25763,G23861,G25781);
  and GNAME25764(G25764,G23781,G25781);
  and GNAME25765(G25765,G23861,G23781);
  or GNAME25766(G25766,G25765,G25764,G25763);
  xor GNAME25776(G25776,G25777,G25811);
  xor GNAME25777(G25777,G23876,G23856);
  and GNAME25778(G25778,G23876,G25811);
  and GNAME25779(G25779,G23856,G25811);
  and GNAME25780(G25780,G23876,G23856);
  or GNAME25781(G25781,G25780,G25779,G25778);
  xor GNAME25791(G25791,G25792,G24101);
  xor GNAME25792(G25792,G23906,G23841);
  and GNAME25793(G25793,G23906,G24101);
  and GNAME25794(G25794,G23841,G24101);
  and GNAME25795(G25795,G23906,G23841);
  or GNAME25796(G25796,G25795,G25794,G25793);
  xor GNAME25806(G25806,G25807,G24116);
  xor GNAME25807(G25807,G23921,G23871);
  and GNAME25808(G25808,G23921,G24116);
  and GNAME25809(G25809,G23871,G24116);
  and GNAME25810(G25810,G23921,G23871);
  or GNAME25811(G25811,G25810,G25809,G25808);
  xor GNAME25821(G25821,G25822,G25841);
  xor GNAME25822(G25822,G24476,G24336);
  and GNAME25823(G25823,G24476,G25841);
  and GNAME25824(G25824,G24336,G25841);
  and GNAME25825(G25825,G24476,G24336);
  or GNAME25826(G25826,G25825,G25824,G25823);
  xor GNAME25836(G25836,G25837,G25856);
  xor GNAME25837(G25837,G24491,G24471);
  and GNAME25838(G25838,G24491,G25856);
  and GNAME25839(G25839,G24471,G25856);
  and GNAME25840(G25840,G24491,G24471);
  or GNAME25841(G25841,G25840,G25839,G25838);
  xor GNAME25851(G25851,G25852,G25871);
  xor GNAME25852(G25852,G24656,G24486);
  and GNAME25853(G25853,G24656,G25871);
  and GNAME25854(G25854,G24486,G25871);
  and GNAME25855(G25855,G24656,G24486);
  or GNAME25856(G25856,G25855,G25854,G25853);
  xor GNAME25866(G25866,G25867,G25886);
  xor GNAME25867(G25867,G24671,G24651);
  and GNAME25868(G25868,G24671,G25886);
  and GNAME25869(G25869,G24651,G25886);
  and GNAME25870(G25870,G24671,G24651);
  or GNAME25871(G25871,G25870,G25869,G25868);
  xor GNAME25881(G25881,G25882,G25901);
  xor GNAME25882(G25882,G24836,G24666);
  and GNAME25883(G25883,G24836,G25901);
  and GNAME25884(G25884,G24666,G25901);
  and GNAME25885(G25885,G24836,G24666);
  or GNAME25886(G25886,G25885,G25884,G25883);
  xor GNAME25896(G25896,G25897,G25916);
  xor GNAME25897(G25897,G24851,G24831);
  and GNAME25898(G25898,G24851,G25916);
  and GNAME25899(G25899,G24831,G25916);
  and GNAME25900(G25900,G24851,G24831);
  or GNAME25901(G25901,G25900,G25899,G25898);
  xor GNAME25911(G25911,G25912,G25931);
  xor GNAME25912(G25912,G24926,G24846);
  and GNAME25913(G25913,G24926,G25931);
  and GNAME25914(G25914,G24846,G25931);
  and GNAME25915(G25915,G24926,G24846);
  or GNAME25916(G25916,G25915,G25914,G25913);
  xor GNAME25926(G25926,G25927,G25286);
  xor GNAME25927(G25927,G24941,G24921);
  and GNAME25928(G25928,G24941,G25286);
  and GNAME25929(G25929,G24921,G25286);
  and GNAME25930(G25930,G24941,G24921);
  or GNAME25931(G25931,G25930,G25929,G25928);
  xor GNAME25941(G25941,G25942,G25976);
  xor GNAME25942(G25942,G24506,G24351);
  and GNAME25943(G25943,G24506,G25976);
  and GNAME25944(G25944,G24351,G25976);
  and GNAME25945(G25945,G24506,G24351);
  or GNAME25946(G25946,G25945,G25944,G25943);
  xor GNAME25956(G25956,G25957,G26006);
  xor GNAME25957(G25957,G24521,G24366);
  and GNAME25958(G25958,G24521,G26006);
  and GNAME25959(G25959,G24366,G26006);
  and GNAME25960(G25960,G24521,G24366);
  or GNAME25961(G25961,G25960,G25959,G25958);
  xor GNAME25971(G25971,G25972,G25991);
  xor GNAME25972(G25972,G24536,G24501);
  and GNAME25973(G25973,G24536,G25991);
  and GNAME25974(G25974,G24501,G25991);
  and GNAME25975(G25975,G24536,G24501);
  or GNAME25976(G25976,G25975,G25974,G25973);
  xor GNAME25986(G25986,G25987,G26036);
  xor GNAME25987(G25987,G24686,G24531);
  and GNAME25988(G25988,G24686,G26036);
  and GNAME25989(G25989,G24531,G26036);
  and GNAME25990(G25990,G24686,G24531);
  or GNAME25991(G25991,G25990,G25989,G25988);
  xor GNAME26001(G26001,G26002,G26021);
  xor GNAME26002(G26002,G24551,G24516);
  and GNAME26003(G26003,G24551,G26021);
  and GNAME26004(G26004,G24516,G26021);
  and GNAME26005(G26005,G24551,G24516);
  or GNAME26006(G26006,G26005,G26004,G26003);
  xor GNAME26016(G26016,G26017,G26066);
  xor GNAME26017(G26017,G24701,G24546);
  and GNAME26018(G26018,G24701,G26066);
  and GNAME26019(G26019,G24546,G26066);
  and GNAME26020(G26020,G24701,G24546);
  or GNAME26021(G26021,G26020,G26019,G26018);
  xor GNAME26031(G26031,G26032,G26051);
  xor GNAME26032(G26032,G24716,G24681);
  and GNAME26033(G26033,G24716,G26051);
  and GNAME26034(G26034,G24681,G26051);
  and GNAME26035(G26035,G24716,G24681);
  or GNAME26036(G26036,G26035,G26034,G26033);
  xor GNAME26046(G26046,G26047,G26096);
  xor GNAME26047(G26047,G24866,G24711);
  and GNAME26048(G26048,G24866,G26096);
  and GNAME26049(G26049,G24711,G26096);
  and GNAME26050(G26050,G24866,G24711);
  or GNAME26051(G26051,G26050,G26049,G26048);
  xor GNAME26061(G26061,G26062,G26081);
  xor GNAME26062(G26062,G24731,G24696);
  and GNAME26063(G26063,G24731,G26081);
  and GNAME26064(G26064,G24696,G26081);
  and GNAME26065(G26065,G24731,G24696);
  or GNAME26066(G26066,G26065,G26064,G26063);
  xor GNAME26076(G26076,G26077,G26126);
  xor GNAME26077(G26077,G24881,G24726);
  and GNAME26078(G26078,G24881,G26126);
  and GNAME26079(G26079,G24726,G26126);
  and GNAME26080(G26080,G24881,G24726);
  or GNAME26081(G26081,G26080,G26079,G26078);
  xor GNAME26091(G26091,G26092,G26111);
  xor GNAME26092(G26092,G24896,G24861);
  and GNAME26093(G26093,G24896,G26111);
  and GNAME26094(G26094,G24861,G26111);
  and GNAME26095(G26095,G24896,G24861);
  or GNAME26096(G26096,G26095,G26094,G26093);
  xor GNAME26106(G26106,G26107,G26156);
  xor GNAME26107(G26107,G24956,G24891);
  and GNAME26108(G26108,G24956,G26156);
  and GNAME26109(G26109,G24891,G26156);
  and GNAME26110(G26110,G24956,G24891);
  or GNAME26111(G26111,G26110,G26109,G26108);
  xor GNAME26121(G26121,G26122,G26141);
  xor GNAME26122(G26122,G24911,G24876);
  and GNAME26123(G26123,G24911,G26141);
  and GNAME26124(G26124,G24876,G26141);
  and GNAME26125(G26125,G24911,G24876);
  or GNAME26126(G26126,G26125,G26124,G26123);
  xor GNAME26136(G26136,G26137,G26171);
  xor GNAME26137(G26137,G24971,G24906);
  and GNAME26138(G26138,G24971,G26171);
  and GNAME26139(G26139,G24906,G26171);
  and GNAME26140(G26140,G24971,G24906);
  or GNAME26141(G26141,G26140,G26139,G26138);
  xor GNAME26151(G26151,G26152,G25586);
  xor GNAME26152(G26152,G24986,G24951);
  and GNAME26153(G26153,G24986,G25586);
  and GNAME26154(G26154,G24951,G25586);
  and GNAME26155(G26155,G24986,G24951);
  or GNAME26156(G26156,G26155,G26154,G26153);
  xor GNAME26166(G26166,G26167,G25601);
  xor GNAME26167(G26167,G25001,G24966);
  and GNAME26168(G26168,G25001,G25601);
  and GNAME26169(G26169,G24966,G25601);
  and GNAME26170(G26170,G25001,G24966);
  or GNAME26171(G26171,G26170,G26169,G26168);
  xor GNAME26181(G26181,G26182,G26681);
  xor GNAME26182(G26182,G33942,G3531);
  and GNAME26183(G26183,G33942,G26681);
  and GNAME26184(G26184,G3531,G26681);
  and GNAME26185(G26185,G33942,G3531);
  or GNAME26186(G26186,G26185,G26184,G26183);
  xor GNAME26196(G26196,G26197,G27506);
  xor GNAME26197(G26197,G34436,G34462);
  and GNAME26198(G26198,G34436,G27506);
  and GNAME26199(G26199,G34462,G27506);
  and GNAME26200(G26200,G34436,G34462);
  or GNAME26201(G26201,G26200,G26199,G26198);
  xor GNAME26211(G26211,G26212,G27569);
  xor GNAME26212(G26212,G31771,G2781);
  and GNAME26213(G26213,G31771,G27569);
  and GNAME26214(G26214,G2781,G27569);
  and GNAME26215(G26215,G31771,G2781);
  or GNAME26216(G26216,G26215,G26214,G26213);
  xor GNAME26226(G26226,G26227,G27568);
  xor GNAME26227(G26227,G31797,G31810);
  and GNAME26228(G26228,G31797,G27568);
  and GNAME26229(G26229,G31810,G27568);
  and GNAME26230(G26230,G31797,G31810);
  or GNAME26231(G26231,G26230,G26229,G26228);
  xor GNAME26241(G26241,G26242,G27567);
  xor GNAME26242(G26242,G27851,G27854);
  and GNAME26243(G26243,G27851,G27567);
  and GNAME26244(G26244,G27854,G27567);
  and GNAME26245(G26245,G27851,G27854);
  or GNAME26246(G26246,G26245,G26244,G26243);
  xor GNAME26256(G26256,G26257,G26216);
  xor GNAME26257(G26257,G31784,G2802);
  and GNAME26258(G26258,G31784,G26216);
  and GNAME26259(G26259,G2802,G26216);
  and GNAME26260(G26260,G31784,G2802);
  or GNAME26261(G26261,G26260,G26259,G26258);
  xor GNAME26271(G26271,G26272,G26261);
  xor GNAME26272(G26272,G31875,G2823);
  and GNAME26273(G26273,G31875,G26261);
  and GNAME26274(G26274,G2823,G26261);
  and GNAME26275(G26275,G31875,G2823);
  or GNAME26276(G26276,G26275,G26274,G26273);
  xor GNAME26286(G26286,G26287,G26276);
  xor GNAME26287(G26287,G31888,G2844);
  and GNAME26288(G26288,G31888,G26276);
  and GNAME26289(G26289,G2844,G26276);
  and GNAME26290(G26290,G31888,G2844);
  or GNAME26291(G26291,G26290,G26289,G26288);
  xor GNAME26301(G26301,G26302,G26291);
  xor GNAME26302(G26302,G32005,G2865);
  and GNAME26303(G26303,G32005,G26291);
  and GNAME26304(G26304,G2865,G26291);
  and GNAME26305(G26305,G32005,G2865);
  or GNAME26306(G26306,G26305,G26304,G26303);
  xor GNAME26316(G26316,G26317,G26306);
  xor GNAME26317(G26317,G32018,G2886);
  and GNAME26318(G26318,G32018,G26306);
  and GNAME26319(G26319,G2886,G26306);
  and GNAME26320(G26320,G32018,G2886);
  or GNAME26321(G26321,G26320,G26319,G26318);
  xor GNAME26331(G26331,G26332,G26321);
  xor GNAME26332(G26332,G32135,G2907);
  and GNAME26333(G26333,G32135,G26321);
  and GNAME26334(G26334,G2907,G26321);
  and GNAME26335(G26335,G32135,G2907);
  or GNAME26336(G26336,G26335,G26334,G26333);
  xor GNAME26346(G26346,G26347,G26336);
  xor GNAME26347(G26347,G32148,G2968);
  and GNAME26348(G26348,G32148,G26336);
  and GNAME26349(G26349,G2968,G26336);
  and GNAME26350(G26350,G32148,G2968);
  or GNAME26351(G26351,G26350,G26349,G26348);
  xor GNAME26361(G26361,G26362,G26351);
  xor GNAME26362(G26362,G32265,G2989);
  and GNAME26363(G26363,G32265,G26351);
  and GNAME26364(G26364,G2989,G26351);
  and GNAME26365(G26365,G32265,G2989);
  or GNAME26366(G26366,G26365,G26364,G26363);
  xor GNAME26376(G26376,G26377,G26366);
  xor GNAME26377(G26377,G32278,G3010);
  and GNAME26378(G26378,G32278,G26366);
  and GNAME26379(G26379,G3010,G26366);
  and GNAME26380(G26380,G32278,G3010);
  or GNAME26381(G26381,G26380,G26379,G26378);
  xor GNAME26391(G26391,G26392,G26381);
  xor GNAME26392(G26392,G32395,G3031);
  and GNAME26393(G26393,G32395,G26381);
  and GNAME26394(G26394,G3031,G26381);
  and GNAME26395(G26395,G32395,G3031);
  or GNAME26396(G26396,G26395,G26394,G26393);
  xor GNAME26406(G26406,G26407,G26396);
  xor GNAME26407(G26407,G32408,G3052);
  and GNAME26408(G26408,G32408,G26396);
  and GNAME26409(G26409,G3052,G26396);
  and GNAME26410(G26410,G32408,G3052);
  or GNAME26411(G26411,G26410,G26409,G26408);
  xor GNAME26421(G26421,G26422,G26411);
  xor GNAME26422(G26422,G32525,G3073);
  and GNAME26423(G26423,G32525,G26411);
  and GNAME26424(G26424,G3073,G26411);
  and GNAME26425(G26425,G32525,G3073);
  or GNAME26426(G26426,G26425,G26424,G26423);
  xor GNAME26436(G26436,G26437,G26426);
  xor GNAME26437(G26437,G32538,G3094);
  and GNAME26438(G26438,G32538,G26426);
  and GNAME26439(G26439,G3094,G26426);
  and GNAME26440(G26440,G32538,G3094);
  or GNAME26441(G26441,G26440,G26439,G26438);
  xor GNAME26451(G26451,G26452,G26441);
  xor GNAME26452(G26452,G32655,G3115);
  and GNAME26453(G26453,G32655,G26441);
  and GNAME26454(G26454,G3115,G26441);
  and GNAME26455(G26455,G32655,G3115);
  or GNAME26456(G26456,G26455,G26454,G26453);
  xor GNAME26466(G26466,G26467,G26456);
  xor GNAME26467(G26467,G32668,G3176);
  and GNAME26468(G26468,G32668,G26456);
  and GNAME26469(G26469,G3176,G26456);
  and GNAME26470(G26470,G32668,G3176);
  or GNAME26471(G26471,G26470,G26469,G26468);
  xor GNAME26481(G26481,G26482,G26471);
  xor GNAME26482(G26482,G32785,G3197);
  and GNAME26483(G26483,G32785,G26471);
  and GNAME26484(G26484,G3197,G26471);
  and GNAME26485(G26485,G32785,G3197);
  or GNAME26486(G26486,G26485,G26484,G26483);
  xor GNAME26496(G26496,G26497,G26486);
  xor GNAME26497(G26497,G32798,G3218);
  and GNAME26498(G26498,G32798,G26486);
  and GNAME26499(G26499,G3218,G26486);
  and GNAME26500(G26500,G32798,G3218);
  or GNAME26501(G26501,G26500,G26499,G26498);
  xor GNAME26511(G26511,G26512,G26501);
  xor GNAME26512(G26512,G32980,G3239);
  and GNAME26513(G26513,G32980,G26501);
  and GNAME26514(G26514,G3239,G26501);
  and GNAME26515(G26515,G32980,G3239);
  or GNAME26516(G26516,G26515,G26514,G26513);
  xor GNAME26526(G26526,G26527,G26516);
  xor GNAME26527(G26527,G32993,G3260);
  and GNAME26528(G26528,G32993,G26516);
  and GNAME26529(G26529,G3260,G26516);
  and GNAME26530(G26530,G32993,G3260);
  or GNAME26531(G26531,G26530,G26529,G26528);
  xor GNAME26541(G26541,G26542,G26531);
  xor GNAME26542(G26542,G33162,G3281);
  and GNAME26543(G26543,G33162,G26531);
  and GNAME26544(G26544,G3281,G26531);
  and GNAME26545(G26545,G33162,G3281);
  or GNAME26546(G26546,G26545,G26544,G26543);
  xor GNAME26556(G26556,G26557,G26546);
  xor GNAME26557(G26557,G33175,G3302);
  and GNAME26558(G26558,G33175,G26546);
  and GNAME26559(G26559,G3302,G26546);
  and GNAME26560(G26560,G33175,G3302);
  or GNAME26561(G26561,G26560,G26559,G26558);
  xor GNAME26571(G26571,G26572,G26561);
  xor GNAME26572(G26572,G33188,G3323);
  and GNAME26573(G26573,G33188,G26561);
  and GNAME26574(G26574,G3323,G26561);
  and GNAME26575(G26575,G33188,G3323);
  or GNAME26576(G26576,G26575,G26574,G26573);
  xor GNAME26586(G26586,G26587,G26576);
  xor GNAME26587(G26587,G33370,G3384);
  and GNAME26588(G26588,G33370,G26576);
  and GNAME26589(G26589,G3384,G26576);
  and GNAME26590(G26590,G33370,G3384);
  or GNAME26591(G26591,G26590,G26589,G26588);
  xor GNAME26601(G26601,G26602,G26591);
  xor GNAME26602(G26602,G33383,G3405);
  and GNAME26603(G26603,G33383,G26591);
  and GNAME26604(G26604,G3405,G26591);
  and GNAME26605(G26605,G33383,G3405);
  or GNAME26606(G26606,G26605,G26604,G26603);
  xor GNAME26616(G26616,G26617,G26606);
  xor GNAME26617(G26617,G33552,G3426);
  and GNAME26618(G26618,G33552,G26606);
  and GNAME26619(G26619,G3426,G26606);
  and GNAME26620(G26620,G33552,G3426);
  or GNAME26621(G26621,G26620,G26619,G26618);
  xor GNAME26631(G26631,G26632,G26621);
  xor GNAME26632(G26632,G33565,G3447);
  and GNAME26633(G26633,G33565,G26621);
  and GNAME26634(G26634,G3447,G26621);
  and GNAME26635(G26635,G33565,G3447);
  or GNAME26636(G26636,G26635,G26634,G26633);
  xor GNAME26646(G26646,G26647,G26636);
  xor GNAME26647(G26647,G33747,G3468);
  and GNAME26648(G26648,G33747,G26636);
  and GNAME26649(G26649,G3468,G26636);
  and GNAME26650(G26650,G33747,G3468);
  or GNAME26651(G26651,G26650,G26649,G26648);
  xor GNAME26661(G26661,G26662,G26651);
  xor GNAME26662(G26662,G33760,G3489);
  and GNAME26663(G26663,G33760,G26651);
  and GNAME26664(G26664,G3489,G26651);
  and GNAME26665(G26665,G33760,G3489);
  or GNAME26666(G26666,G26665,G26664,G26663);
  xor GNAME26676(G26676,G26677,G26666);
  xor GNAME26677(G26677,G33929,G3510);
  and GNAME26678(G26678,G33929,G26666);
  and GNAME26679(G26679,G3510,G26666);
  and GNAME26680(G26680,G33929,G3510);
  or GNAME26681(G26681,G26680,G26679,G26678);
  xor GNAME26691(G26691,G26692,G26231);
  xor GNAME26692(G26692,G31901,G31927);
  and GNAME26693(G26693,G31901,G26231);
  and GNAME26694(G26694,G31927,G26231);
  and GNAME26695(G26695,G31901,G31927);
  or GNAME26696(G26696,G26695,G26694,G26693);
  xor GNAME26706(G26706,G26707,G26696);
  xor GNAME26707(G26707,G31914,G31940);
  and GNAME26708(G26708,G31914,G26696);
  and GNAME26709(G26709,G31940,G26696);
  and GNAME26710(G26710,G31914,G31940);
  or GNAME26711(G26711,G26710,G26709,G26708);
  xor GNAME26721(G26721,G26722,G26711);
  xor GNAME26722(G26722,G32031,G32057);
  and GNAME26723(G26723,G32031,G26711);
  and GNAME26724(G26724,G32057,G26711);
  and GNAME26725(G26725,G32031,G32057);
  or GNAME26726(G26726,G26725,G26724,G26723);
  xor GNAME26736(G26736,G26737,G26246);
  xor GNAME26737(G26737,G27845,G27848);
  and GNAME26738(G26738,G27845,G26246);
  and GNAME26739(G26739,G27848,G26246);
  and GNAME26740(G26740,G27845,G27848);
  or GNAME26741(G26741,G26740,G26739,G26738);
  xor GNAME26751(G26751,G26752,G26726);
  xor GNAME26752(G26752,G32044,G32070);
  and GNAME26753(G26753,G32044,G26726);
  and GNAME26754(G26754,G32070,G26726);
  and GNAME26755(G26755,G32044,G32070);
  or GNAME26756(G26756,G26755,G26754,G26753);
  xor GNAME26766(G26766,G26767,G26756);
  xor GNAME26767(G26767,G32161,G32187);
  and GNAME26768(G26768,G32161,G26756);
  and GNAME26769(G26769,G32187,G26756);
  and GNAME26770(G26770,G32161,G32187);
  or GNAME26771(G26771,G26770,G26769,G26768);
  xor GNAME26781(G26781,G26782,G26741);
  xor GNAME26782(G26782,G27839,G27842);
  and GNAME26783(G26783,G27839,G26741);
  and GNAME26784(G26784,G27842,G26741);
  and GNAME26785(G26785,G27839,G27842);
  or GNAME26786(G26786,G26785,G26784,G26783);
  xor GNAME26796(G26796,G26797,G26786);
  xor GNAME26797(G26797,G27833,G27836);
  and GNAME26798(G26798,G27833,G26786);
  and GNAME26799(G26799,G27836,G26786);
  and GNAME26800(G26800,G27833,G27836);
  or GNAME26801(G26801,G26800,G26799,G26798);
  xor GNAME26811(G26811,G26812,G26771);
  xor GNAME26812(G26812,G32174,G32200);
  and GNAME26813(G26813,G32174,G26771);
  and GNAME26814(G26814,G32200,G26771);
  and GNAME26815(G26815,G32174,G32200);
  or GNAME26816(G26816,G26815,G26814,G26813);
  xor GNAME26826(G26826,G26827,G26816);
  xor GNAME26827(G26827,G32291,G32317);
  and GNAME26828(G26828,G32291,G26816);
  and GNAME26829(G26829,G32317,G26816);
  and GNAME26830(G26830,G32291,G32317);
  or GNAME26831(G26831,G26830,G26829,G26828);
  xor GNAME26841(G26841,G26842,G26801);
  xor GNAME26842(G26842,G27827,G27830);
  and GNAME26843(G26843,G27827,G26801);
  and GNAME26844(G26844,G27830,G26801);
  and GNAME26845(G26845,G27827,G27830);
  or GNAME26846(G26846,G26845,G26844,G26843);
  xor GNAME26856(G26856,G26857,G26846);
  xor GNAME26857(G26857,G27821,G27824);
  and GNAME26858(G26858,G27821,G26846);
  and GNAME26859(G26859,G27824,G26846);
  and GNAME26860(G26860,G27821,G27824);
  or GNAME26861(G26861,G26860,G26859,G26858);
  xor GNAME26871(G26871,G26872,G26831);
  xor GNAME26872(G26872,G32304,G32330);
  and GNAME26873(G26873,G32304,G26831);
  and GNAME26874(G26874,G32330,G26831);
  and GNAME26875(G26875,G32304,G32330);
  or GNAME26876(G26876,G26875,G26874,G26873);
  xor GNAME26886(G26886,G26887,G26876);
  xor GNAME26887(G26887,G32421,G32447);
  and GNAME26888(G26888,G32421,G26876);
  and GNAME26889(G26889,G32447,G26876);
  and GNAME26890(G26890,G32421,G32447);
  or GNAME26891(G26891,G26890,G26889,G26888);
  xor GNAME26901(G26901,G26902,G26861);
  xor GNAME26902(G26902,G27815,G27818);
  and GNAME26903(G26903,G27815,G26861);
  and GNAME26904(G26904,G27818,G26861);
  and GNAME26905(G26905,G27815,G27818);
  or GNAME26906(G26906,G26905,G26904,G26903);
  xor GNAME26916(G26916,G26917,G26906);
  xor GNAME26917(G26917,G27809,G27812);
  and GNAME26918(G26918,G27809,G26906);
  and GNAME26919(G26919,G27812,G26906);
  and GNAME26920(G26920,G27809,G27812);
  or GNAME26921(G26921,G26920,G26919,G26918);
  xor GNAME26931(G26931,G26932,G26921);
  xor GNAME26932(G26932,G27803,G27806);
  and GNAME26933(G26933,G27803,G26921);
  and GNAME26934(G26934,G27806,G26921);
  and GNAME26935(G26935,G27803,G27806);
  or GNAME26936(G26936,G26935,G26934,G26933);
  xor GNAME26946(G26946,G26947,G26891);
  xor GNAME26947(G26947,G32434,G32460);
  and GNAME26948(G26948,G32434,G26891);
  and GNAME26949(G26949,G32460,G26891);
  and GNAME26950(G26950,G32434,G32460);
  or GNAME26951(G26951,G26950,G26949,G26948);
  xor GNAME26961(G26961,G26962,G26951);
  xor GNAME26962(G26962,G32551,G32577);
  and GNAME26963(G26963,G32551,G26951);
  and GNAME26964(G26964,G32577,G26951);
  and GNAME26965(G26965,G32551,G32577);
  or GNAME26966(G26966,G26965,G26964,G26963);
  xor GNAME26976(G26976,G26977,G26936);
  xor GNAME26977(G26977,G27797,G27800);
  and GNAME26978(G26978,G27797,G26936);
  and GNAME26979(G26979,G27800,G26936);
  and GNAME26980(G26980,G27797,G27800);
  or GNAME26981(G26981,G26980,G26979,G26978);
  xor GNAME26991(G26991,G26992,G26981);
  xor GNAME26992(G26992,G27791,G27794);
  and GNAME26993(G26993,G27791,G26981);
  and GNAME26994(G26994,G27794,G26981);
  and GNAME26995(G26995,G27791,G27794);
  or GNAME26996(G26996,G26995,G26994,G26993);
  xor GNAME27006(G27006,G27007,G26966);
  xor GNAME27007(G27007,G32564,G32590);
  and GNAME27008(G27008,G32564,G26966);
  and GNAME27009(G27009,G32590,G26966);
  and GNAME27010(G27010,G32564,G32590);
  or GNAME27011(G27011,G27010,G27009,G27008);
  xor GNAME27021(G27021,G27022,G27011);
  xor GNAME27022(G27022,G32681,G32707);
  and GNAME27023(G27023,G32681,G27011);
  and GNAME27024(G27024,G32707,G27011);
  and GNAME27025(G27025,G32681,G32707);
  or GNAME27026(G27026,G27025,G27024,G27023);
  xor GNAME27036(G27036,G27037,G26996);
  xor GNAME27037(G27037,G27785,G27788);
  and GNAME27038(G27038,G27785,G26996);
  and GNAME27039(G27039,G27788,G26996);
  and GNAME27040(G27040,G27785,G27788);
  or GNAME27041(G27041,G27040,G27039,G27038);
  xor GNAME27051(G27051,G27052,G27041);
  xor GNAME27052(G27052,G27779,G27782);
  and GNAME27053(G27053,G27779,G27041);
  and GNAME27054(G27054,G27782,G27041);
  and GNAME27055(G27055,G27779,G27782);
  or GNAME27056(G27056,G27055,G27054,G27053);
  xor GNAME27066(G27066,G27067,G27026);
  xor GNAME27067(G27067,G32694,G32720);
  and GNAME27068(G27068,G32694,G27026);
  and GNAME27069(G27069,G32720,G27026);
  and GNAME27070(G27070,G32694,G32720);
  or GNAME27071(G27071,G27070,G27069,G27068);
  xor GNAME27081(G27081,G27082,G27071);
  xor GNAME27082(G27082,G32811,G32837);
  and GNAME27083(G27083,G32811,G27071);
  and GNAME27084(G27084,G32837,G27071);
  and GNAME27085(G27085,G32811,G32837);
  or GNAME27086(G27086,G27085,G27084,G27083);
  xor GNAME27096(G27096,G27097,G27056);
  xor GNAME27097(G27097,G27773,G27776);
  and GNAME27098(G27098,G27773,G27056);
  and GNAME27099(G27099,G27776,G27056);
  and GNAME27100(G27100,G27773,G27776);
  or GNAME27101(G27101,G27100,G27099,G27098);
  xor GNAME27111(G27111,G27112,G27101);
  xor GNAME27112(G27112,G27767,G27770);
  and GNAME27113(G27113,G27767,G27101);
  and GNAME27114(G27114,G27770,G27101);
  and GNAME27115(G27115,G27767,G27770);
  or GNAME27116(G27116,G27115,G27114,G27113);
  xor GNAME27126(G27126,G27127,G27086);
  xor GNAME27127(G27127,G32824,G32850);
  and GNAME27128(G27128,G32824,G27086);
  and GNAME27129(G27129,G32850,G27086);
  and GNAME27130(G27130,G32824,G32850);
  or GNAME27131(G27131,G27130,G27129,G27128);
  xor GNAME27141(G27141,G27142,G27131);
  xor GNAME27142(G27142,G33006,G33032);
  and GNAME27143(G27143,G33006,G27131);
  and GNAME27144(G27144,G33032,G27131);
  and GNAME27145(G27145,G33006,G33032);
  or GNAME27146(G27146,G27145,G27144,G27143);
  xor GNAME27156(G27156,G27157,G27116);
  xor GNAME27157(G27157,G27761,G27764);
  and GNAME27158(G27158,G27761,G27116);
  and GNAME27159(G27159,G27764,G27116);
  and GNAME27160(G27160,G27761,G27764);
  or GNAME27161(G27161,G27160,G27159,G27158);
  xor GNAME27171(G27171,G27172,G27161);
  xor GNAME27172(G27172,G27755,G27758);
  and GNAME27173(G27173,G27755,G27161);
  and GNAME27174(G27174,G27758,G27161);
  and GNAME27175(G27175,G27755,G27758);
  or GNAME27176(G27176,G27175,G27174,G27173);
  xor GNAME27186(G27186,G27187,G27146);
  xor GNAME27187(G27187,G33019,G33045);
  and GNAME27188(G27188,G33019,G27146);
  and GNAME27189(G27189,G33045,G27146);
  and GNAME27190(G27190,G33019,G33045);
  or GNAME27191(G27191,G27190,G27189,G27188);
  xor GNAME27201(G27201,G27202,G27191);
  xor GNAME27202(G27202,G33201,G33227);
  and GNAME27203(G27203,G33201,G27191);
  and GNAME27204(G27204,G33227,G27191);
  and GNAME27205(G27205,G33201,G33227);
  or GNAME27206(G27206,G27205,G27204,G27203);
  xor GNAME27216(G27216,G27217,G27206);
  xor GNAME27217(G27217,G33214,G33240);
  and GNAME27218(G27218,G33214,G27206);
  and GNAME27219(G27219,G33240,G27206);
  and GNAME27220(G27220,G33214,G33240);
  or GNAME27221(G27221,G27220,G27219,G27218);
  xor GNAME27231(G27231,G27232,G27176);
  xor GNAME27232(G27232,G27749,G27752);
  and GNAME27233(G27233,G27749,G27176);
  and GNAME27234(G27234,G27752,G27176);
  and GNAME27235(G27235,G27749,G27752);
  or GNAME27236(G27236,G27235,G27234,G27233);
  xor GNAME27246(G27246,G27247,G27236);
  xor GNAME27247(G27247,G27743,G27746);
  and GNAME27248(G27248,G27743,G27236);
  and GNAME27249(G27249,G27746,G27236);
  and GNAME27250(G27250,G27743,G27746);
  or GNAME27251(G27251,G27250,G27249,G27248);
  xor GNAME27261(G27261,G27262,G27221);
  xor GNAME27262(G27262,G33396,G33422);
  and GNAME27263(G27263,G33396,G27221);
  and GNAME27264(G27264,G33422,G27221);
  and GNAME27265(G27265,G33396,G33422);
  or GNAME27266(G27266,G27265,G27264,G27263);
  xor GNAME27276(G27276,G27277,G27266);
  xor GNAME27277(G27277,G33409,G33435);
  and GNAME27278(G27278,G33409,G27266);
  and GNAME27279(G27279,G33435,G27266);
  and GNAME27280(G27280,G33409,G33435);
  or GNAME27281(G27281,G27280,G27279,G27278);
  xor GNAME27291(G27291,G27292,G27251);
  xor GNAME27292(G27292,G27737,G27740);
  and GNAME27293(G27293,G27737,G27251);
  and GNAME27294(G27294,G27740,G27251);
  and GNAME27295(G27295,G27737,G27740);
  or GNAME27296(G27296,G27295,G27294,G27293);
  xor GNAME27306(G27306,G27307,G27296);
  xor GNAME27307(G27307,G27731,G27734);
  and GNAME27308(G27308,G27731,G27296);
  and GNAME27309(G27309,G27734,G27296);
  and GNAME27310(G27310,G27731,G27734);
  or GNAME27311(G27311,G27310,G27309,G27308);
  xor GNAME27321(G27321,G27322,G27281);
  xor GNAME27322(G27322,G33578,G33604);
  and GNAME27323(G27323,G33578,G27281);
  and GNAME27324(G27324,G33604,G27281);
  and GNAME27325(G27325,G33578,G33604);
  or GNAME27326(G27326,G27325,G27324,G27323);
  xor GNAME27336(G27336,G27337,G27326);
  xor GNAME27337(G27337,G33591,G33617);
  and GNAME27338(G27338,G33591,G27326);
  and GNAME27339(G27339,G33617,G27326);
  and GNAME27340(G27340,G33591,G33617);
  or GNAME27341(G27341,G27340,G27339,G27338);
  xor GNAME27351(G27351,G27352,G27311);
  xor GNAME27352(G27352,G27725,G27728);
  and GNAME27353(G27353,G27725,G27311);
  and GNAME27354(G27354,G27728,G27311);
  and GNAME27355(G27355,G27725,G27728);
  or GNAME27356(G27356,G27355,G27354,G27353);
  xor GNAME27366(G27366,G27367,G27356);
  xor GNAME27367(G27367,G27719,G27722);
  and GNAME27368(G27368,G27719,G27356);
  and GNAME27369(G27369,G27722,G27356);
  and GNAME27370(G27370,G27719,G27722);
  or GNAME27371(G27371,G27370,G27369,G27368);
  xor GNAME27381(G27381,G27382,G27341);
  xor GNAME27382(G27382,G33773,G33799);
  and GNAME27383(G27383,G33773,G27341);
  and GNAME27384(G27384,G33799,G27341);
  and GNAME27385(G27385,G33773,G33799);
  or GNAME27386(G27386,G27385,G27384,G27383);
  xor GNAME27396(G27396,G27397,G27386);
  xor GNAME27397(G27397,G33786,G33812);
  and GNAME27398(G27398,G33786,G27386);
  and GNAME27399(G27399,G33812,G27386);
  and GNAME27400(G27400,G33786,G33812);
  or GNAME27401(G27401,G27400,G27399,G27398);
  xor GNAME27411(G27411,G27412,G27371);
  xor GNAME27412(G27412,G27713,G27716);
  and GNAME27413(G27413,G27713,G27371);
  and GNAME27414(G27414,G27716,G27371);
  and GNAME27415(G27415,G27713,G27716);
  or GNAME27416(G27416,G27415,G27414,G27413);
  xor GNAME27426(G27426,G27427,G27416);
  xor GNAME27427(G27427,G27707,G27710);
  and GNAME27428(G27428,G27707,G27416);
  and GNAME27429(G27429,G27710,G27416);
  and GNAME27430(G27430,G27707,G27710);
  or GNAME27431(G27431,G27430,G27429,G27428);
  xor GNAME27441(G27441,G27442,G27401);
  xor GNAME27442(G27442,G33955,G33981);
  and GNAME27443(G27443,G33955,G27401);
  and GNAME27444(G27444,G33981,G27401);
  and GNAME27445(G27445,G33955,G33981);
  or GNAME27446(G27446,G27445,G27444,G27443);
  xor GNAME27456(G27456,G27457,G27446);
  xor GNAME27457(G27457,G33968,G33994);
  and GNAME27458(G27458,G33968,G27446);
  and GNAME27459(G27459,G33994,G27446);
  and GNAME27460(G27460,G33968,G33994);
  or GNAME27461(G27461,G27460,G27459,G27458);
  xor GNAME27471(G27471,G27472,G27431);
  xor GNAME27472(G27472,G27701,G27704);
  and GNAME27473(G27473,G27701,G27431);
  and GNAME27474(G27474,G27704,G27431);
  and GNAME27475(G27475,G27701,G27704);
  or GNAME27476(G27476,G27475,G27474,G27473);
  xor GNAME27486(G27486,G27487,G27476);
  xor GNAME27487(G27487,G27695,G27698);
  and GNAME27488(G27488,G27695,G27476);
  and GNAME27489(G27489,G27698,G27476);
  and GNAME27490(G27490,G27695,G27698);
  or GNAME27491(G27491,G27490,G27489,G27488);
  xor GNAME27501(G27501,G27502,G27461);
  xor GNAME27502(G27502,G34423,G34449);
  and GNAME27503(G27503,G34423,G27461);
  and GNAME27504(G27504,G34449,G27461);
  and GNAME27505(G27505,G34423,G34449);
  or GNAME27506(G27506,G27505,G27504,G27503);
  xor GNAME27516(G27516,G27517,G27491);
  xor GNAME27517(G27517,G27689,G27692);
  and GNAME27518(G27518,G27689,G27491);
  and GNAME27519(G27519,G27692,G27491);
  and GNAME27520(G27520,G27689,G27692);
  or GNAME27521(G27521,G27520,G27519,G27518);
  xor GNAME27531(G27531,G27532,G27521);
  xor GNAME27532(G27532,G27683,G27686);
  and GNAME27533(G27533,G27683,G27521);
  and GNAME27534(G27534,G27686,G27521);
  and GNAME27535(G27535,G27683,G27686);
  or GNAME27536(G27536,G27535,G27534,G27533);
  xor GNAME27546(G27546,G27547,G27536);
  xor GNAME27547(G27547,G27677,G27680);
  and GNAME27548(G27548,G27677,G27536);
  and GNAME27549(G27549,G27680,G27536);
  and GNAME27550(G27550,G27677,G27680);
  or GNAME27551(G27551,G27550,G27549,G27548);
  xor GNAME27561(G27561,G27562,G27551);
  xor GNAME27562(G27562,G27671,G27674);
  and GNAME27563(G27563,G27671,G27551);
  and GNAME27564(G27564,G27674,G27551);
  and GNAME27565(G27565,G27671,G27674);
  or GNAME27566(G27566,G27565,G27564,G27563);
  and GNAME27567(G27567,G27860,G27857);
  and GNAME27568(G27568,G31680,G31706);
  and GNAME27569(G27569,G2760,G31693);
  and GNAME27570(G27570,G29944,G29953);
  and GNAME27571(G27571,G29947,G29956);
  and GNAME27572(G27572,G29950,G29959);
  and GNAME27573(G27573,G28618,G34596);
  and GNAME27574(G27574,G32941,G31442);
  or GNAME27575(G27575,G27574,G27573);
  and GNAME27576(G27576,G28612,G34596);
  and GNAME27577(G27577,G32928,G31442);
  or GNAME27578(G27578,G27577,G27576);
  and GNAME27579(G27579,G28606,G34596);
  and GNAME27580(G27580,G32915,G31442);
  or GNAME27581(G27581,G27580,G27579);
  and GNAME27582(G27582,G28594,G34596);
  and GNAME27583(G27583,G32902,G31442);
  or GNAME27584(G27584,G27583,G27582);
  and GNAME27585(G27585,G31436,G34596);
  and GNAME27586(G27586,G32863,G31442);
  or GNAME27587(G27587,G27586,G27585);
  and GNAME27588(G27588,G28636,G34596);
  and GNAME27589(G27589,G33110,G31442);
  or GNAME27590(G27590,G27589,G27588);
  and GNAME27591(G27591,G28630,G34596);
  and GNAME27592(G27592,G33097,G31442);
  or GNAME27593(G27593,G27592,G27591);
  and GNAME27594(G27594,G28624,G34596);
  and GNAME27595(G27595,G33084,G31442);
  or GNAME27596(G27596,G27595,G27594);
  and GNAME27597(G27597,G28642,G34597);
  and GNAME27598(G27598,G33123,G31442);
  or GNAME27599(G27599,G27598,G27597);
  and GNAME27600(G27600,G34597,G28648);
  and GNAME27601(G27601,G33279,G31442);
  or GNAME27602(G27602,G27601,G27600);
  and GNAME27603(G27603,G28672,G34596);
  and GNAME27604(G27604,G33331,G31442);
  or GNAME27605(G27605,G27604,G27603);
  and GNAME27606(G27606,G28666,G34596);
  and GNAME27607(G27607,G33318,G31442);
  or GNAME27608(G27608,G27607,G27606);
  and GNAME27609(G27609,G28660,G34596);
  and GNAME27610(G27610,G33305,G31442);
  or GNAME27611(G27611,G27610,G27609);
  and GNAME27612(G27612,G28654,G34596);
  and GNAME27613(G27613,G33292,G31442);
  or GNAME27614(G27614,G27613,G27612);
  and GNAME27615(G27615,G28702,G34596);
  and GNAME27616(G27616,G33656,G31442);
  or GNAME27617(G27617,G27616,G27615);
  and GNAME27618(G27618,G28696,G34596);
  and GNAME27619(G27619,G33513,G31442);
  or GNAME27620(G27620,G27619,G27618);
  and GNAME27621(G27621,G28690,G34596);
  and GNAME27622(G27622,G33500,G31442);
  or GNAME27623(G27623,G27622,G27621);
  and GNAME27624(G27624,G28684,G34596);
  and GNAME27625(G27625,G33487,G31442);
  or GNAME27626(G27626,G27625,G27624);
  and GNAME27627(G27627,G28678,G34596);
  and GNAME27628(G27628,G33474,G31442);
  or GNAME27629(G27629,G27628,G27627);
  and GNAME27630(G27630,G28726,G34596);
  and GNAME27631(G27631,G33708,G31442);
  or GNAME27632(G27632,G27631,G27630);
  and GNAME27633(G27633,G28720,G34596);
  and GNAME27634(G27634,G33695,G31442);
  or GNAME27635(G27635,G27634,G27633);
  and GNAME27636(G27636,G28714,G34596);
  and GNAME27637(G27637,G33682,G31442);
  or GNAME27638(G27638,G27637,G27636);
  and GNAME27639(G27639,G28708,G34596);
  and GNAME27640(G27640,G33669,G31442);
  or GNAME27641(G27641,G27640,G27639);
  and GNAME27642(G27642,G28756,G34596);
  and GNAME27643(G27643,G34371,G31442);
  or GNAME27644(G27644,G27643,G27642);
  and GNAME27645(G27645,G28750,G34596);
  and GNAME27646(G27646,G33890,G31442);
  or GNAME27647(G27647,G27646,G27645);
  and GNAME27648(G27648,G28744,G34596);
  and GNAME27649(G27649,G33877,G31442);
  or GNAME27650(G27650,G27649,G27648);
  and GNAME27651(G27651,G28738,G34596);
  and GNAME27652(G27652,G33864,G31442);
  or GNAME27653(G27653,G27652,G27651);
  and GNAME27654(G27654,G28732,G34596);
  and GNAME27655(G27655,G33851,G31442);
  or GNAME27656(G27656,G27655,G27654);
  and GNAME27657(G27657,G31584,G34596);
  and GNAME27658(G27658,G34345,G31442);
  or GNAME27659(G27659,G27658,G27657);
  and GNAME27660(G27660,G28600,G34596);
  and GNAME27661(G27661,G34410,G31442);
  or GNAME27662(G27662,G27661,G27660);
  and GNAME27663(G27663,G28768,G34596);
  and GNAME27664(G27664,G34397,G31442);
  or GNAME27665(G27665,G27664,G27663);
  and GNAME27666(G27666,G28762,G34596);
  and GNAME27667(G27667,G34384,G31442);
  or GNAME27668(G27668,G27667,G27666);
  and GNAME27669(G27669,G31585,G34653);
  and GNAME27670(G27670,G34332,G31519);
  or GNAME27671(G27671,G27670,G27669);
  and GNAME27672(G27672,G31586,G34652);
  and GNAME27673(G27673,G34358,G31518);
  or GNAME27674(G27674,G27673,G27672);
  and GNAME27675(G27675,G28582,G34653);
  and GNAME27676(G27676,G33838,G31519);
  or GNAME27677(G27677,G27676,G27675);
  and GNAME27678(G27678,G28588,G34652);
  and GNAME27679(G27679,G33916,G31518);
  or GNAME27680(G27680,G27679,G27678);
  and GNAME27681(G27681,G28570,G34653);
  and GNAME27682(G27682,G33825,G31519);
  or GNAME27683(G27683,G27682,G27681);
  and GNAME27684(G27684,G28576,G34652);
  and GNAME27685(G27685,G33903,G31518);
  or GNAME27686(G27686,G27685,G27684);
  and GNAME27687(G27687,G28558,G34653);
  and GNAME27688(G27688,G33643,G31519);
  or GNAME27689(G27689,G27688,G27687);
  and GNAME27690(G27690,G28564,G34652);
  and GNAME27691(G27691,G33734,G31518);
  or GNAME27692(G27692,G27691,G27690);
  and GNAME27693(G27693,G28546,G34653);
  and GNAME27694(G27694,G33630,G31519);
  or GNAME27695(G27695,G27694,G27693);
  and GNAME27696(G27696,G28552,G34652);
  and GNAME27697(G27697,G33721,G31518);
  or GNAME27698(G27698,G27697,G27696);
  and GNAME27699(G27699,G28534,G34653);
  and GNAME27700(G27700,G33461,G31519);
  or GNAME27701(G27701,G27700,G27699);
  and GNAME27702(G27702,G28540,G34652);
  and GNAME27703(G27703,G33539,G31518);
  or GNAME27704(G27704,G27703,G27702);
  and GNAME27705(G27705,G28522,G34653);
  and GNAME27706(G27706,G33448,G31519);
  or GNAME27707(G27707,G27706,G27705);
  and GNAME27708(G27708,G28528,G34652);
  and GNAME27709(G27709,G33526,G31518);
  or GNAME27710(G27710,G27709,G27708);
  and GNAME27711(G27711,G28510,G34653);
  and GNAME27712(G27712,G33266,G31519);
  or GNAME27713(G27713,G27712,G27711);
  and GNAME27714(G27714,G28516,G34652);
  and GNAME27715(G27715,G33357,G31518);
  or GNAME27716(G27716,G27715,G27714);
  and GNAME27717(G27717,G28498,G34653);
  and GNAME27718(G27718,G33253,G31519);
  or GNAME27719(G27719,G27718,G27717);
  and GNAME27720(G27720,G28504,G34652);
  and GNAME27721(G27721,G33344,G31518);
  or GNAME27722(G27722,G27721,G27720);
  and GNAME27723(G27723,G28486,G34653);
  and GNAME27724(G27724,G33071,G31519);
  or GNAME27725(G27725,G27724,G27723);
  and GNAME27726(G27726,G28492,G34652);
  and GNAME27727(G27727,G33149,G31518);
  or GNAME27728(G27728,G27727,G27726);
  and GNAME27729(G27729,G28474,G34653);
  and GNAME27730(G27730,G33058,G31519);
  or GNAME27731(G27731,G27730,G27729);
  and GNAME27732(G27732,G28480,G34652);
  and GNAME27733(G27733,G33136,G31518);
  or GNAME27734(G27734,G27733,G27732);
  and GNAME27735(G27735,G28462,G34653);
  and GNAME27736(G27736,G32889,G31519);
  or GNAME27737(G27737,G27736,G27735);
  and GNAME27738(G27738,G28468,G34652);
  and GNAME27739(G27739,G32967,G31518);
  or GNAME27740(G27740,G27739,G27738);
  and GNAME27741(G27741,G28450,G34653);
  and GNAME27742(G27742,G32876,G31519);
  or GNAME27743(G27743,G27742,G27741);
  and GNAME27744(G27744,G28456,G34652);
  and GNAME27745(G27745,G32954,G31518);
  or GNAME27746(G27746,G27745,G27744);
  and GNAME27747(G27747,G28438,G34653);
  and GNAME27748(G27748,G32746,G31519);
  or GNAME27749(G27749,G27748,G27747);
  and GNAME27750(G27750,G28444,G34652);
  and GNAME27751(G27751,G32772,G31518);
  or GNAME27752(G27752,G27751,G27750);
  and GNAME27753(G27753,G28426,G34653);
  and GNAME27754(G27754,G32733,G31519);
  or GNAME27755(G27755,G27754,G27753);
  and GNAME27756(G27756,G28432,G34652);
  and GNAME27757(G27757,G32759,G31518);
  or GNAME27758(G27758,G27757,G27756);
  and GNAME27759(G27759,G28414,G34653);
  and GNAME27760(G27760,G32616,G31519);
  or GNAME27761(G27761,G27760,G27759);
  and GNAME27762(G27762,G28420,G34652);
  and GNAME27763(G27763,G32642,G31518);
  or GNAME27764(G27764,G27763,G27762);
  and GNAME27765(G27765,G28402,G34653);
  and GNAME27766(G27766,G32603,G31519);
  or GNAME27767(G27767,G27766,G27765);
  and GNAME27768(G27768,G28408,G34652);
  and GNAME27769(G27769,G32629,G31518);
  or GNAME27770(G27770,G27769,G27768);
  and GNAME27771(G27771,G28390,G34653);
  and GNAME27772(G27772,G32486,G31519);
  or GNAME27773(G27773,G27772,G27771);
  and GNAME27774(G27774,G28396,G34652);
  and GNAME27775(G27775,G32512,G31518);
  or GNAME27776(G27776,G27775,G27774);
  and GNAME27777(G27777,G28378,G34653);
  and GNAME27778(G27778,G32473,G31519);
  or GNAME27779(G27779,G27778,G27777);
  and GNAME27780(G27780,G28384,G34652);
  and GNAME27781(G27781,G32499,G31518);
  or GNAME27782(G27782,G27781,G27780);
  and GNAME27783(G27783,G28366,G34653);
  and GNAME27784(G27784,G32356,G31519);
  or GNAME27785(G27785,G27784,G27783);
  and GNAME27786(G27786,G28372,G34652);
  and GNAME27787(G27787,G32382,G31518);
  or GNAME27788(G27788,G27787,G27786);
  and GNAME27789(G27789,G28342,G34653);
  and GNAME27790(G27790,G32343,G31519);
  or GNAME27791(G27791,G27790,G27789);
  and GNAME27792(G27792,G28348,G34652);
  and GNAME27793(G27793,G32369,G31518);
  or GNAME27794(G27794,G27793,G27792);
  and GNAME27795(G27795,G28330,G34653);
  and GNAME27796(G27796,G32226,G31519);
  or GNAME27797(G27797,G27796,G27795);
  and GNAME27798(G27798,G28336,G34652);
  and GNAME27799(G27799,G32252,G31518);
  or GNAME27800(G27800,G27799,G27798);
  and GNAME27801(G27801,G34661,G28354);
  and GNAME27802(G27802,G32213,G31519);
  or GNAME27803(G27803,G27802,G27801);
  and GNAME27804(G27804,G34660,G28360);
  and GNAME27805(G27805,G32239,G31518);
  or GNAME27806(G27806,G27805,G27804);
  and GNAME27807(G27807,G28318,G34661);
  and GNAME27808(G27808,G32096,G31519);
  or GNAME27809(G27809,G27808,G27807);
  and GNAME27810(G27810,G28324,G34660);
  and GNAME27811(G27811,G32122,G31518);
  or GNAME27812(G27812,G27811,G27810);
  and GNAME27813(G27813,G28306,G34653);
  and GNAME27814(G27814,G32083,G31519);
  or GNAME27815(G27815,G27814,G27813);
  and GNAME27816(G27816,G28312,G34652);
  and GNAME27817(G27817,G32109,G31518);
  or GNAME27818(G27818,G27817,G27816);
  and GNAME27819(G27819,G28294,G34653);
  and GNAME27820(G27820,G31966,G31519);
  or GNAME27821(G27821,G27820,G27819);
  and GNAME27822(G27822,G28300,G34652);
  and GNAME27823(G27823,G31992,G31518);
  or GNAME27824(G27824,G27823,G27822);
  and GNAME27825(G27825,G28282,G34653);
  and GNAME27826(G27826,G31953,G31519);
  or GNAME27827(G27827,G27826,G27825);
  and GNAME27828(G27828,G28288,G34652);
  and GNAME27829(G27829,G31979,G31518);
  or GNAME27830(G27830,G27829,G27828);
  and GNAME27831(G27831,G28270,G34653);
  and GNAME27832(G27832,G31836,G31519);
  or GNAME27833(G27833,G27832,G27831);
  and GNAME27834(G27834,G28276,G34652);
  and GNAME27835(G27835,G31862,G31518);
  or GNAME27836(G27836,G27835,G27834);
  and GNAME27837(G27837,G28258,G34653);
  and GNAME27838(G27838,G31823,G31519);
  or GNAME27839(G27839,G27838,G27837);
  and GNAME27840(G27840,G28264,G34652);
  and GNAME27841(G27841,G31849,G31518);
  or GNAME27842(G27842,G27841,G27840);
  and GNAME27843(G27843,G28246,G34653);
  and GNAME27844(G27844,G31732,G31519);
  or GNAME27845(G27845,G27844,G27843);
  and GNAME27846(G27846,G28252,G34652);
  and GNAME27847(G27847,G31758,G31518);
  or GNAME27848(G27848,G27847,G27846);
  and GNAME27849(G27849,G28234,G34653);
  and GNAME27850(G27850,G31719,G31519);
  or GNAME27851(G27851,G27850,G27849);
  and GNAME27852(G27852,G28240,G34652);
  and GNAME27853(G27853,G31745,G31518);
  or GNAME27854(G27854,G27853,G27852);
  and GNAME27855(G27855,G31437,G34653);
  and GNAME27856(G27856,G31628,G31519);
  or GNAME27857(G27857,G27856,G27855);
  and GNAME27858(G27858,G31438,G34652);
  and GNAME27859(G27859,G31641,G31518);
  or GNAME27860(G27860,G27859,G27858);
  not GNAME27861(G27861,G27863);
  not GNAME27862(G27862,G34677);
  and GNAME27863(G27863,G34654,G27862);
  not GNAME27864(G27864,G27866);
  not GNAME27865(G27865,G34678);
  and GNAME27866(G27866,G34655,G27865);
  not GNAME27867(G27867,G27869);
  not GNAME27868(G27868,G34679);
  and GNAME27869(G27869,G34656,G27868);
  not GNAME27870(G27870,G27872);
  not GNAME27871(G27871,G34677);
  and GNAME27872(G27872,G34657,G27871);
  not GNAME27873(G27873,G27875);
  not GNAME27874(G27874,G34678);
  and GNAME27875(G27875,G34658,G27874);
  not GNAME27876(G27876,G27878);
  not GNAME27877(G27877,G34679);
  and GNAME27878(G27878,G34659,G27877);
  not GNAME27879(G27879,G27881);
  not GNAME27880(G27880,G34677);
  and GNAME27881(G27881,G34674,G27880);
  not GNAME27882(G27882,G27884);
  not GNAME27883(G27883,G34678);
  and GNAME27884(G27884,G34675,G27883);
  not GNAME27885(G27885,G27887);
  not GNAME27886(G27886,G34679);
  and GNAME27887(G27887,G34676,G27886);
  not GNAME27888(G27888,G27890);
  not GNAME27889(G27889,G34710);
  and GNAME27890(G27890,G34689,G27889);
  not GNAME27891(G27891,G27893);
  not GNAME27892(G27892,G34711);
  and GNAME27893(G27893,G34690,G27892);
  not GNAME27894(G27894,G27896);
  not GNAME27895(G27895,G34712);
  and GNAME27896(G27896,G34691,G27895);
  not GNAME27897(G27897,G27899);
  not GNAME27898(G27898,G34710);
  and GNAME27899(G27899,G34704,G27898);
  not GNAME27900(G27900,G27902);
  not GNAME27901(G27901,G34711);
  and GNAME27902(G27902,G34705,G27901);
  not GNAME27903(G27903,G27905);
  not GNAME27904(G27904,G34712);
  and GNAME27905(G27905,G34706,G27904);
  not GNAME27906(G27906,G27908);
  not GNAME27907(G27907,G34710);
  and GNAME27908(G27908,G34719,G27907);
  not GNAME27909(G27909,G27911);
  not GNAME27910(G27910,G34711);
  and GNAME27911(G27911,G34720,G27910);
  not GNAME27912(G27912,G27914);
  not GNAME27913(G27913,G34712);
  and GNAME27914(G27914,G34721,G27913);
  not GNAME27915(G27915,G27917);
  not GNAME27916(G27916,G34710);
  and GNAME27917(G27917,G34707,G27916);
  not GNAME27918(G27918,G27920);
  not GNAME27919(G27919,G34711);
  and GNAME27920(G27920,G34708,G27919);
  not GNAME27921(G27921,G27923);
  not GNAME27922(G27922,G34712);
  and GNAME27923(G27923,G34709,G27922);
  not GNAME27924(G27924,G27926);
  not GNAME27925(G27925,G34710);
  and GNAME27926(G27926,G34722,G27925);
  not GNAME27927(G27927,G27929);
  not GNAME27928(G27928,G34711);
  and GNAME27929(G27929,G34723,G27928);
  not GNAME27930(G27930,G27932);
  not GNAME27931(G27931,G34712);
  and GNAME27932(G27932,G34724,G27931);
  xor GNAME27933(G27933,G27934,G28921);
  xor GNAME27934(G27934,G29589,G28987);
  xor GNAME27935(G27935,G27936,G28922);
  xor GNAME27936(G27936,G29591,G28988);
  xor GNAME27937(G27937,G27938,G28923);
  xor GNAME27938(G27938,G29593,G28989);
  xor GNAME27939(G27939,G27940,G26186);
  xor GNAME27940(G27940,G34475,G3552);
  not GNAME27941(G27941,G27943);
  not GNAME27942(G27942,G34677);
  or GNAME27943(G27943,G34785,G27942);
  not GNAME27944(G27944,G27946);
  not GNAME27945(G27945,G34678);
  or GNAME27946(G27946,G34786,G27945);
  not GNAME27947(G27947,G27949);
  not GNAME27948(G27948,G34679);
  or GNAME27949(G27949,G34787,G27948);
  not GNAME27950(G27950,G27952);
  not GNAME27951(G27951,G34677);
  or GNAME27952(G27952,G34731,G27951);
  not GNAME27953(G27953,G27955);
  not GNAME27954(G27954,G34678);
  or GNAME27955(G27955,G34732,G27954);
  not GNAME27956(G27956,G27958);
  not GNAME27957(G27957,G34679);
  or GNAME27958(G27958,G34733,G27957);
  not GNAME27959(G27959,G27961);
  not GNAME27960(G27960,G26451);
  or GNAME27961(G27961,G34725,G27960);
  not GNAME27962(G27962,G27964);
  not GNAME27963(G27963,G26436);
  or GNAME27964(G27964,G34725,G27963);
  not GNAME27965(G27965,G27967);
  not GNAME27966(G27966,G26421);
  or GNAME27967(G27967,G34725,G27966);
  not GNAME27968(G27968,G27970);
  not GNAME27969(G27969,G26406);
  or GNAME27970(G27970,G34725,G27969);
  not GNAME27971(G27971,G27973);
  not GNAME27972(G27972,G26391);
  or GNAME27973(G27973,G34725,G27972);
  not GNAME27974(G27974,G27976);
  not GNAME27975(G27975,G26376);
  or GNAME27976(G27976,G34725,G27975);
  not GNAME27977(G27977,G27979);
  not GNAME27978(G27978,G26361);
  or GNAME27979(G27979,G34729,G27978);
  not GNAME27980(G27980,G27982);
  not GNAME27981(G27981,G26346);
  or GNAME27982(G27982,G34729,G27981);
  not GNAME27983(G27983,G27985);
  not GNAME27984(G27984,G26571);
  or GNAME27985(G27985,G34730,G27984);
  not GNAME27986(G27986,G27988);
  not GNAME27987(G27987,G26556);
  or GNAME27988(G27988,G34730,G27987);
  not GNAME27989(G27989,G27991);
  not GNAME27990(G27990,G26541);
  or GNAME27991(G27991,G34730,G27990);
  not GNAME27992(G27992,G27994);
  not GNAME27993(G27993,G26526);
  or GNAME27994(G27994,G34730,G27993);
  not GNAME27995(G27995,G27997);
  not GNAME27996(G27996,G26511);
  or GNAME27997(G27997,G34730,G27996);
  not GNAME27998(G27998,G28000);
  not GNAME27999(G27999,G26496);
  or GNAME28000(G28000,G34730,G27999);
  not GNAME28001(G28001,G28003);
  not GNAME28002(G28002,G26481);
  or GNAME28003(G28003,G34730,G28002);
  not GNAME28004(G28004,G28006);
  not GNAME28005(G28005,G26466);
  or GNAME28006(G28006,G34730,G28005);
  not GNAME28007(G28007,G28009);
  not GNAME28008(G28008,G26331);
  or GNAME28009(G28009,G34729,G28008);
  not GNAME28010(G28010,G28012);
  not GNAME28011(G28011,G26316);
  or GNAME28012(G28012,G34729,G28011);
  not GNAME28013(G28013,G28015);
  not GNAME28014(G28014,G26301);
  or GNAME28015(G28015,G34729,G28014);
  not GNAME28016(G28016,G28018);
  not GNAME28017(G28017,G26286);
  or GNAME28018(G28018,G34729,G28017);
  not GNAME28019(G28019,G28021);
  not GNAME28020(G28020,G26271);
  or GNAME28021(G28021,G34729,G28020);
  not GNAME28022(G28022,G28024);
  not GNAME28023(G28023,G26256);
  or GNAME28024(G28024,G34729,G28023);
  not GNAME28025(G28025,G28027);
  not GNAME28026(G28026,G26211);
  or GNAME28027(G28027,G34730,G28026);
  not GNAME28028(G28028,G28030);
  not GNAME28029(G28029,G26676);
  or GNAME28030(G28030,G34729,G28029);
  not GNAME28031(G28031,G28033);
  not GNAME28032(G28032,G26661);
  or GNAME28033(G28033,G34729,G28032);
  not GNAME28034(G28034,G28036);
  not GNAME28035(G28035,G26646);
  or GNAME28036(G28036,G34729,G28035);
  not GNAME28037(G28037,G28039);
  not GNAME28038(G28038,G26631);
  or GNAME28039(G28039,G34729,G28038);
  not GNAME28040(G28040,G28042);
  not GNAME28041(G28041,G26616);
  or GNAME28042(G28042,G34730,G28041);
  not GNAME28043(G28043,G28045);
  not GNAME28044(G28044,G26601);
  or GNAME28045(G28045,G34730,G28044);
  not GNAME28046(G28046,G28048);
  not GNAME28047(G28047,G26586);
  or GNAME28048(G28048,G34730,G28047);
  not GNAME28049(G28049,G28051);
  not GNAME28050(G28050,G34677);
  or GNAME28051(G28051,G34737,G28050);
  not GNAME28052(G28052,G28054);
  not GNAME28053(G28053,G34678);
  or GNAME28054(G28054,G34738,G28053);
  not GNAME28055(G28055,G28057);
  not GNAME28056(G28056,G34679);
  or GNAME28057(G28057,G34739,G28056);
  not GNAME28058(G28058,G28060);
  not GNAME28059(G28059,G34677);
  or GNAME28060(G28060,G34746,G28059);
  not GNAME28061(G28061,G28063);
  not GNAME28062(G28062,G34678);
  or GNAME28063(G28063,G34747,G28062);
  not GNAME28064(G28064,G28066);
  not GNAME28065(G28065,G34679);
  or GNAME28066(G28066,G34748,G28065);
  not GNAME28067(G28067,G28069);
  not GNAME28068(G28068,G34677);
  or GNAME28069(G28069,G34809,G28068);
  not GNAME28070(G28070,G28072);
  not GNAME28071(G28071,G34678);
  or GNAME28072(G28072,G34810,G28071);
  not GNAME28073(G28073,G28075);
  not GNAME28074(G28074,G34679);
  or GNAME28075(G28075,G34811,G28074);
  not GNAME28076(G28076,G28078);
  not GNAME28077(G28077,G34710);
  or GNAME28078(G28078,G34812,G28077);
  not GNAME28079(G28079,G28081);
  not GNAME28080(G28080,G34711);
  or GNAME28081(G28081,G34813,G28080);
  not GNAME28082(G28082,G28084);
  not GNAME28083(G28083,G34712);
  or GNAME28084(G28084,G34814,G28083);
  not GNAME28085(G28085,G28087);
  not GNAME28086(G28086,G34710);
  or GNAME28087(G28087,G34773,G28086);
  not GNAME28088(G28088,G28090);
  not GNAME28089(G28089,G34711);
  or GNAME28090(G28090,G34775,G28089);
  not GNAME28091(G28091,G28093);
  not GNAME28092(G28092,G34712);
  or GNAME28093(G28093,G34777,G28092);
  not GNAME28094(G28094,G28096);
  not GNAME28095(G28095,G34710);
  or GNAME28096(G28096,G34774,G28095);
  not GNAME28097(G28097,G28099);
  not GNAME28098(G28098,G34711);
  or GNAME28099(G28099,G34776,G28098);
  not GNAME28100(G28100,G28102);
  not GNAME28101(G28101,G34712);
  or GNAME28102(G28102,G34778,G28101);
  or GNAME28103(G28103,G26181,G27939);
  xor GNAME28108(G28108,G29737,G29740);
  and GNAME28109(G28109,G29737,G29740);
  xor GNAME28114(G28114,G29743,G29746);
  and GNAME28115(G28115,G29743,G29746);
  xor GNAME28120(G28120,G29749,G29752);
  and GNAME28121(G28121,G29749,G29752);
  xor GNAME28126(G28126,G29755,G29758);
  and GNAME28127(G28127,G29755,G29758);
  xor GNAME28132(G28132,G29761,G29764);
  and GNAME28133(G28133,G29761,G29764);
  xor GNAME28138(G28138,G29767,G29770);
  and GNAME28139(G28139,G29767,G29770);
  xor GNAME28144(G28144,G29791,G29794);
  and GNAME28145(G28145,G29791,G29794);
  xor GNAME28150(G28150,G29797,G29800);
  and GNAME28151(G28151,G29797,G29800);
  xor GNAME28156(G28156,G29803,G29806);
  and GNAME28157(G28157,G29803,G29806);
  xor GNAME28162(G28162,G29827,G29830);
  and GNAME28163(G28163,G29827,G29830);
  xor GNAME28168(G28168,G29833,G29836);
  and GNAME28169(G28169,G29833,G29836);
  xor GNAME28174(G28174,G29839,G29842);
  and GNAME28175(G28175,G29839,G29842);
  xor GNAME28180(G28180,G29863,G29866);
  and GNAME28181(G28181,G29863,G29866);
  xor GNAME28186(G28186,G29869,G29872);
  and GNAME28187(G28187,G29869,G29872);
  xor GNAME28192(G28192,G29875,G29878);
  and GNAME28193(G28193,G29875,G29878);
  xor GNAME28198(G28198,G29962,G31429);
  and GNAME28199(G28199,G29962,G31429);
  xor GNAME28204(G28204,G29965,G31432);
  and GNAME28205(G28205,G29965,G31432);
  xor GNAME28210(G28210,G29968,G31435);
  and GNAME28211(G28211,G29968,G31435);
  xor GNAME28216(G28216,G31411,G31414);
  and GNAME28217(G28217,G31411,G31414);
  xor GNAME28222(G28222,G31417,G31420);
  and GNAME28223(G28223,G31417,G31420);
  xor GNAME28228(G28228,G31423,G31426);
  and GNAME28229(G28229,G31423,G31426);
  xor GNAME28234(G28234,G31719,G31628);
  and GNAME28235(G28235,G31719,G31628);
  xor GNAME28240(G28240,G31745,G31641);
  and GNAME28241(G28241,G31745,G31641);
  xor GNAME28246(G28246,G31732,G28235);
  and GNAME28247(G28247,G31732,G28235);
  xor GNAME28252(G28252,G31758,G28241);
  and GNAME28253(G28253,G31758,G28241);
  xor GNAME28258(G28258,G31823,G28247);
  and GNAME28259(G28259,G31823,G28247);
  xor GNAME28264(G28264,G31849,G28253);
  and GNAME28265(G28265,G31849,G28253);
  xor GNAME28270(G28270,G31836,G28259);
  and GNAME28271(G28271,G31836,G28259);
  xor GNAME28276(G28276,G31862,G28265);
  and GNAME28277(G28277,G31862,G28265);
  xor GNAME28282(G28282,G31953,G28271);
  and GNAME28283(G28283,G31953,G28271);
  xor GNAME28288(G28288,G31979,G28277);
  and GNAME28289(G28289,G31979,G28277);
  xor GNAME28294(G28294,G31966,G28283);
  and GNAME28295(G28295,G31966,G28283);
  xor GNAME28300(G28300,G31992,G28289);
  and GNAME28301(G28301,G31992,G28289);
  xor GNAME28306(G28306,G32083,G28295);
  and GNAME28307(G28307,G32083,G28295);
  xor GNAME28312(G28312,G32109,G28301);
  and GNAME28313(G28313,G32109,G28301);
  xor GNAME28318(G28318,G32096,G28307);
  and GNAME28319(G28319,G32096,G28307);
  xor GNAME28324(G28324,G32122,G28313);
  and GNAME28325(G28325,G32122,G28313);
  xor GNAME28330(G28330,G32226,G28355);
  and GNAME28331(G28331,G32226,G28355);
  xor GNAME28336(G28336,G32252,G28361);
  and GNAME28337(G28337,G32252,G28361);
  xor GNAME28342(G28342,G32343,G28331);
  and GNAME28343(G28343,G32343,G28331);
  xor GNAME28348(G28348,G32369,G28337);
  and GNAME28349(G28349,G32369,G28337);
  xor GNAME28354(G28354,G32213,G28319);
  and GNAME28355(G28355,G32213,G28319);
  xor GNAME28360(G28360,G32239,G28325);
  and GNAME28361(G28361,G32239,G28325);
  xor GNAME28366(G28366,G32356,G28343);
  and GNAME28367(G28367,G32356,G28343);
  xor GNAME28372(G28372,G32382,G28349);
  and GNAME28373(G28373,G32382,G28349);
  xor GNAME28378(G28378,G32473,G28367);
  and GNAME28379(G28379,G32473,G28367);
  xor GNAME28384(G28384,G32499,G28373);
  and GNAME28385(G28385,G32499,G28373);
  xor GNAME28390(G28390,G32486,G28379);
  and GNAME28391(G28391,G32486,G28379);
  xor GNAME28396(G28396,G32512,G28385);
  and GNAME28397(G28397,G32512,G28385);
  xor GNAME28402(G28402,G32603,G28391);
  and GNAME28403(G28403,G32603,G28391);
  xor GNAME28408(G28408,G32629,G28397);
  and GNAME28409(G28409,G32629,G28397);
  xor GNAME28414(G28414,G32616,G28403);
  and GNAME28415(G28415,G32616,G28403);
  xor GNAME28420(G28420,G32642,G28409);
  and GNAME28421(G28421,G32642,G28409);
  xor GNAME28426(G28426,G32733,G28415);
  and GNAME28427(G28427,G32733,G28415);
  xor GNAME28432(G28432,G32759,G28421);
  and GNAME28433(G28433,G32759,G28421);
  xor GNAME28438(G28438,G32746,G28427);
  and GNAME28439(G28439,G32746,G28427);
  xor GNAME28444(G28444,G32772,G28433);
  and GNAME28445(G28445,G32772,G28433);
  xor GNAME28450(G28450,G32876,G28439);
  and GNAME28451(G28451,G32876,G28439);
  xor GNAME28456(G28456,G32954,G28445);
  and GNAME28457(G28457,G32954,G28445);
  xor GNAME28462(G28462,G32889,G28451);
  and GNAME28463(G28463,G32889,G28451);
  xor GNAME28468(G28468,G32967,G28457);
  and GNAME28469(G28469,G32967,G28457);
  xor GNAME28474(G28474,G33058,G28463);
  and GNAME28475(G28475,G33058,G28463);
  xor GNAME28480(G28480,G33136,G28469);
  and GNAME28481(G28481,G33136,G28469);
  xor GNAME28486(G28486,G33071,G28475);
  and GNAME28487(G28487,G33071,G28475);
  xor GNAME28492(G28492,G33149,G28481);
  and GNAME28493(G28493,G33149,G28481);
  xor GNAME28498(G28498,G33253,G28487);
  and GNAME28499(G28499,G33253,G28487);
  xor GNAME28504(G28504,G33344,G28493);
  and GNAME28505(G28505,G33344,G28493);
  xor GNAME28510(G28510,G33266,G28499);
  and GNAME28511(G28511,G33266,G28499);
  xor GNAME28516(G28516,G33357,G28505);
  and GNAME28517(G28517,G33357,G28505);
  xor GNAME28522(G28522,G33448,G28511);
  and GNAME28523(G28523,G33448,G28511);
  xor GNAME28528(G28528,G33526,G28517);
  and GNAME28529(G28529,G33526,G28517);
  xor GNAME28534(G28534,G33461,G28523);
  and GNAME28535(G28535,G33461,G28523);
  xor GNAME28540(G28540,G33539,G28529);
  and GNAME28541(G28541,G33539,G28529);
  xor GNAME28546(G28546,G33630,G28535);
  and GNAME28547(G28547,G33630,G28535);
  xor GNAME28552(G28552,G33721,G28541);
  and GNAME28553(G28553,G33721,G28541);
  xor GNAME28558(G28558,G33643,G28547);
  and GNAME28559(G28559,G33643,G28547);
  xor GNAME28564(G28564,G33734,G28553);
  and GNAME28565(G28565,G33734,G28553);
  xor GNAME28570(G28570,G33825,G28559);
  and GNAME28571(G28571,G33825,G28559);
  xor GNAME28576(G28576,G33903,G28565);
  and GNAME28577(G28577,G33903,G28565);
  xor GNAME28582(G28582,G33838,G28571);
  and GNAME28583(G28583,G33838,G28571);
  xor GNAME28588(G28588,G33916,G28577);
  and GNAME28589(G28589,G33916,G28577);
  xor GNAME28594(G28594,G32902,G32863);
  and GNAME28595(G28595,G32902,G32863);
  xor GNAME28600(G28600,G34410,G28769);
  and GNAME28601(G28601,G34410,G28769);
  xor GNAME28606(G28606,G32915,G28595);
  and GNAME28607(G28607,G32915,G28595);
  xor GNAME28612(G28612,G32928,G28607);
  and GNAME28613(G28613,G32928,G28607);
  xor GNAME28618(G28618,G32941,G28613);
  and GNAME28619(G28619,G32941,G28613);
  xor GNAME28624(G28624,G33084,G28619);
  and GNAME28625(G28625,G33084,G28619);
  xor GNAME28630(G28630,G33097,G28625);
  and GNAME28631(G28631,G33097,G28625);
  xor GNAME28636(G28636,G33110,G28631);
  and GNAME28637(G28637,G33110,G28631);
  xor GNAME28642(G28642,G33123,G28637);
  and GNAME28643(G28643,G33123,G28637);
  xor GNAME28648(G28648,G33279,G28643);
  and GNAME28649(G28649,G33279,G28643);
  xor GNAME28654(G28654,G33292,G28649);
  and GNAME28655(G28655,G33292,G28649);
  xor GNAME28660(G28660,G33305,G28655);
  and GNAME28661(G28661,G33305,G28655);
  xor GNAME28666(G28666,G33318,G28661);
  and GNAME28667(G28667,G33318,G28661);
  xor GNAME28672(G28672,G33331,G28667);
  and GNAME28673(G28673,G33331,G28667);
  xor GNAME28678(G28678,G33474,G28673);
  and GNAME28679(G28679,G33474,G28673);
  xor GNAME28684(G28684,G33487,G28679);
  and GNAME28685(G28685,G33487,G28679);
  xor GNAME28690(G28690,G33500,G28685);
  and GNAME28691(G28691,G33500,G28685);
  xor GNAME28696(G28696,G33513,G28691);
  and GNAME28697(G28697,G33513,G28691);
  xor GNAME28702(G28702,G33656,G28697);
  and GNAME28703(G28703,G33656,G28697);
  xor GNAME28708(G28708,G33669,G28703);
  and GNAME28709(G28709,G33669,G28703);
  xor GNAME28714(G28714,G33682,G28709);
  and GNAME28715(G28715,G33682,G28709);
  xor GNAME28720(G28720,G33695,G28715);
  and GNAME28721(G28721,G33695,G28715);
  xor GNAME28726(G28726,G33708,G28721);
  and GNAME28727(G28727,G33708,G28721);
  xor GNAME28732(G28732,G33851,G28727);
  and GNAME28733(G28733,G33851,G28727);
  xor GNAME28738(G28738,G33864,G28733);
  and GNAME28739(G28739,G33864,G28733);
  xor GNAME28744(G28744,G33877,G28739);
  and GNAME28745(G28745,G33877,G28739);
  xor GNAME28750(G28750,G33890,G28745);
  and GNAME28751(G28751,G33890,G28745);
  xor GNAME28756(G28756,G34371,G28751);
  and GNAME28757(G28757,G34371,G28751);
  xor GNAME28762(G28762,G34384,G28757);
  and GNAME28763(G28763,G34384,G28757);
  xor GNAME28768(G28768,G34397,G28763);
  and GNAME28769(G28769,G34397,G28763);
  and GNAME28776(G28776,G27570,G28094);
  and GNAME28777(G28777,G29935,G27570);
  and GNAME28778(G28778,G28094,G29935);
  or GNAME28779(G28779,G28778,G28777,G28776);
  and GNAME28786(G28786,G27571,G28097);
  and GNAME28787(G28787,G29938,G27571);
  and GNAME28788(G28788,G28097,G29938);
  or GNAME28789(G28789,G28788,G28787,G28786);
  and GNAME28796(G28796,G27572,G28100);
  and GNAME28797(G28797,G29941,G27572);
  and GNAME28798(G28798,G28100,G29941);
  or GNAME28799(G28799,G28798,G28797,G28796);
  and GNAME28806(G28806,G28779,G31402);
  and GNAME28807(G28807,G28198,G28779);
  and GNAME28808(G28808,G31402,G28198);
  or GNAME28809(G28809,G28808,G28807,G28806);
  and GNAME28816(G28816,G28809,G28199);
  and GNAME28817(G28817,G17856,G28809);
  and GNAME28818(G28818,G28199,G17856);
  or GNAME28819(G28819,G28818,G28817,G28816);
  and GNAME28826(G28826,G28789,G31405);
  and GNAME28827(G28827,G28204,G28789);
  and GNAME28828(G28828,G31405,G28204);
  or GNAME28829(G28829,G28828,G28827,G28826);
  and GNAME28836(G28836,G28829,G28205);
  and GNAME28837(G28837,G17871,G28829);
  and GNAME28838(G28838,G28205,G17871);
  or GNAME28839(G28839,G28838,G28837,G28836);
  and GNAME28846(G28846,G28799,G31408);
  and GNAME28847(G28847,G28210,G28799);
  and GNAME28848(G28848,G31408,G28210);
  or GNAME28849(G28849,G28848,G28847,G28846);
  and GNAME28856(G28856,G28849,G28211);
  and GNAME28857(G28857,G17886,G28849);
  and GNAME28858(G28858,G28211,G17886);
  or GNAME28859(G28859,G28858,G28857,G28856);
  and GNAME28866(G28866,G28819,G17861);
  and GNAME28867(G28867,G17811,G28819);
  and GNAME28868(G28868,G17861,G17811);
  or GNAME28869(G28869,G28868,G28867,G28866);
  and GNAME28876(G28876,G28869,G17816);
  and GNAME28877(G28877,G21771,G28869);
  and GNAME28878(G28878,G17816,G21771);
  or GNAME28879(G28879,G28878,G28877,G28876);
  and GNAME28886(G28886,G28839,G17876);
  and GNAME28887(G28887,G17826,G28839);
  and GNAME28888(G28888,G17876,G17826);
  or GNAME28889(G28889,G28888,G28887,G28886);
  and GNAME28896(G28896,G28889,G17831);
  and GNAME28897(G28897,G21801,G28889);
  and GNAME28898(G28898,G17831,G21801);
  or GNAME28899(G28899,G28898,G28897,G28896);
  and GNAME28906(G28906,G28859,G17891);
  and GNAME28907(G28907,G17841,G28859);
  and GNAME28908(G28908,G17891,G17841);
  or GNAME28909(G28909,G28908,G28907,G28906);
  and GNAME28916(G28916,G28909,G17846);
  and GNAME28917(G28917,G21831,G28909);
  and GNAME28918(G28918,G17846,G21831);
  or GNAME28919(G28919,G28918,G28917,G28916);
  nor GNAME28920(G28920,G28990,G34725);
  nor GNAME28921(G28921,G34782,G31446);
  nor GNAME28922(G28922,G34783,G31447);
  nor GNAME28923(G28923,G34784,G31448);
  nor GNAME28924(G28924,G34783,G31449);
  nor GNAME28925(G28925,G34782,G31450);
  nor GNAME28926(G28926,G34784,G31451);
  nor GNAME28927(G28927,G34783,G31452);
  nor GNAME28928(G28928,G34782,G31453);
  nor GNAME28929(G28929,G34784,G31454);
  nor GNAME28930(G28930,G34783,G31455);
  nor GNAME28931(G28931,G34782,G31456);
  nor GNAME28932(G28932,G34784,G31457);
  nor GNAME28933(G28933,G34783,G31458);
  nor GNAME28934(G28934,G34782,G31459);
  nor GNAME28935(G28935,G34784,G31460);
  nor GNAME28936(G28936,G34783,G31461);
  nor GNAME28937(G28937,G34782,G31462);
  nor GNAME28938(G28938,G34784,G31463);
  nor GNAME28939(G28939,G34783,G31464);
  nor GNAME28940(G28940,G34782,G31465);
  nor GNAME28941(G28941,G34784,G31466);
  nor GNAME28942(G28942,G34783,G31467);
  nor GNAME28943(G28943,G34782,G31468);
  nor GNAME28944(G28944,G34784,G31469);
  nor GNAME28945(G28945,G34783,G31470);
  nor GNAME28946(G28946,G34782,G31471);
  nor GNAME28947(G28947,G34784,G31472);
  nor GNAME28948(G28948,G34783,G31473);
  nor GNAME28949(G28949,G34782,G31474);
  nor GNAME28950(G28950,G34784,G31475);
  nor GNAME28951(G28951,G34783,G31476);
  nor GNAME28952(G28952,G34782,G31477);
  nor GNAME28953(G28953,G34784,G31478);
  nor GNAME28954(G28954,G34785,G31482);
  nor GNAME28955(G28955,G34786,G31483);
  nor GNAME28956(G28956,G34787,G31484);
  nor GNAME28957(G28957,G34785,G31485);
  nor GNAME28958(G28958,G34786,G31486);
  nor GNAME28959(G28959,G34787,G31487);
  nor GNAME28960(G28960,G34785,G31488);
  nor GNAME28961(G28961,G34786,G31489);
  nor GNAME28962(G28962,G34787,G31490);
  nor GNAME28963(G28963,G34785,G31479);
  nor GNAME28964(G28964,G34786,G31480);
  nor GNAME28965(G28965,G34787,G31481);
  nor GNAME28966(G28966,G34785,G31491);
  nor GNAME28967(G28967,G34785,G31492);
  nor GNAME28968(G28968,G34786,G31493);
  nor GNAME28969(G28969,G34787,G31494);
  nor GNAME28970(G28970,G34786,G31495);
  nor GNAME28971(G28971,G34787,G31496);
  nor GNAME28972(G28972,G34785,G31497);
  nor GNAME28973(G28973,G34785,G31498);
  nor GNAME28974(G28974,G34786,G31499);
  nor GNAME28975(G28975,G34787,G31500);
  nor GNAME28976(G28976,G34786,G31501);
  nor GNAME28977(G28977,G34787,G31502);
  nor GNAME28978(G28978,G34785,G31503);
  nor GNAME28979(G28979,G34785,G31504);
  nor GNAME28980(G28980,G34786,G31505);
  nor GNAME28981(G28981,G34787,G31506);
  nor GNAME28982(G28982,G34786,G31507);
  nor GNAME28983(G28983,G34787,G31508);
  nor GNAME28984(G28984,G34785,G31509);
  nor GNAME28985(G28985,G34786,G31510);
  nor GNAME28986(G28986,G34787,G31511);
  nor GNAME28987(G28987,G34782,G31443);
  nor GNAME28988(G28988,G34783,G31444);
  nor GNAME28989(G28989,G34784,G31445);
  xnor GNAME28990(G28990,G31693,G2760);
  xnor GNAME28991(G28991,G2678,G2657);
  xnor GNAME28992(G28992,G2262,G2241);
  xnor GNAME28993(G28993,G1846,G1825);
  xnor GNAME28994(G28994,G2636,G2615);
  xnor GNAME28995(G28995,G2220,G2199);
  xnor GNAME28996(G28996,G1804,G1783);
  xnor GNAME28997(G28997,G2552,G2491);
  xnor GNAME28998(G28998,G2136,G2075);
  xnor GNAME28999(G28999,G1720,G1659);
  xnor GNAME29000(G29000,G2594,G2573);
  xnor GNAME29001(G29001,G2178,G2157);
  xnor GNAME29002(G29002,G1762,G1741);
  xnor GNAME29003(G29003,G2470,G2449);
  xnor GNAME29004(G29004,G2054,G2033);
  xnor GNAME29005(G29005,G1638,G1617);
  xnor GNAME29006(G29006,G2428,G2407);
  xnor GNAME29007(G29007,G2012,G1991);
  xnor GNAME29008(G29008,G1596,G1575);
  xnor GNAME29009(G29009,G2386,G2365);
  xnor GNAME29010(G29010,G1970,G1949);
  xnor GNAME29011(G29011,G1554,G1533);
  xnor GNAME29012(G29012,G34598,G34601);
  xnor GNAME29013(G29013,G34598,G34610);
  xnor GNAME29014(G29014,G34599,G34602);
  xnor GNAME29015(G29015,G34599,G34611);
  xnor GNAME29016(G29016,G34600,G34603);
  xnor GNAME29017(G29017,G34600,G34612);
  xnor GNAME29018(G29018,G34598,G34607);
  xnor GNAME29019(G29019,G34604,G34601);
  xnor GNAME29020(G29020,G34604,G34610);
  xnor GNAME29021(G29021,G34598,G34619);
  xnor GNAME29022(G29022,G34599,G34608);
  xnor GNAME29023(G29023,G34605,G34602);
  xnor GNAME29024(G29024,G34605,G34611);
  xnor GNAME29025(G29025,G34599,G34620);
  xnor GNAME29026(G29026,G34600,G34609);
  xnor GNAME29027(G29027,G34606,G34603);
  xnor GNAME29028(G29028,G34606,G34612);
  xnor GNAME29029(G29029,G34600,G34621);
  xnor GNAME29030(G29030,G34598,G34628);
  xnor GNAME29031(G29031,G34604,G34619);
  xnor GNAME29032(G29032,G34599,G34629);
  xnor GNAME29033(G29033,G34605,G34620);
  xnor GNAME29034(G29034,G34600,G34630);
  xnor GNAME29035(G29035,G34606,G34621);
  xnor GNAME29036(G29036,G34604,G34607);
  xnor GNAME29037(G29037,G34613,G34601);
  xnor GNAME29038(G29038,G34598,G34616);
  xnor GNAME29039(G29039,G34605,G34608);
  xnor GNAME29040(G29040,G34614,G34602);
  xnor GNAME29041(G29041,G34606,G34609);
  xnor GNAME29042(G29042,G34615,G34603);
  xnor GNAME29043(G29043,G34599,G34617);
  xnor GNAME29044(G29044,G34600,G34618);
  xnor GNAME29045(G29045,G34613,G34610);
  xnor GNAME29046(G29046,G34613,G34607);
  xnor GNAME29047(G29047,G34622,G34601);
  xnor GNAME29048(G29048,G34598,G34625);
  xnor GNAME29049(G29049,G34604,G34616);
  xnor GNAME29050(G29050,G34614,G34611);
  xnor GNAME29051(G29051,G34614,G34608);
  xnor GNAME29052(G29052,G34623,G34602);
  xnor GNAME29053(G29053,G34615,G34612);
  xnor GNAME29054(G29054,G34615,G34609);
  xnor GNAME29055(G29055,G34624,G34603);
  xnor GNAME29056(G29056,G34599,G34626);
  xnor GNAME29057(G29057,G34605,G34617);
  xnor GNAME29058(G29058,G34600,G34627);
  xnor GNAME29059(G29059,G34606,G34618);
  xnor GNAME29060(G29060,G34613,G34619);
  xnor GNAME29061(G29061,G34598,G34637);
  xnor GNAME29062(G29062,G34604,G34628);
  xnor GNAME29063(G29063,G34604,G34625);
  xnor GNAME29064(G29064,G34631,G34601);
  xnor GNAME29065(G29065,G34614,G34620);
  xnor GNAME29066(G29066,G34599,G34638);
  xnor GNAME29067(G29067,G34605,G34629);
  xnor GNAME29068(G29068,G34615,G34621);
  xnor GNAME29069(G29069,G34600,G34639);
  xnor GNAME29070(G29070,G34606,G34630);
  xnor GNAME29071(G29071,G34605,G34626);
  xnor GNAME29072(G29072,G34632,G34602);
  xnor GNAME29073(G29073,G34606,G34627);
  xnor GNAME29074(G29074,G34633,G34603);
  xnor GNAME29075(G29075,G34613,G34616);
  xnor GNAME29076(G29076,G34598,G34634);
  xnor GNAME29077(G29077,G34622,G34610);
  xnor GNAME29078(G29078,G34622,G34607);
  xnor GNAME29079(G29079,G34614,G34617);
  xnor GNAME29080(G29080,G34599,G34635);
  xnor GNAME29081(G29081,G34623,G34611);
  xnor GNAME29082(G29082,G34623,G34608);
  xnor GNAME29083(G29083,G34615,G34618);
  xnor GNAME29084(G29084,G34600,G34636);
  xnor GNAME29085(G29085,G34624,G34612);
  xnor GNAME29086(G29086,G34624,G34609);
  xnor GNAME29087(G29087,G34604,G34637);
  xnor GNAME29088(G29088,G34605,G34638);
  xnor GNAME29089(G29089,G34606,G34639);
  xnor GNAME29090(G29090,G34622,G34619);
  xnor GNAME29091(G29091,G34598,G34644);
  xnor GNAME29092(G29092,G34613,G34628);
  xnor GNAME29093(G29093,G34631,G34610);
  xnor GNAME29094(G29094,G34631,G34607);
  xnor GNAME29095(G29095,G34640,G34601);
  xnor GNAME29096(G29096,G34613,G34625);
  xnor GNAME29097(G29097,G34598,G34643);
  xnor GNAME29098(G29098,G34622,G34616);
  xnor GNAME29099(G29099,G34604,G34634);
  xnor GNAME29100(G29100,G34623,G34620);
  xnor GNAME29101(G29101,G34599,G34646);
  xnor GNAME29102(G29102,G34614,G34629);
  xnor GNAME29103(G29103,G34624,G34621);
  xnor GNAME29104(G29104,G34600,G34648);
  xnor GNAME29105(G29105,G34615,G34630);
  xnor GNAME29106(G29106,G34632,G34611);
  xnor GNAME29107(G29107,G34632,G34608);
  xnor GNAME29108(G29108,G34641,G34602);
  xnor GNAME29109(G29109,G34614,G34626);
  xnor GNAME29110(G29110,G34599,G34645);
  xnor GNAME29111(G29111,G34623,G34617);
  xnor GNAME29112(G29112,G34605,G34635);
  xnor GNAME29113(G29113,G34633,G34612);
  xnor GNAME29114(G29114,G34633,G34609);
  xnor GNAME29115(G29115,G34642,G34603);
  xnor GNAME29116(G29116,G34615,G34627);
  xnor GNAME29117(G29117,G34600,G34647);
  xnor GNAME29118(G29118,G34624,G34618);
  xnor GNAME29119(G29119,G34606,G34636);
  xnor GNAME29120(G29120,G34631,G34619);
  xnor GNAME29121(G29121,G34598,G34662);
  xnor GNAME29122(G29122,G34640,G34610);
  xnor GNAME29123(G29123,G34622,G34628);
  xnor GNAME29124(G29124,G34604,G34644);
  xnor GNAME29125(G29125,G34613,G34637);
  xnor GNAME29126(G29126,G34622,G34625);
  xnor GNAME29127(G29127,G34613,G34634);
  xnor GNAME29128(G29128,G34631,G34616);
  xnor GNAME29129(G29129,G34604,G34643);
  xnor GNAME29130(G29130,G34598,G34663);
  xnor GNAME29131(G29131,G34640,G34607);
  xnor GNAME29132(G29132,G34649,G34601);
  xnor GNAME29133(G29133,G34632,G34620);
  xnor GNAME29134(G29134,G34599,G34665);
  xnor GNAME29135(G29135,G34641,G34611);
  xnor GNAME29136(G29136,G34623,G34629);
  xnor GNAME29137(G29137,G34605,G34646);
  xnor GNAME29138(G29138,G34614,G34638);
  xnor GNAME29139(G29139,G34633,G34621);
  xnor GNAME29140(G29140,G34600,G34667);
  xnor GNAME29141(G29141,G34642,G34612);
  xnor GNAME29142(G29142,G34624,G34630);
  xnor GNAME29143(G29143,G34606,G34648);
  xnor GNAME29144(G29144,G34615,G34639);
  xnor GNAME29145(G29145,G34623,G34626);
  xnor GNAME29146(G29146,G34614,G34635);
  xnor GNAME29147(G29147,G34632,G34617);
  xnor GNAME29148(G29148,G34605,G34645);
  xnor GNAME29149(G29149,G34599,G34666);
  xnor GNAME29150(G29150,G34641,G34608);
  xnor GNAME29151(G29151,G34650,G34602);
  xnor GNAME29152(G29152,G34624,G34627);
  xnor GNAME29153(G29153,G34615,G34636);
  xnor GNAME29154(G29154,G34633,G34618);
  xnor GNAME29155(G29155,G34606,G34647);
  xnor GNAME29156(G29156,G34600,G34668);
  xnor GNAME29157(G29157,G34642,G34609);
  xnor GNAME29158(G29158,G34651,G34603);
  xnor GNAME29159(G29159,G34654,G34664);
  xnor GNAME29160(G29160,G34622,G34637);
  xnor GNAME29161(G29161,G34640,G34619);
  xnor GNAME29162(G29162,G34613,G34644);
  xnor GNAME29163(G29163,G34649,G34610);
  xnor GNAME29164(G29164,G34631,G34628);
  xnor GNAME29165(G29165,G34604,G34662);
  xnor GNAME29166(G29166,G34622,G34634);
  xnor GNAME29167(G29167,G34613,G34643);
  xnor GNAME29168(G29168,G34631,G34625);
  xnor GNAME29169(G29169,G34604,G34663);
  xnor GNAME29170(G29170,G34654,G34686);
  xnor GNAME29171(G29171,G34640,G34616);
  xnor GNAME29172(G29172,G34649,G34607);
  xnor GNAME29173(G29173,G34655,G34669);
  xnor GNAME29174(G29174,G34623,G34638);
  xnor GNAME29175(G29175,G34641,G34620);
  xnor GNAME29176(G29176,G34614,G34646);
  xnor GNAME29177(G29177,G34650,G34611);
  xnor GNAME29178(G29178,G34632,G34629);
  xnor GNAME29179(G29179,G34605,G34665);
  xnor GNAME29180(G29180,G34656,G34670);
  xnor GNAME29181(G29181,G34624,G34639);
  xnor GNAME29182(G29182,G34642,G34621);
  xnor GNAME29183(G29183,G34615,G34648);
  xnor GNAME29184(G29184,G34651,G34612);
  xnor GNAME29185(G29185,G34633,G34630);
  xnor GNAME29186(G29186,G34606,G34667);
  xnor GNAME29187(G29187,G34623,G34635);
  xnor GNAME29188(G29188,G34614,G34645);
  xnor GNAME29189(G29189,G34632,G34626);
  xnor GNAME29190(G29190,G34605,G34666);
  xnor GNAME29191(G29191,G34655,G34687);
  xnor GNAME29192(G29192,G34641,G34617);
  xnor GNAME29193(G29193,G34650,G34608);
  xnor GNAME29194(G29194,G34624,G34636);
  xnor GNAME29195(G29195,G34615,G34647);
  xnor GNAME29196(G29196,G34633,G34627);
  xnor GNAME29197(G29197,G34606,G34668);
  xnor GNAME29198(G29198,G34656,G34688);
  xnor GNAME29199(G29199,G34642,G34618);
  xnor GNAME29200(G29200,G34651,G34609);
  xnor GNAME29201(G29201,G34671,G34601);
  xnor GNAME29202(G29202,G34672,G34602);
  xnor GNAME29203(G29203,G34673,G34603);
  xnor GNAME29204(G29204,G34622,G34644);
  xnor GNAME29205(G29205,G34613,G34662);
  xnor GNAME29206(G29206,G34631,G34637);
  xnor GNAME29207(G29207,G34657,G34664);
  xnor GNAME29208(G29208,G34654,G34681);
  xnor GNAME29209(G29209,G34640,G34628);
  xnor GNAME29210(G29210,G34649,G34619);
  xnor GNAME29211(G29211,G34622,G34643);
  xnor GNAME29212(G29212,G34613,G34663);
  xnor GNAME29213(G29213,G34631,G34634);
  xnor GNAME29214(G29214,G34657,G34686);
  xnor GNAME29215(G29215,G34654,G34680);
  xnor GNAME29216(G29216,G34640,G34625);
  xnor GNAME29217(G29217,G34649,G34616);
  xnor GNAME29218(G29218,G34623,G34646);
  xnor GNAME29219(G29219,G34614,G34665);
  xnor GNAME29220(G29220,G34632,G34638);
  xnor GNAME29221(G29221,G34658,G34669);
  xnor GNAME29222(G29222,G34655,G34683);
  xnor GNAME29223(G29223,G34641,G34629);
  xnor GNAME29224(G29224,G34650,G34620);
  xnor GNAME29225(G29225,G34624,G34648);
  xnor GNAME29226(G29226,G34615,G34667);
  xnor GNAME29227(G29227,G34633,G34639);
  xnor GNAME29228(G29228,G34659,G34670);
  xnor GNAME29229(G29229,G34656,G34685);
  xnor GNAME29230(G29230,G34642,G34630);
  xnor GNAME29231(G29231,G34651,G34621);
  xnor GNAME29232(G29232,G34623,G34645);
  xnor GNAME29233(G29233,G34614,G34666);
  xnor GNAME29234(G29234,G34632,G34635);
  xnor GNAME29235(G29235,G34658,G34687);
  xnor GNAME29236(G29236,G34655,G34682);
  xnor GNAME29237(G29237,G34641,G34626);
  xnor GNAME29238(G29238,G34650,G34617);
  xnor GNAME29239(G29239,G34624,G34647);
  xnor GNAME29240(G29240,G34615,G34668);
  xnor GNAME29241(G29241,G34633,G34636);
  xnor GNAME29242(G29242,G34659,G34688);
  xnor GNAME29243(G29243,G34656,G34684);
  xnor GNAME29244(G29244,G34642,G34627);
  xnor GNAME29245(G29245,G34651,G34618);
  xnor GNAME29246(G29246,G34671,G34610);
  xnor GNAME29247(G29247,G34671,G34607);
  xnor GNAME29248(G29248,G34672,G34611);
  xnor GNAME29249(G29249,G34673,G34612);
  xnor GNAME29250(G29250,G34672,G34608);
  xnor GNAME29251(G29251,G34673,G34609);
  xnor GNAME29252(G29252,G34622,G34662);
  xnor GNAME29253(G29253,G34674,G34664);
  xnor GNAME29254(G29254,G34631,G34644);
  xnor GNAME29255(G29255,G34657,G34681);
  xnor GNAME29256(G29256,G34654,G34695);
  xnor GNAME29257(G29257,G34640,G34637);
  xnor GNAME29258(G29258,G34649,G34628);
  xnor GNAME29259(G29259,G34622,G34663);
  xnor GNAME29260(G29260,G34674,G34686);
  xnor GNAME29261(G29261,G34631,G34643);
  xnor GNAME29262(G29262,G34657,G34680);
  xnor GNAME29263(G29263,G34654,G34692);
  xnor GNAME29264(G29264,G34640,G34634);
  xnor GNAME29265(G29265,G34649,G34625);
  xnor GNAME29266(G29266,G34623,G34665);
  xnor GNAME29267(G29267,G34675,G34669);
  xnor GNAME29268(G29268,G34632,G34646);
  xnor GNAME29269(G29269,G34658,G34683);
  xnor GNAME29270(G29270,G34655,G34696);
  xnor GNAME29271(G29271,G34641,G34638);
  xnor GNAME29272(G29272,G34650,G34629);
  xnor GNAME29273(G29273,G34624,G34667);
  xnor GNAME29274(G29274,G34676,G34670);
  xnor GNAME29275(G29275,G34633,G34648);
  xnor GNAME29276(G29276,G34659,G34685);
  xnor GNAME29277(G29277,G34656,G34697);
  xnor GNAME29278(G29278,G34642,G34639);
  xnor GNAME29279(G29279,G34651,G34630);
  xnor GNAME29280(G29280,G34623,G34666);
  xnor GNAME29281(G29281,G34675,G34687);
  xnor GNAME29282(G29282,G34632,G34645);
  xnor GNAME29283(G29283,G34658,G34682);
  xnor GNAME29284(G29284,G34655,G34700);
  xnor GNAME29285(G29285,G34641,G34635);
  xnor GNAME29286(G29286,G34650,G34626);
  xnor GNAME29287(G29287,G34624,G34668);
  xnor GNAME29288(G29288,G34676,G34688);
  xnor GNAME29289(G29289,G34633,G34647);
  xnor GNAME29290(G29290,G34659,G34684);
  xnor GNAME29291(G29291,G34656,G34703);
  xnor GNAME29292(G29292,G34642,G34636);
  xnor GNAME29293(G29293,G34651,G34627);
  xnor GNAME29294(G29294,G34671,G34619);
  xnor GNAME29295(G29295,G34671,G34616);
  xnor GNAME29296(G29296,G34672,G34620);
  xnor GNAME29297(G29297,G34673,G34621);
  xnor GNAME29298(G29298,G34672,G34617);
  xnor GNAME29299(G29299,G34673,G34618);
  xnor GNAME29300(G29300,G34689,G34664);
  xnor GNAME29301(G29301,G34674,G34681);
  xnor GNAME29302(G29302,G34631,G34662);
  xnor GNAME29303(G29303,G34657,G34695);
  xnor GNAME29304(G29304,G34654,G34693);
  xnor GNAME29305(G29305,G34640,G34644);
  xnor GNAME29306(G29306,G34649,G34637);
  xnor GNAME29307(G29307,G34689,G34686);
  xnor GNAME29308(G29308,G34674,G34680);
  xnor GNAME29309(G29309,G34631,G34663);
  xnor GNAME29310(G29310,G34657,G34692);
  xnor GNAME29311(G29311,G34654,G34694);
  xnor GNAME29312(G29312,G34640,G34643);
  xnor GNAME29313(G29313,G34649,G34634);
  xnor GNAME29314(G29314,G34690,G34669);
  xnor GNAME29315(G29315,G34675,G34683);
  xnor GNAME29316(G29316,G34632,G34665);
  xnor GNAME29317(G29317,G34658,G34696);
  xnor GNAME29318(G29318,G34655,G34699);
  xnor GNAME29319(G29319,G34641,G34646);
  xnor GNAME29320(G29320,G34650,G34638);
  xnor GNAME29321(G29321,G34691,G34670);
  xnor GNAME29322(G29322,G34676,G34685);
  xnor GNAME29323(G29323,G34633,G34667);
  xnor GNAME29324(G29324,G34659,G34697);
  xnor GNAME29325(G29325,G34656,G34702);
  xnor GNAME29326(G29326,G34642,G34648);
  xnor GNAME29327(G29327,G34651,G34639);
  xnor GNAME29328(G29328,G34690,G34687);
  xnor GNAME29329(G29329,G34675,G34682);
  xnor GNAME29330(G29330,G34632,G34666);
  xnor GNAME29331(G29331,G34658,G34700);
  xnor GNAME29332(G29332,G34655,G34698);
  xnor GNAME29333(G29333,G34641,G34645);
  xnor GNAME29334(G29334,G34650,G34635);
  xnor GNAME29335(G29335,G34691,G34688);
  xnor GNAME29336(G29336,G34676,G34684);
  xnor GNAME29337(G29337,G34633,G34668);
  xnor GNAME29338(G29338,G34659,G34703);
  xnor GNAME29339(G29339,G34656,G34701);
  xnor GNAME29340(G29340,G34642,G34647);
  xnor GNAME29341(G29341,G34651,G34636);
  xnor GNAME29342(G29342,G34671,G34628);
  xnor GNAME29343(G29343,G34671,G34625);
  xnor GNAME29344(G29344,G34672,G34629);
  xnor GNAME29345(G29345,G34673,G34630);
  xnor GNAME29346(G29346,G34672,G34626);
  xnor GNAME29347(G29347,G34673,G34627);
  xnor GNAME29348(G29348,G34640,G34663);
  xnor GNAME29349(G29349,G34641,G34666);
  xnor GNAME29350(G29350,G34642,G34668);
  xnor GNAME29351(G29351,G34689,G34681);
  xnor GNAME29352(G29352,G34674,G34695);
  xnor GNAME29353(G29353,G34704,G34664);
  xnor GNAME29354(G29354,G34657,G34693);
  xnor GNAME29355(G29355,G34654,G34713);
  xnor GNAME29356(G29356,G34640,G34662);
  xnor GNAME29357(G29357,G34649,G34644);
  xnor GNAME29358(G29358,G34689,G34680);
  xnor GNAME29359(G29359,G34674,G34692);
  xnor GNAME29360(G29360,G34704,G34686);
  xnor GNAME29361(G29361,G34657,G34694);
  xnor GNAME29362(G29362,G34649,G34643);
  xnor GNAME29363(G29363,G34690,G34683);
  xnor GNAME29364(G29364,G34675,G34696);
  xnor GNAME29365(G29365,G34705,G34669);
  xnor GNAME29366(G29366,G34658,G34699);
  xnor GNAME29367(G29367,G34655,G34715);
  xnor GNAME29368(G29368,G34641,G34665);
  xnor GNAME29369(G29369,G34650,G34646);
  xnor GNAME29370(G29370,G34691,G34685);
  xnor GNAME29371(G29371,G34676,G34697);
  xnor GNAME29372(G29372,G34706,G34670);
  xnor GNAME29373(G29373,G34659,G34702);
  xnor GNAME29374(G29374,G34656,G34717);
  xnor GNAME29375(G29375,G34642,G34667);
  xnor GNAME29376(G29376,G34651,G34648);
  xnor GNAME29377(G29377,G34690,G34682);
  xnor GNAME29378(G29378,G34675,G34700);
  xnor GNAME29379(G29379,G34705,G34687);
  xnor GNAME29380(G29380,G34658,G34698);
  xnor GNAME29381(G29381,G34650,G34645);
  xnor GNAME29382(G29382,G34691,G34684);
  xnor GNAME29383(G29383,G34676,G34703);
  xnor GNAME29384(G29384,G34706,G34688);
  xnor GNAME29385(G29385,G34659,G34701);
  xnor GNAME29386(G29386,G34651,G34647);
  xnor GNAME29387(G29387,G34671,G34637);
  xnor GNAME29388(G29388,G34672,G34638);
  xnor GNAME29389(G29389,G34673,G34639);
  xnor GNAME29390(G29390,G34657,G34677);
  xnor GNAME29391(G29391,G34658,G34678);
  xnor GNAME29392(G29392,G34659,G34679);
  xnor GNAME29393(G29393,G34654,G34677);
  xnor GNAME29394(G29394,G34655,G34678);
  xnor GNAME29395(G29395,G34656,G34679);
  xnor GNAME29396(G29396,G34704,G34695);
  xnor GNAME29397(G29397,G34705,G34696);
  xnor GNAME29398(G29398,G34706,G34697);
  xnor GNAME29399(G29399,G34654,G34714);
  xnor GNAME29400(G29400,G34704,G34681);
  xnor GNAME29401(G29401,G34649,G34662);
  xnor GNAME29402(G29402,G34674,G34693);
  xnor GNAME29403(G29403,G34657,G34713);
  xnor GNAME29404(G29404,G34689,G34695);
  xnor GNAME29405(G29405,G34649,G34663);
  xnor GNAME29406(G29406,G34674,G34694);
  xnor GNAME29407(G29407,G34657,G34714);
  xnor GNAME29408(G29408,G34707,G34664);
  xnor GNAME29409(G29409,G34707,G34686);
  xnor GNAME29410(G29410,G34689,G34692);
  xnor GNAME29411(G29411,G34704,G34680);
  xnor GNAME29412(G29412,G34655,G34716);
  xnor GNAME29413(G29413,G34705,G34683);
  xnor GNAME29414(G29414,G34650,G34665);
  xnor GNAME29415(G29415,G34675,G34699);
  xnor GNAME29416(G29416,G34658,G34715);
  xnor GNAME29417(G29417,G34690,G34696);
  xnor GNAME29418(G29418,G34656,G34718);
  xnor GNAME29419(G29419,G34706,G34685);
  xnor GNAME29420(G29420,G34651,G34667);
  xnor GNAME29421(G29421,G34676,G34702);
  xnor GNAME29422(G29422,G34659,G34717);
  xnor GNAME29423(G29423,G34691,G34697);
  xnor GNAME29424(G29424,G34650,G34666);
  xnor GNAME29425(G29425,G34675,G34698);
  xnor GNAME29426(G29426,G34658,G34716);
  xnor GNAME29427(G29427,G34708,G34669);
  xnor GNAME29428(G29428,G34708,G34687);
  xnor GNAME29429(G29429,G34690,G34700);
  xnor GNAME29430(G29430,G34705,G34682);
  xnor GNAME29431(G29431,G34651,G34668);
  xnor GNAME29432(G29432,G34676,G34701);
  xnor GNAME29433(G29433,G34659,G34718);
  xnor GNAME29434(G29434,G34709,G34670);
  xnor GNAME29435(G29435,G34709,G34688);
  xnor GNAME29436(G29436,G34691,G34703);
  xnor GNAME29437(G29437,G34706,G34684);
  xnor GNAME29438(G29438,G34671,G34634);
  xnor GNAME29439(G29439,G34671,G34644);
  xnor GNAME29440(G29440,G34671,G34643);
  xnor GNAME29441(G29441,G34672,G34635);
  xnor GNAME29442(G29442,G34672,G34646);
  xnor GNAME29443(G29443,G34673,G34636);
  xnor GNAME29444(G29444,G34673,G34648);
  xnor GNAME29445(G29445,G34672,G34645);
  xnor GNAME29446(G29446,G34673,G34647);
  xnor GNAME29447(G29447,G34689,G34694);
  xnor GNAME29448(G29448,G34689,G34713);
  xnor GNAME29449(G29449,G34707,G34680);
  xnor GNAME29450(G29450,G34707,G34695);
  xnor GNAME29451(G29451,G34704,G34693);
  xnor GNAME29452(G29452,G34690,G34698);
  xnor GNAME29453(G29453,G34690,G34715);
  xnor GNAME29454(G29454,G34708,G34682);
  xnor GNAME29455(G29455,G34708,G34696);
  xnor GNAME29456(G29456,G34705,G34699);
  xnor GNAME29457(G29457,G34691,G34701);
  xnor GNAME29458(G29458,G34691,G34717);
  xnor GNAME29459(G29459,G34709,G34684);
  xnor GNAME29460(G29460,G34709,G34697);
  xnor GNAME29461(G29461,G34706,G34702);
  xnor GNAME29462(G29462,G34674,G34713);
  xnor GNAME29463(G29463,G34707,G34681);
  xnor GNAME29464(G29464,G34719,G34664);
  xnor GNAME29465(G29465,G34689,G34693);
  xnor GNAME29466(G29466,G34674,G34714);
  xnor GNAME29467(G29467,G34719,G34686);
  xnor GNAME29468(G29468,G34704,G34692);
  xnor GNAME29469(G29469,G34675,G34715);
  xnor GNAME29470(G29470,G34708,G34683);
  xnor GNAME29471(G29471,G34720,G34669);
  xnor GNAME29472(G29472,G34690,G34699);
  xnor GNAME29473(G29473,G34676,G34717);
  xnor GNAME29474(G29474,G34709,G34685);
  xnor GNAME29475(G29475,G34721,G34670);
  xnor GNAME29476(G29476,G34691,G34702);
  xnor GNAME29477(G29477,G34675,G34716);
  xnor GNAME29478(G29478,G34720,G34687);
  xnor GNAME29479(G29479,G34705,G34700);
  xnor GNAME29480(G29480,G34676,G34718);
  xnor GNAME29481(G29481,G34721,G34688);
  xnor GNAME29482(G29482,G34706,G34703);
  xnor GNAME29483(G29483,G34671,G34662);
  xnor GNAME29484(G29484,G34671,G34663);
  xnor GNAME29485(G29485,G34672,G34665);
  xnor GNAME29486(G29486,G34672,G34666);
  xnor GNAME29487(G29487,G34673,G34667);
  xnor GNAME29488(G29488,G34673,G34668);
  xnor GNAME29489(G29489,G34674,G34677);
  xnor GNAME29490(G29490,G34675,G34678);
  xnor GNAME29491(G29491,G34676,G34679);
  xnor GNAME29492(G29492,G34689,G34677);
  xnor GNAME29493(G29493,G34690,G34678);
  xnor GNAME29494(G29494,G34691,G34679);
  xnor GNAME29495(G29495,G34719,G34680);
  xnor GNAME29496(G29496,G34704,G34713);
  xnor GNAME29497(G29497,G34707,G34693);
  xnor GNAME29498(G29498,G34720,G34682);
  xnor GNAME29499(G29499,G34721,G34684);
  xnor GNAME29500(G29500,G34705,G34715);
  xnor GNAME29501(G29501,G34708,G34699);
  xnor GNAME29502(G29502,G34706,G34717);
  xnor GNAME29503(G29503,G34709,G34702);
  xnor GNAME29504(G29504,G34704,G34694);
  xnor GNAME29505(G29505,G34689,G34714);
  xnor GNAME29506(G29506,G34707,G34692);
  xnor GNAME29507(G29507,G34719,G34681);
  xnor GNAME29508(G29508,G34719,G34695);
  xnor GNAME29509(G29509,G34704,G34714);
  xnor GNAME29510(G29510,G34705,G34698);
  xnor GNAME29511(G29511,G34690,G34716);
  xnor GNAME29512(G29512,G34708,G34700);
  xnor GNAME29513(G29513,G34720,G34683);
  xnor GNAME29514(G29514,G34706,G34701);
  xnor GNAME29515(G29515,G34691,G34718);
  xnor GNAME29516(G29516,G34709,G34703);
  xnor GNAME29517(G29517,G34721,G34685);
  xnor GNAME29518(G29518,G34720,G34696);
  xnor GNAME29519(G29519,G34721,G34697);
  xnor GNAME29520(G29520,G34705,G34716);
  xnor GNAME29521(G29521,G34706,G34718);
  xnor GNAME29522(G29522,G34722,G34664);
  xnor GNAME29523(G29523,G34722,G34686);
  xnor GNAME29524(G29524,G34722,G34681);
  xnor GNAME29525(G29525,G34722,G34680);
  xnor GNAME29526(G29526,G34723,G34669);
  xnor GNAME29527(G29527,G34723,G34687);
  xnor GNAME29528(G29528,G34724,G34670);
  xnor GNAME29529(G29529,G34724,G34688);
  xnor GNAME29530(G29530,G34723,G34683);
  xnor GNAME29531(G29531,G34723,G34682);
  xnor GNAME29532(G29532,G34724,G34685);
  xnor GNAME29533(G29533,G34724,G34684);
  xnor GNAME29534(G29534,G34704,G34710);
  xnor GNAME29535(G29535,G34705,G34711);
  xnor GNAME29536(G29536,G34706,G34712);
  xnor GNAME29537(G29537,G34707,G34710);
  xnor GNAME29538(G29538,G34708,G34711);
  xnor GNAME29539(G29539,G34709,G34712);
  xnor GNAME29540(G29540,G34707,G34713);
  xnor GNAME29541(G29541,G34707,G34694);
  xnor GNAME29542(G29542,G34719,G34692);
  xnor GNAME29543(G29543,G34719,G34693);
  xnor GNAME29544(G29544,G34708,G34698);
  xnor GNAME29545(G29545,G34708,G34715);
  xnor GNAME29546(G29546,G34720,G34700);
  xnor GNAME29547(G29547,G34720,G34699);
  xnor GNAME29548(G29548,G34709,G34701);
  xnor GNAME29549(G29549,G34709,G34717);
  xnor GNAME29550(G29550,G34721,G34703);
  xnor GNAME29551(G29551,G34721,G34702);
  xnor GNAME29552(G29552,G34719,G34694);
  xnor GNAME29553(G29553,G34707,G34714);
  xnor GNAME29554(G29554,G34720,G34698);
  xnor GNAME29555(G29555,G34708,G34716);
  xnor GNAME29556(G29556,G34721,G34701);
  xnor GNAME29557(G29557,G34709,G34718);
  xnor GNAME29558(G29558,G34722,G34692);
  xnor GNAME29559(G29559,G34722,G34695);
  xnor GNAME29560(G29560,G34723,G34696);
  xnor GNAME29561(G29561,G34724,G34697);
  xnor GNAME29562(G29562,G34723,G34700);
  xnor GNAME29563(G29563,G34724,G34703);
  xnor GNAME29564(G29564,G34719,G34713);
  xnor GNAME29565(G29565,G34719,G34714);
  xnor GNAME29566(G29566,G34720,G34715);
  xnor GNAME29567(G29567,G34720,G34716);
  xnor GNAME29568(G29568,G34721,G34717);
  xnor GNAME29569(G29569,G34721,G34718);
  xnor GNAME29570(G29570,G34722,G34693);
  xnor GNAME29571(G29571,G34722,G34694);
  xnor GNAME29572(G29572,G34723,G34699);
  xnor GNAME29573(G29573,G34723,G34698);
  xnor GNAME29574(G29574,G34724,G34702);
  xnor GNAME29575(G29575,G34724,G34701);
  xnor GNAME29576(G29576,G34722,G34713);
  xnor GNAME29577(G29577,G34722,G34714);
  xnor GNAME29578(G29578,G34723,G34715);
  xnor GNAME29579(G29579,G34723,G34716);
  xnor GNAME29580(G29580,G34724,G34717);
  xnor GNAME29581(G29581,G34724,G34718);
  xnor GNAME29582(G29582,G34722,G34710);
  xnor GNAME29583(G29583,G34723,G34711);
  xnor GNAME29584(G29584,G34724,G34712);
  xnor GNAME29585(G29585,G34719,G34710);
  xnor GNAME29586(G29586,G34720,G34711);
  xnor GNAME29587(G29587,G34721,G34712);
  and GNAME29588(G29588,G34795,G34727);
  or GNAME29589(G29589,G31512,G29588);
  and GNAME29590(G29590,G34794,G34726);
  or GNAME29591(G29591,G31513,G29590);
  and GNAME29592(G29592,G34796,G34728);
  or GNAME29593(G29593,G31514,G29592);
  and GNAME29594(G29594,G34800,G34734);
  or GNAME29595(G29595,G31515,G29594);
  and GNAME29596(G29596,G34801,G34735);
  or GNAME29597(G29597,G31516,G29596);
  and GNAME29598(G29598,G34802,G34736);
  or GNAME29599(G29599,G31517,G29598);
  and GNAME29600(G29600,G34749,G34740);
  or GNAME29601(G29601,G31520,G29600);
  and GNAME29602(G29602,G34751,G34742);
  or GNAME29603(G29603,G31522,G29602);
  and GNAME29604(G29604,G34752,G34743);
  or GNAME29605(G29605,G31523,G29604);
  and GNAME29606(G29606,G34750,G34741);
  or GNAME29607(G29607,G31521,G29606);
  and GNAME29608(G29608,G34753,G34744);
  or GNAME29609(G29609,G31524,G29608);
  and GNAME29610(G29610,G34754,G34745);
  or GNAME29611(G29611,G31525,G29610);
  and GNAME29612(G29612,G34827,G34803);
  or GNAME29613(G29613,G31526,G29612);
  and GNAME29614(G29614,G34828,G34804);
  or GNAME29615(G29615,G31527,G29614);
  and GNAME29616(G29616,G34829,G34805);
  or GNAME29617(G29617,G31528,G29616);
  and GNAME29618(G29618,G34824,G34806);
  or GNAME29619(G29619,G31532,G29618);
  and GNAME29620(G29620,G34825,G34807);
  or GNAME29621(G29621,G31529,G29620);
  and GNAME29622(G29622,G34826,G34808);
  or GNAME29623(G29623,G31530,G29622);
  and GNAME29624(G29624,G34779,G34761);
  or GNAME29625(G29625,G31531,G29624);
  and GNAME29626(G29626,G34780,G34762);
  or GNAME29627(G29627,G31533,G29626);
  and GNAME29628(G29628,G34781,G34763);
  or GNAME29629(G29629,G31534,G29628);
  and GNAME29630(G29630,G34764,G34758);
  or GNAME29631(G29631,G31535,G29630);
  and GNAME29632(G29632,G34765,G34759);
  or GNAME29633(G29633,G31536,G29632);
  and GNAME29634(G29634,G34766,G34760);
  or GNAME29635(G29635,G31537,G29634);
  or GNAME29636(G29636,G34794,G29012);
  or GNAME29637(G29637,G34726,G29013);
  nand GNAME29638(G29638,G29637,G29636);
  or GNAME29639(G29639,G34795,G29014);
  or GNAME29640(G29640,G34727,G29015);
  nand GNAME29641(G29641,G29640,G29639);
  or GNAME29642(G29642,G34796,G29016);
  or GNAME29643(G29643,G34728,G29017);
  nand GNAME29644(G29644,G29643,G29642);
  or GNAME29645(G29645,G34800,G29019);
  or GNAME29646(G29646,G34734,G29020);
  nand GNAME29647(G29647,G29646,G29645);
  or GNAME29648(G29648,G34801,G29023);
  or GNAME29649(G29649,G34735,G29024);
  nand GNAME29650(G29650,G29649,G29648);
  or GNAME29651(G29651,G34802,G29027);
  or GNAME29652(G29652,G34736,G29028);
  nand GNAME29653(G29653,G29652,G29651);
  or GNAME29654(G29654,G34749,G29037);
  or GNAME29655(G29655,G34740,G29045);
  nand GNAME29656(G29656,G29655,G29654);
  or GNAME29657(G29657,G34751,G29040);
  or GNAME29658(G29658,G34742,G29050);
  nand GNAME29659(G29659,G29658,G29657);
  or GNAME29660(G29660,G34752,G29042);
  or GNAME29661(G29661,G34743,G29053);
  nand GNAME29662(G29662,G29661,G29660);
  or GNAME29663(G29663,G34749,G29046);
  or GNAME29664(G29664,G34740,G29060);
  nand GNAME29665(G29665,G29664,G29663);
  or GNAME29666(G29666,G34751,G29051);
  or GNAME29667(G29667,G34742,G29065);
  nand GNAME29668(G29668,G29667,G29666);
  or GNAME29669(G29669,G34752,G29054);
  or GNAME29670(G29670,G34743,G29068);
  nand GNAME29671(G29671,G29670,G29669);
  or GNAME29672(G29672,G34750,G29078);
  or GNAME29673(G29673,G34741,G29090);
  nand GNAME29674(G29674,G29673,G29672);
  or GNAME29675(G29675,G34753,G29082);
  or GNAME29676(G29676,G34744,G29100);
  nand GNAME29677(G29677,G29676,G29675);
  or GNAME29678(G29678,G34754,G29086);
  or GNAME29679(G29679,G34745,G29103);
  nand GNAME29680(G29680,G29679,G29678);
  or GNAME29681(G29681,G34750,G29098);
  or GNAME29682(G29682,G34741,G29123);
  nand GNAME29683(G29683,G29682,G29681);
  or GNAME29684(G29684,G34753,G29111);
  or GNAME29685(G29685,G34744,G29136);
  nand GNAME29686(G29686,G29685,G29684);
  or GNAME29687(G29687,G34754,G29118);
  or GNAME29688(G29688,G34745,G29142);
  nand GNAME29689(G29689,G29688,G29687);
  or GNAME29690(G29690,G34779,G31531);
  or GNAME29691(G29691,G34761,G29132);
  nand GNAME29692(G29692,G29691,G29690);
  or GNAME29693(G29693,G34780,G31533);
  or GNAME29694(G29694,G34762,G29151);
  nand GNAME29695(G29695,G29694,G29693);
  or GNAME29696(G29696,G34781,G31534);
  or GNAME29697(G29697,G34763,G29158);
  nand GNAME29698(G29698,G29697,G29696);
  or GNAME29699(G29699,G34779,G29357);
  or GNAME29700(G29700,G34761,G29362);
  nand GNAME29701(G29701,G29700,G29699);
  or GNAME29702(G29702,G29387,G34764);
  or GNAME29703(G29703,G34758,G29438);
  nand GNAME29704(G29704,G29703,G29702);
  or GNAME29705(G29705,G34780,G29369);
  or GNAME29706(G29706,G34762,G29381);
  nand GNAME29707(G29707,G29706,G29705);
  or GNAME29708(G29708,G29388,G34765);
  or GNAME29709(G29709,G34759,G29441);
  nand GNAME29710(G29710,G29709,G29708);
  or GNAME29711(G29711,G34781,G29376);
  or GNAME29712(G29712,G34763,G29386);
  nand GNAME29713(G29713,G29712,G29711);
  or GNAME29714(G29714,G29389,G34766);
  or GNAME29715(G29715,G34760,G29443);
  nand GNAME29716(G29716,G29715,G29714);
  or GNAME29717(G29717,G34774,G29401);
  or GNAME29718(G29718,G34770,G29405);
  nand GNAME29719(G29719,G29718,G29717);
  or GNAME29720(G29720,G29439,G34764);
  or GNAME29721(G29721,G34758,G29440);
  nand GNAME29722(G29722,G29721,G29720);
  or GNAME29723(G29723,G34776,G29414);
  or GNAME29724(G29724,G34771,G29424);
  nand GNAME29725(G29725,G29724,G29723);
  or GNAME29726(G29726,G29442,G34765);
  or GNAME29727(G29727,G34759,G29445);
  nand GNAME29728(G29728,G29727,G29726);
  or GNAME29729(G29729,G34778,G29420);
  or GNAME29730(G29730,G34772,G29431);
  nand GNAME29731(G29731,G29730,G29729);
  or GNAME29732(G29732,G29444,G34766);
  or GNAME29733(G29733,G34760,G29446);
  nand GNAME29734(G29734,G29733,G29732);
  or GNAME29735(G29735,G34737,G29407);
  or GNAME29736(G29736,G34789,G29390);
  nand GNAME29737(G29737,G29736,G29735);
  or GNAME29738(G29738,G29440,G34764);
  or GNAME29739(G29739,G34767,G29483);
  nand GNAME29740(G29740,G29739,G29738);
  or GNAME29741(G29741,G34738,G29426);
  or GNAME29742(G29742,G34792,G29391);
  nand GNAME29743(G29743,G29742,G29741);
  or GNAME29744(G29744,G29445,G34765);
  or GNAME29745(G29745,G34768,G29485);
  nand GNAME29746(G29746,G29745,G29744);
  or GNAME29747(G29747,G34739,G29433);
  or GNAME29748(G29748,G34793,G29392);
  nand GNAME29749(G29749,G29748,G29747);
  or GNAME29750(G29750,G29446,G34766);
  or GNAME29751(G29751,G34769,G29487);
  nand GNAME29752(G29752,G29751,G29750);
  or GNAME29753(G29753,G34731,G29399);
  or GNAME29754(G29754,G34788,G29393);
  nand GNAME29755(G29755,G29754,G29753);
  or GNAME29756(G29756,G29438,G34764);
  or GNAME29757(G29757,G34758,G29439);
  nand GNAME29758(G29758,G29757,G29756);
  or GNAME29759(G29759,G34732,G29412);
  or GNAME29760(G29760,G34790,G29394);
  nand GNAME29761(G29761,G29760,G29759);
  or GNAME29762(G29762,G29441,G34765);
  or GNAME29763(G29763,G34759,G29442);
  nand GNAME29764(G29764,G29763,G29762);
  or GNAME29765(G29765,G34733,G29418);
  or GNAME29766(G29766,G34791,G29395);
  nand GNAME29767(G29767,G29766,G29765);
  or GNAME29768(G29768,G29443,G34766);
  or GNAME29769(G29769,G34760,G29444);
  nand GNAME29770(G29770,G29769,G29768);
  or GNAME29771(G29771,G34774,G29464);
  or GNAME29772(G29772,G34770,G29467);
  nand GNAME29773(G29773,G29772,G29771);
  or GNAME29774(G29774,G29483,G34755);
  or GNAME29775(G29775,G34767,G29484);
  nand GNAME29776(G29776,G29775,G29774);
  or GNAME29777(G29777,G34776,G29471);
  or GNAME29778(G29778,G34771,G29478);
  nand GNAME29779(G29779,G29778,G29777);
  or GNAME29780(G29780,G29485,G34756);
  or GNAME29781(G29781,G34768,G29486);
  nand GNAME29782(G29782,G29781,G29780);
  or GNAME29783(G29783,G34778,G29475);
  or GNAME29784(G29784,G34772,G29481);
  nand GNAME29785(G29785,G29784,G29783);
  or GNAME29786(G29786,G29487,G34757);
  or GNAME29787(G29787,G34769,G29488);
  nand GNAME29788(G29788,G29787,G29786);
  or GNAME29789(G29789,G34746,G29466);
  or GNAME29790(G29790,G34797,G29489);
  nand GNAME29791(G29791,G29790,G29789);
  or GNAME29792(G29792,G29484,G34755);
  or GNAME29793(G29793,G34767,G29522);
  nand GNAME29794(G29794,G29793,G29792);
  or GNAME29795(G29795,G34747,G29477);
  or GNAME29796(G29796,G34798,G29490);
  nand GNAME29797(G29797,G29796,G29795);
  or GNAME29798(G29798,G29486,G34756);
  or GNAME29799(G29799,G34768,G29526);
  nand GNAME29800(G29800,G29799,G29798);
  or GNAME29801(G29801,G34748,G29480);
  or GNAME29802(G29802,G34799,G29491);
  nand GNAME29803(G29803,G29802,G29801);
  or GNAME29804(G29804,G29488,G34757);
  or GNAME29805(G29805,G34769,G29528);
  nand GNAME29806(G29806,G29805,G29804);
  or GNAME29807(G29807,G34774,G29507);
  or GNAME29808(G29808,G34770,G29495);
  nand GNAME29809(G29809,G29808,G29807);
  or GNAME29810(G29810,G29522,G34755);
  or GNAME29811(G29811,G34767,G29523);
  nand GNAME29812(G29812,G29811,G29810);
  or GNAME29813(G29813,G34776,G29513);
  or GNAME29814(G29814,G34771,G29498);
  nand GNAME29815(G29815,G29814,G29813);
  or GNAME29816(G29816,G29526,G34756);
  or GNAME29817(G29817,G34768,G29527);
  nand GNAME29818(G29818,G29817,G29816);
  or GNAME29819(G29819,G34778,G29517);
  or GNAME29820(G29820,G34772,G29499);
  nand GNAME29821(G29821,G29820,G29819);
  or GNAME29822(G29822,G29528,G34757);
  or GNAME29823(G29823,G34769,G29529);
  nand GNAME29824(G29824,G29823,G29822);
  or GNAME29825(G29825,G34809,G29505);
  or GNAME29826(G29826,G34815,G29492);
  nand GNAME29827(G29827,G29826,G29825);
  or GNAME29828(G29828,G29523,G34755);
  or GNAME29829(G29829,G34767,G29524);
  nand GNAME29830(G29830,G29829,G29828);
  or GNAME29831(G29831,G34810,G29511);
  or GNAME29832(G29832,G34816,G29493);
  nand GNAME29833(G29833,G29832,G29831);
  or GNAME29834(G29834,G29527,G34756);
  or GNAME29835(G29835,G34768,G29530);
  nand GNAME29836(G29836,G29835,G29834);
  or GNAME29837(G29837,G34811,G29515);
  or GNAME29838(G29838,G34817,G29494);
  nand GNAME29839(G29839,G29838,G29837);
  or GNAME29840(G29840,G29529,G34757);
  or GNAME29841(G29841,G34769,G29532);
  nand GNAME29842(G29842,G29841,G29840);
  or GNAME29843(G29843,G34774,G29508);
  or GNAME29844(G29844,G34770,G29542);
  nand GNAME29845(G29845,G29844,G29843);
  or GNAME29846(G29846,G29524,G34755);
  or GNAME29847(G29847,G34767,G29525);
  nand GNAME29848(G29848,G29847,G29846);
  or GNAME29849(G29849,G34776,G29518);
  or GNAME29850(G29850,G34771,G29546);
  nand GNAME29851(G29851,G29850,G29849);
  or GNAME29852(G29852,G29530,G34756);
  or GNAME29853(G29853,G34768,G29531);
  nand GNAME29854(G29854,G29853,G29852);
  or GNAME29855(G29855,G34778,G29519);
  or GNAME29856(G29856,G34772,G29550);
  nand GNAME29857(G29857,G29856,G29855);
  or GNAME29858(G29858,G29532,G34757);
  or GNAME29859(G29859,G34769,G29533);
  nand GNAME29860(G29860,G29859,G29858);
  or GNAME29861(G29861,G34812,G29509);
  or GNAME29862(G29862,G34821,G29534);
  nand GNAME29863(G29863,G29862,G29861);
  or GNAME29864(G29864,G29525,G34755);
  or GNAME29865(G29865,G34767,G29559);
  nand GNAME29866(G29866,G29865,G29864);
  or GNAME29867(G29867,G34813,G29520);
  or GNAME29868(G29868,G34822,G29535);
  nand GNAME29869(G29869,G29868,G29867);
  or GNAME29870(G29870,G29531,G34756);
  or GNAME29871(G29871,G34768,G29560);
  nand GNAME29872(G29872,G29871,G29870);
  or GNAME29873(G29873,G34814,G29521);
  or GNAME29874(G29874,G34823,G29536);
  nand GNAME29875(G29875,G29874,G29873);
  or GNAME29876(G29876,G29533,G34757);
  or GNAME29877(G29877,G34769,G29561);
  nand GNAME29878(G29878,G29877,G29876);
  or GNAME29879(G29879,G34774,G29543);
  or GNAME29880(G29880,G34770,G29552);
  nand GNAME29881(G29881,G29880,G29879);
  or GNAME29882(G29882,G29559,G34755);
  or GNAME29883(G29883,G34767,G29558);
  nand GNAME29884(G29884,G29883,G29882);
  or GNAME29885(G29885,G34776,G29547);
  or GNAME29886(G29886,G34771,G29554);
  nand GNAME29887(G29887,G29886,G29885);
  or GNAME29888(G29888,G29560,G34756);
  or GNAME29889(G29889,G34768,G29562);
  nand GNAME29890(G29890,G29889,G29888);
  or GNAME29891(G29891,G34778,G29551);
  or GNAME29892(G29892,G34772,G29556);
  nand GNAME29893(G29893,G29892,G29891);
  or GNAME29894(G29894,G29561,G34757);
  or GNAME29895(G29895,G34769,G29563);
  nand GNAME29896(G29896,G29895,G29894);
  or GNAME29897(G29897,G34773,G29553);
  or GNAME29898(G29898,G34818,G29537);
  nand GNAME29899(G29899,G29898,G29897);
  or GNAME29900(G29900,G34824,G27915);
  or GNAME29901(G29901,G34806,G31532);
  nand GNAME29902(G29902,G29901,G29900);
  or GNAME29903(G29903,G34775,G29555);
  or GNAME29904(G29904,G34819,G29538);
  nand GNAME29905(G29905,G29904,G29903);
  or GNAME29906(G29906,G34825,G27918);
  or GNAME29907(G29907,G34807,G31529);
  nand GNAME29908(G29908,G29907,G29906);
  or GNAME29909(G29909,G34777,G29557);
  or GNAME29910(G29910,G34820,G29539);
  nand GNAME29911(G29911,G29910,G29909);
  or GNAME29912(G29912,G34826,G27921);
  or GNAME29913(G29913,G34808,G31530);
  nand GNAME29914(G29914,G29913,G29912);
  or GNAME29915(G29915,G34774,G29564);
  or GNAME29916(G29916,G34770,G29565);
  nand GNAME29917(G29917,G29916,G29915);
  or GNAME29918(G29918,G29570,G34755);
  or GNAME29919(G29919,G34767,G29571);
  nand GNAME29920(G29920,G29919,G29918);
  or GNAME29921(G29921,G34776,G29566);
  or GNAME29922(G29922,G34771,G29567);
  nand GNAME29923(G29923,G29922,G29921);
  or GNAME29924(G29924,G29572,G34756);
  or GNAME29925(G29925,G34768,G29573);
  nand GNAME29926(G29926,G29925,G29924);
  or GNAME29927(G29927,G34778,G29568);
  or GNAME29928(G29928,G34772,G29569);
  nand GNAME29929(G29929,G29928,G29927);
  or GNAME29930(G29930,G29574,G34757);
  or GNAME29931(G29931,G34769,G29575);
  nand GNAME29932(G29932,G29931,G29930);
  or GNAME29933(G29933,G29576,G34755);
  or GNAME29934(G29934,G34767,G29577);
  nand GNAME29935(G29935,G29934,G29933);
  or GNAME29936(G29936,G29578,G34756);
  or GNAME29937(G29937,G34768,G29579);
  nand GNAME29938(G29938,G29937,G29936);
  or GNAME29939(G29939,G29580,G34757);
  or GNAME29940(G29940,G34769,G29581);
  nand GNAME29941(G29941,G29940,G29939);
  or GNAME29942(G29942,G29577,G34755);
  or GNAME29943(G29943,G34767,G29582);
  nand GNAME29944(G29944,G29943,G29942);
  or GNAME29945(G29945,G29579,G34756);
  or GNAME29946(G29946,G34768,G29583);
  nand GNAME29947(G29947,G29946,G29945);
  or GNAME29948(G29948,G29581,G34757);
  or GNAME29949(G29949,G34769,G29584);
  nand GNAME29950(G29950,G29949,G29948);
  or GNAME29951(G29951,G27924,G34764);
  or GNAME29952(G29952,G34758,G31535);
  nand GNAME29953(G29953,G29952,G29951);
  or GNAME29954(G29954,G27927,G34765);
  or GNAME29955(G29955,G34759,G31536);
  nand GNAME29956(G29956,G29955,G29954);
  or GNAME29957(G29957,G27930,G34766);
  or GNAME29958(G29958,G34760,G31537);
  nand GNAME29959(G29959,G29958,G29957);
  or GNAME29960(G29960,G34774,G29565);
  or GNAME29961(G29961,G34770,G29585);
  nand GNAME29962(G29962,G29961,G29960);
  or GNAME29963(G29963,G34776,G29567);
  or GNAME29964(G29964,G34771,G29586);
  nand GNAME29965(G29965,G29964,G29963);
  or GNAME29966(G29966,G34778,G29569);
  or GNAME29967(G29967,G34772,G29587);
  nand GNAME29968(G29968,G29967,G29966);
  or GNAME29969(G29969,G34794,G31513);
  or GNAME29970(G29970,G34726,G29012);
  nand GNAME29971(G29971,G29970,G29969);
  or GNAME29972(G29972,G34795,G31512);
  or GNAME29973(G29973,G34727,G29014);
  nand GNAME29974(G29974,G29973,G29972);
  or GNAME29975(G29975,G34796,G31514);
  or GNAME29976(G29976,G34728,G29016);
  nand GNAME29977(G29977,G29976,G29975);
  or GNAME29978(G29978,G34800,G31515);
  or GNAME29979(G29979,G34734,G29019);
  nand GNAME29980(G29980,G29979,G29978);
  or GNAME29981(G29981,G34794,G29013);
  or GNAME29982(G29982,G34726,G29018);
  nand GNAME29983(G29983,G29982,G29981);
  or GNAME29984(G29984,G34801,G31516);
  or GNAME29985(G29985,G34735,G29023);
  nand GNAME29986(G29986,G29985,G29984);
  or GNAME29987(G29987,G34795,G29015);
  or GNAME29988(G29988,G34727,G29022);
  nand GNAME29989(G29989,G29988,G29987);
  or GNAME29990(G29990,G34802,G31517);
  or GNAME29991(G29991,G34736,G29027);
  nand GNAME29992(G29992,G29991,G29990);
  or GNAME29993(G29993,G34796,G29017);
  or GNAME29994(G29994,G34728,G29026);
  nand GNAME29995(G29995,G29994,G29993);
  or GNAME29996(G29996,G34794,G29018);
  or GNAME29997(G29997,G34726,G29021);
  nand GNAME29998(G29998,G29997,G29996);
  or GNAME29999(G29999,G34795,G29022);
  or GNAME30000(G30000,G34727,G29025);
  nand GNAME30001(G30001,G30000,G29999);
  or GNAME30002(G30002,G34796,G29026);
  or GNAME30003(G30003,G34728,G29029);
  nand GNAME30004(G30004,G30003,G30002);
  or GNAME30005(G30005,G34794,G29021);
  or GNAME30006(G30006,G34726,G29038);
  nand GNAME30007(G30007,G30006,G30005);
  or GNAME30008(G30008,G34795,G29025);
  or GNAME30009(G30009,G34727,G29043);
  nand GNAME30010(G30010,G30009,G30008);
  or GNAME30011(G30011,G34796,G29029);
  or GNAME30012(G30012,G34728,G29044);
  nand GNAME30013(G30013,G30012,G30011);
  or GNAME30014(G30014,G34749,G31520);
  or GNAME30015(G30015,G34740,G29037);
  nand GNAME30016(G30016,G30015,G30014);
  or GNAME30017(G30017,G34800,G29020);
  or GNAME30018(G30018,G34734,G29036);
  nand GNAME30019(G30019,G30018,G30017);
  or GNAME30020(G30020,G34751,G31522);
  or GNAME30021(G30021,G34742,G29040);
  nand GNAME30022(G30022,G30021,G30020);
  or GNAME30023(G30023,G34801,G29024);
  or GNAME30024(G30024,G34735,G29039);
  nand GNAME30025(G30025,G30024,G30023);
  or GNAME30026(G30026,G34752,G31523);
  or GNAME30027(G30027,G34743,G29042);
  nand GNAME30028(G30028,G30027,G30026);
  or GNAME30029(G30029,G34802,G29028);
  or GNAME30030(G30030,G34736,G29041);
  nand GNAME30031(G30031,G30030,G30029);
  or GNAME30032(G30032,G34794,G29038);
  or GNAME30033(G30033,G34726,G29030);
  nand GNAME30034(G30034,G30033,G30032);
  or GNAME30035(G30035,G34800,G29036);
  or GNAME30036(G30036,G34734,G29031);
  nand GNAME30037(G30037,G30036,G30035);
  or GNAME30038(G30038,G34795,G29043);
  or GNAME30039(G30039,G34727,G29032);
  nand GNAME30040(G30040,G30039,G30038);
  or GNAME30041(G30041,G34801,G29039);
  or GNAME30042(G30042,G34735,G29033);
  nand GNAME30043(G30043,G30042,G30041);
  or GNAME30044(G30044,G34796,G29044);
  or GNAME30045(G30045,G34728,G29034);
  nand GNAME30046(G30046,G30045,G30044);
  or GNAME30047(G30047,G34802,G29041);
  or GNAME30048(G30048,G34736,G29035);
  nand GNAME30049(G30049,G30048,G30047);
  or GNAME30050(G30050,G34750,G31521);
  or GNAME30051(G30051,G34741,G29047);
  nand GNAME30052(G30052,G30051,G30050);
  or GNAME30053(G30053,G34749,G29045);
  or GNAME30054(G30054,G34740,G29046);
  nand GNAME30055(G30055,G30054,G30053);
  or GNAME30056(G30056,G34753,G31524);
  or GNAME30057(G30057,G34744,G29052);
  nand GNAME30058(G30058,G30057,G30056);
  or GNAME30059(G30059,G34751,G29050);
  or GNAME30060(G30060,G34742,G29051);
  nand GNAME30061(G30061,G30060,G30059);
  or GNAME30062(G30062,G34754,G31525);
  or GNAME30063(G30063,G34745,G29055);
  nand GNAME30064(G30064,G30063,G30062);
  or GNAME30065(G30065,G34752,G29053);
  or GNAME30066(G30066,G34743,G29054);
  nand GNAME30067(G30067,G30066,G30065);
  or GNAME30068(G30068,G34800,G29031);
  or GNAME30069(G30069,G34734,G29049);
  nand GNAME30070(G30070,G30069,G30068);
  or GNAME30071(G30071,G34794,G29030);
  or GNAME30072(G30072,G34726,G29048);
  nand GNAME30073(G30073,G30072,G30071);
  or GNAME30074(G30074,G34801,G29033);
  or GNAME30075(G30075,G34735,G29057);
  nand GNAME30076(G30076,G30075,G30074);
  or GNAME30077(G30077,G34795,G29032);
  or GNAME30078(G30078,G34727,G29056);
  nand GNAME30079(G30079,G30078,G30077);
  or GNAME30080(G30080,G34802,G29035);
  or GNAME30081(G30081,G34736,G29059);
  nand GNAME30082(G30082,G30081,G30080);
  or GNAME30083(G30083,G34796,G29034);
  or GNAME30084(G30084,G34728,G29058);
  nand GNAME30085(G30085,G30084,G30083);
  or GNAME30086(G30086,G34827,G31526);
  or GNAME30087(G30087,G34803,G29064);
  nand GNAME30088(G30088,G30087,G30086);
  or GNAME30089(G30089,G34750,G29077);
  or GNAME30090(G30090,G34741,G29078);
  nand GNAME30091(G30091,G30090,G30089);
  or GNAME30092(G30092,G34828,G31527);
  or GNAME30093(G30093,G34804,G29072);
  nand GNAME30094(G30094,G30093,G30092);
  or GNAME30095(G30095,G34753,G29081);
  or GNAME30096(G30096,G34744,G29082);
  nand GNAME30097(G30097,G30096,G30095);
  or GNAME30098(G30098,G34829,G31528);
  or GNAME30099(G30099,G34805,G29074);
  nand GNAME30100(G30100,G30099,G30098);
  or GNAME30101(G30101,G34754,G29085);
  or GNAME30102(G30102,G34745,G29086);
  nand GNAME30103(G30103,G30102,G30101);
  or GNAME30104(G30104,G34750,G29047);
  or GNAME30105(G30105,G34741,G29077);
  nand GNAME30106(G30106,G30105,G30104);
  or GNAME30107(G30107,G34753,G29052);
  or GNAME30108(G30108,G34744,G29081);
  nand GNAME30109(G30109,G30108,G30107);
  or GNAME30110(G30110,G34754,G29055);
  or GNAME30111(G30111,G34745,G29085);
  nand GNAME30112(G30112,G30111,G30110);
  or GNAME30113(G30113,G34794,G29061);
  or GNAME30114(G30114,G34726,G29076);
  nand GNAME30115(G30115,G30114,G30113);
  or GNAME30116(G30116,G34800,G29062);
  or GNAME30117(G30117,G34734,G29063);
  nand GNAME30118(G30118,G30117,G30116);
  or GNAME30119(G30119,G34749,G29060);
  or GNAME30120(G30120,G34740,G29075);
  nand GNAME30121(G30121,G30120,G30119);
  or GNAME30122(G30122,G34795,G29066);
  or GNAME30123(G30123,G34727,G29080);
  nand GNAME30124(G30124,G30123,G30122);
  or GNAME30125(G30125,G34801,G29067);
  or GNAME30126(G30126,G34735,G29071);
  nand GNAME30127(G30127,G30126,G30125);
  or GNAME30128(G30128,G34751,G29065);
  or GNAME30129(G30129,G34742,G29079);
  nand GNAME30130(G30130,G30129,G30128);
  or GNAME30131(G30131,G34796,G29069);
  or GNAME30132(G30132,G34728,G29084);
  nand GNAME30133(G30133,G30132,G30131);
  or GNAME30134(G30134,G34802,G29070);
  or GNAME30135(G30135,G34736,G29073);
  nand GNAME30136(G30136,G30135,G30134);
  or GNAME30137(G30137,G34752,G29068);
  or GNAME30138(G30138,G34743,G29083);
  nand GNAME30139(G30139,G30138,G30137);
  or GNAME30140(G30140,G34800,G29049);
  or GNAME30141(G30141,G34734,G29062);
  nand GNAME30142(G30142,G30141,G30140);
  or GNAME30143(G30143,G34794,G29048);
  or GNAME30144(G30144,G34726,G29061);
  nand GNAME30145(G30145,G30144,G30143);
  or GNAME30146(G30146,G34801,G29057);
  or GNAME30147(G30147,G34735,G29067);
  nand GNAME30148(G30148,G30147,G30146);
  or GNAME30149(G30149,G34795,G29056);
  or GNAME30150(G30150,G34727,G29066);
  nand GNAME30151(G30151,G30150,G30149);
  or GNAME30152(G30152,G34802,G29059);
  or GNAME30153(G30153,G34736,G29070);
  nand GNAME30154(G30154,G30153,G30152);
  or GNAME30155(G30155,G34796,G29058);
  or GNAME30156(G30156,G34728,G29069);
  nand GNAME30157(G30157,G30156,G30155);
  or GNAME30158(G30158,G34749,G29075);
  or GNAME30159(G30159,G34740,G29092);
  nand GNAME30160(G30160,G30159,G30158);
  or GNAME30161(G30161,G34794,G29076);
  or GNAME30162(G30162,G34726,G29091);
  nand GNAME30163(G30163,G30162,G30161);
  or GNAME30164(G30164,G34751,G29079);
  or GNAME30165(G30165,G34742,G29102);
  nand GNAME30166(G30166,G30165,G30164);
  or GNAME30167(G30167,G34795,G29080);
  or GNAME30168(G30168,G34727,G29101);
  nand GNAME30169(G30169,G30168,G30167);
  or GNAME30170(G30170,G34752,G29083);
  or GNAME30171(G30171,G34743,G29105);
  nand GNAME30172(G30172,G30171,G30170);
  or GNAME30173(G30173,G34796,G29084);
  or GNAME30174(G30174,G34728,G29104);
  nand GNAME30175(G30175,G30174,G30173);
  or GNAME30176(G30176,G34827,G29064);
  or GNAME30177(G30177,G34803,G29093);
  nand GNAME30178(G30178,G30177,G30176);
  or GNAME30179(G30179,G34800,G29063);
  or GNAME30180(G30180,G34734,G29087);
  nand GNAME30181(G30181,G30180,G30179);
  or GNAME30182(G30182,G34828,G29072);
  or GNAME30183(G30183,G34804,G29106);
  nand GNAME30184(G30184,G30183,G30182);
  or GNAME30185(G30185,G34801,G29071);
  or GNAME30186(G30186,G34735,G29088);
  nand GNAME30187(G30187,G30186,G30185);
  or GNAME30188(G30188,G34829,G29074);
  or GNAME30189(G30189,G34805,G29113);
  nand GNAME30190(G30190,G30189,G30188);
  or GNAME30191(G30191,G34802,G29073);
  or GNAME30192(G30192,G34736,G29089);
  nand GNAME30193(G30193,G30192,G30191);
  or GNAME30194(G30194,G34824,G31532);
  or GNAME30195(G30195,G34806,G29095);
  nand GNAME30196(G30196,G30195,G30194);
  or GNAME30197(G30197,G34827,G29093);
  or GNAME30198(G30198,G34803,G29094);
  nand GNAME30199(G30199,G30198,G30197);
  or GNAME30200(G30200,G34825,G31529);
  or GNAME30201(G30201,G34807,G29108);
  nand GNAME30202(G30202,G30201,G30200);
  or GNAME30203(G30203,G34828,G29106);
  or GNAME30204(G30204,G34804,G29107);
  nand GNAME30205(G30205,G30204,G30203);
  or GNAME30206(G30206,G34826,G31530);
  or GNAME30207(G30207,G34808,G29115);
  nand GNAME30208(G30208,G30207,G30206);
  or GNAME30209(G30209,G34829,G29113);
  or GNAME30210(G30210,G34805,G29114);
  nand GNAME30211(G30211,G30210,G30209);
  or GNAME30212(G30212,G34750,G29090);
  or GNAME30213(G30213,G34741,G29098);
  nand GNAME30214(G30214,G30213,G30212);
  or GNAME30215(G30215,G34794,G29091);
  or GNAME30216(G30216,G34726,G29097);
  nand GNAME30217(G30217,G30216,G30215);
  or GNAME30218(G30218,G34749,G29092);
  or GNAME30219(G30219,G34740,G29096);
  nand GNAME30220(G30220,G30219,G30218);
  or GNAME30221(G30221,G34753,G29100);
  or GNAME30222(G30222,G34744,G29111);
  nand GNAME30223(G30223,G30222,G30221);
  or GNAME30224(G30224,G34795,G29101);
  or GNAME30225(G30225,G34727,G29110);
  nand GNAME30226(G30226,G30225,G30224);
  or GNAME30227(G30227,G34751,G29102);
  or GNAME30228(G30228,G34742,G29109);
  nand GNAME30229(G30229,G30228,G30227);
  or GNAME30230(G30230,G34754,G29103);
  or GNAME30231(G30231,G34745,G29118);
  nand GNAME30232(G30232,G30231,G30230);
  or GNAME30233(G30233,G34796,G29104);
  or GNAME30234(G30234,G34728,G29117);
  nand GNAME30235(G30235,G30234,G30233);
  or GNAME30236(G30236,G34752,G29105);
  or GNAME30237(G30237,G34743,G29116);
  nand GNAME30238(G30238,G30237,G30236);
  or GNAME30239(G30239,G34749,G29096);
  or GNAME30240(G30240,G34740,G29125);
  nand GNAME30241(G30241,G30240,G30239);
  or GNAME30242(G30242,G34800,G29099);
  or GNAME30243(G30243,G34734,G29124);
  nand GNAME30244(G30244,G30243,G30242);
  or GNAME30245(G30245,G34751,G29109);
  or GNAME30246(G30246,G34742,G29138);
  nand GNAME30247(G30247,G30246,G30245);
  or GNAME30248(G30248,G34801,G29112);
  or GNAME30249(G30249,G34735,G29137);
  nand GNAME30250(G30250,G30249,G30248);
  or GNAME30251(G30251,G34752,G29116);
  or GNAME30252(G30252,G34743,G29144);
  nand GNAME30253(G30253,G30252,G30251);
  or GNAME30254(G30254,G34802,G29119);
  or GNAME30255(G30255,G34736,G29143);
  nand GNAME30256(G30256,G30255,G30254);
  or GNAME30257(G30257,G34800,G29087);
  or GNAME30258(G30258,G34734,G29099);
  nand GNAME30259(G30259,G30258,G30257);
  or GNAME30260(G30260,G34801,G29088);
  or GNAME30261(G30261,G34735,G29112);
  nand GNAME30262(G30262,G30261,G30260);
  or GNAME30263(G30263,G34802,G29089);
  or GNAME30264(G30264,G34736,G29119);
  nand GNAME30265(G30265,G30264,G30263);
  or GNAME30266(G30266,G34824,G29095);
  or GNAME30267(G30267,G34806,G29122);
  nand GNAME30268(G30268,G30267,G30266);
  or GNAME30269(G30269,G34794,G29097);
  or GNAME30270(G30270,G34788,G29121);
  nand GNAME30271(G30271,G30270,G30269);
  or GNAME30272(G30272,G34827,G29094);
  or GNAME30273(G30273,G34803,G29120);
  nand GNAME30274(G30274,G30273,G30272);
  or GNAME30275(G30275,G34827,G29120);
  or GNAME30276(G30276,G34803,G29128);
  nand GNAME30277(G30277,G30276,G30275);
  or GNAME30278(G30278,G34749,G29125);
  or GNAME30279(G30279,G34740,G29127);
  nand GNAME30280(G30280,G30279,G30278);
  or GNAME30281(G30281,G34750,G29123);
  or GNAME30282(G30282,G34741,G29126);
  nand GNAME30283(G30283,G30282,G30281);
  or GNAME30284(G30284,G34825,G29108);
  or GNAME30285(G30285,G34807,G29135);
  nand GNAME30286(G30286,G30285,G30284);
  or GNAME30287(G30287,G34795,G29110);
  or GNAME30288(G30288,G34790,G29134);
  nand GNAME30289(G30289,G30288,G30287);
  or GNAME30290(G30290,G34828,G29107);
  or GNAME30291(G30291,G34804,G29133);
  nand GNAME30292(G30292,G30291,G30290);
  or GNAME30293(G30293,G34826,G29115);
  or GNAME30294(G30294,G34808,G29141);
  nand GNAME30295(G30295,G30294,G30293);
  or GNAME30296(G30296,G34796,G29117);
  or GNAME30297(G30297,G34791,G29140);
  nand GNAME30298(G30298,G30297,G30296);
  or GNAME30299(G30299,G34829,G29114);
  or GNAME30300(G30300,G34805,G29139);
  nand GNAME30301(G30301,G30300,G30299);
  or GNAME30302(G30302,G34828,G29133);
  or GNAME30303(G30303,G34804,G29147);
  nand GNAME30304(G30304,G30303,G30302);
  or GNAME30305(G30305,G34751,G29138);
  or GNAME30306(G30306,G34742,G29146);
  nand GNAME30307(G30307,G30306,G30305);
  or GNAME30308(G30308,G34753,G29136);
  or GNAME30309(G30309,G34744,G29145);
  nand GNAME30310(G30310,G30309,G30308);
  or GNAME30311(G30311,G34829,G29139);
  or GNAME30312(G30312,G34805,G29154);
  nand GNAME30313(G30313,G30312,G30311);
  or GNAME30314(G30314,G34752,G29144);
  or GNAME30315(G30315,G34743,G29153);
  nand GNAME30316(G30316,G30315,G30314);
  or GNAME30317(G30317,G34754,G29142);
  or GNAME30318(G30318,G34745,G29152);
  nand GNAME30319(G30319,G30318,G30317);
  or GNAME30320(G30320,G34824,G29122);
  or GNAME30321(G30321,G34806,G29131);
  nand GNAME30322(G30322,G30321,G30320);
  or GNAME30323(G30323,G34731,G29121);
  or GNAME30324(G30324,G34788,G29130);
  nand GNAME30325(G30325,G30324,G30323);
  or GNAME30326(G30326,G34800,G29124);
  or GNAME30327(G30327,G34734,G29129);
  nand GNAME30328(G30328,G30327,G30326);
  or GNAME30329(G30329,G34825,G29135);
  or GNAME30330(G30330,G34807,G29150);
  nand GNAME30331(G30331,G30330,G30329);
  or GNAME30332(G30332,G34732,G29134);
  or GNAME30333(G30333,G34790,G29149);
  nand GNAME30334(G30334,G30333,G30332);
  or GNAME30335(G30335,G34801,G29137);
  or GNAME30336(G30336,G34735,G29148);
  nand GNAME30337(G30337,G30336,G30335);
  or GNAME30338(G30338,G34826,G29141);
  or GNAME30339(G30339,G34808,G29157);
  nand GNAME30340(G30340,G30339,G30338);
  or GNAME30341(G30341,G34733,G29140);
  or GNAME30342(G30342,G34791,G29156);
  nand GNAME30343(G30343,G30342,G30341);
  or GNAME30344(G30344,G34802,G29143);
  or GNAME30345(G30345,G34736,G29155);
  nand GNAME30346(G30346,G30345,G30344);
  or GNAME30347(G30347,G34750,G29126);
  or GNAME30348(G30348,G34741,G29160);
  nand GNAME30349(G30349,G30348,G30347);
  or GNAME30350(G30350,G34731,G29130);
  or GNAME30351(G30351,G34788,G29159);
  nand GNAME30352(G30352,G30351,G30350);
  or GNAME30353(G30353,G34753,G29145);
  or GNAME30354(G30354,G34744,G29174);
  nand GNAME30355(G30355,G30354,G30353);
  or GNAME30356(G30356,G34732,G29149);
  or GNAME30357(G30357,G34790,G29173);
  nand GNAME30358(G30358,G30357,G30356);
  or GNAME30359(G30359,G34754,G29152);
  or GNAME30360(G30360,G34745,G29181);
  nand GNAME30361(G30361,G30360,G30359);
  or GNAME30362(G30362,G34733,G29156);
  or GNAME30363(G30363,G34791,G29180);
  nand GNAME30364(G30364,G30363,G30362);
  or GNAME30365(G30365,G34827,G29164);
  or GNAME30366(G30366,G34803,G29168);
  nand GNAME30367(G30367,G30366,G30365);
  or GNAME30368(G30368,G34749,G29162);
  or GNAME30369(G30369,G34740,G29167);
  nand GNAME30370(G30370,G30369,G30368);
  or GNAME30371(G30371,G34750,G29160);
  or GNAME30372(G30372,G34741,G29166);
  nand GNAME30373(G30373,G30372,G30371);
  or GNAME30374(G30374,G34828,G29178);
  or GNAME30375(G30375,G34804,G29189);
  nand GNAME30376(G30376,G30375,G30374);
  or GNAME30377(G30377,G34751,G29176);
  or GNAME30378(G30378,G34742,G29188);
  nand GNAME30379(G30379,G30378,G30377);
  or GNAME30380(G30380,G34753,G29174);
  or GNAME30381(G30381,G34744,G29187);
  nand GNAME30382(G30382,G30381,G30380);
  or GNAME30383(G30383,G34829,G29185);
  or GNAME30384(G30384,G34805,G29196);
  nand GNAME30385(G30385,G30384,G30383);
  or GNAME30386(G30386,G34752,G29183);
  or GNAME30387(G30387,G34743,G29195);
  nand GNAME30388(G30388,G30387,G30386);
  or GNAME30389(G30389,G34754,G29181);
  or GNAME30390(G30390,G34745,G29194);
  nand GNAME30391(G30391,G30390,G30389);
  or GNAME30392(G30392,G34779,G29163);
  or GNAME30393(G30393,G34761,G29172);
  nand GNAME30394(G30394,G30393,G30392);
  or GNAME30395(G30395,G31535,G34764);
  or GNAME30396(G30396,G34758,G29201);
  nand GNAME30397(G30397,G30396,G30395);
  or GNAME30398(G30398,G34780,G29177);
  or GNAME30399(G30399,G34762,G29193);
  nand GNAME30400(G30400,G30399,G30398);
  or GNAME30401(G30401,G31536,G34765);
  or GNAME30402(G30402,G34759,G29202);
  nand GNAME30403(G30403,G30402,G30401);
  or GNAME30404(G30404,G34781,G29184);
  or GNAME30405(G30405,G34763,G29200);
  nand GNAME30406(G30406,G30405,G30404);
  or GNAME30407(G30407,G31537,G34766);
  or GNAME30408(G30408,G34760,G29203);
  nand GNAME30409(G30409,G30408,G30407);
  or GNAME30410(G30410,G34800,G29129);
  or GNAME30411(G30411,G34789,G29165);
  nand GNAME30412(G30412,G30411,G30410);
  or GNAME30413(G30413,G34827,G29128);
  or GNAME30414(G30414,G34803,G29164);
  nand GNAME30415(G30415,G30414,G30413);
  or GNAME30416(G30416,G34801,G29148);
  or GNAME30417(G30417,G34792,G29179);
  nand GNAME30418(G30418,G30417,G30416);
  or GNAME30419(G30419,G34828,G29147);
  or GNAME30420(G30420,G34804,G29178);
  nand GNAME30421(G30421,G30420,G30419);
  or GNAME30422(G30422,G34802,G29155);
  or GNAME30423(G30423,G34793,G29186);
  nand GNAME30424(G30424,G30423,G30422);
  or GNAME30425(G30425,G34829,G29154);
  or GNAME30426(G30426,G34805,G29185);
  nand GNAME30427(G30427,G30426,G30425);
  or GNAME30428(G30428,G34779,G29132);
  or GNAME30429(G30429,G34761,G29163);
  nand GNAME30430(G30430,G30429,G30428);
  or GNAME30431(G30431,G34749,G29127);
  or GNAME30432(G30432,G34740,G29162);
  nand GNAME30433(G30433,G30432,G30431);
  or GNAME30434(G30434,G34824,G29131);
  or GNAME30435(G30435,G34806,G29161);
  nand GNAME30436(G30436,G30435,G30434);
  or GNAME30437(G30437,G34824,G29161);
  or GNAME30438(G30438,G34806,G29171);
  nand GNAME30439(G30439,G30438,G30437);
  or GNAME30440(G30440,G34731,G29159);
  or GNAME30441(G30441,G34788,G29170);
  nand GNAME30442(G30442,G30441,G30440);
  or GNAME30443(G30443,G34737,G29165);
  or GNAME30444(G30444,G34789,G29169);
  nand GNAME30445(G30445,G30444,G30443);
  or GNAME30446(G30446,G34780,G29151);
  or GNAME30447(G30447,G34762,G29177);
  nand GNAME30448(G30448,G30447,G30446);
  or GNAME30449(G30449,G34751,G29146);
  or GNAME30450(G30450,G34742,G29176);
  nand GNAME30451(G30451,G30450,G30449);
  or GNAME30452(G30452,G34825,G29150);
  or GNAME30453(G30453,G34807,G29175);
  nand GNAME30454(G30454,G30453,G30452);
  or GNAME30455(G30455,G34781,G29158);
  or GNAME30456(G30456,G34763,G29184);
  nand GNAME30457(G30457,G30456,G30455);
  or GNAME30458(G30458,G34752,G29153);
  or GNAME30459(G30459,G34743,G29183);
  nand GNAME30460(G30460,G30459,G30458);
  or GNAME30461(G30461,G34826,G29157);
  or GNAME30462(G30462,G34808,G29182);
  nand GNAME30463(G30463,G30462,G30461);
  or GNAME30464(G30464,G34825,G29175);
  or GNAME30465(G30465,G34807,G29192);
  nand GNAME30466(G30466,G30465,G30464);
  or GNAME30467(G30467,G34732,G29173);
  or GNAME30468(G30468,G34790,G29191);
  nand GNAME30469(G30469,G30468,G30467);
  or GNAME30470(G30470,G34738,G29179);
  or GNAME30471(G30471,G34792,G29190);
  nand GNAME30472(G30472,G30471,G30470);
  or GNAME30473(G30473,G34826,G29182);
  or GNAME30474(G30474,G34808,G29199);
  nand GNAME30475(G30475,G30474,G30473);
  or GNAME30476(G30476,G34733,G29180);
  or GNAME30477(G30477,G34791,G29198);
  nand GNAME30478(G30478,G30477,G30476);
  or GNAME30479(G30479,G34739,G29186);
  or GNAME30480(G30480,G34793,G29197);
  nand GNAME30481(G30481,G30480,G30479);
  or GNAME30482(G30482,G34827,G29168);
  or GNAME30483(G30483,G34803,G29206);
  nand GNAME30484(G30484,G30483,G30482);
  or GNAME30485(G30485,G34749,G29167);
  or GNAME30486(G30486,G34797,G29205);
  nand GNAME30487(G30487,G30486,G30485);
  or GNAME30488(G30488,G34750,G29166);
  or GNAME30489(G30489,G34741,G29204);
  nand GNAME30490(G30490,G30489,G30488);
  or GNAME30491(G30491,G34827,G29206);
  or GNAME30492(G30492,G34803,G29213);
  nand GNAME30493(G30493,G30492,G30491);
  or GNAME30494(G30494,G34746,G29205);
  or GNAME30495(G30495,G34797,G29212);
  nand GNAME30496(G30496,G30495,G30494);
  or GNAME30497(G30497,G34750,G29204);
  or GNAME30498(G30498,G34741,G29211);
  nand GNAME30499(G30499,G30498,G30497);
  or GNAME30500(G30500,G34828,G29189);
  or GNAME30501(G30501,G34804,G29220);
  nand GNAME30502(G30502,G30501,G30500);
  or GNAME30503(G30503,G34751,G29188);
  or GNAME30504(G30504,G34798,G29219);
  nand GNAME30505(G30505,G30504,G30503);
  or GNAME30506(G30506,G34753,G29187);
  or GNAME30507(G30507,G34744,G29218);
  nand GNAME30508(G30508,G30507,G30506);
  or GNAME30509(G30509,G34829,G29196);
  or GNAME30510(G30510,G34805,G29227);
  nand GNAME30511(G30511,G30510,G30509);
  or GNAME30512(G30512,G34752,G29195);
  or GNAME30513(G30513,G34799,G29226);
  nand GNAME30514(G30514,G30513,G30512);
  or GNAME30515(G30515,G34754,G29194);
  or GNAME30516(G30516,G34745,G29225);
  nand GNAME30517(G30517,G30516,G30515);
  or GNAME30518(G30518,G34828,G29220);
  or GNAME30519(G30519,G34804,G29234);
  nand GNAME30520(G30520,G30519,G30518);
  or GNAME30521(G30521,G34747,G29219);
  or GNAME30522(G30522,G34798,G29233);
  nand GNAME30523(G30523,G30522,G30521);
  or GNAME30524(G30524,G34753,G29218);
  or GNAME30525(G30525,G34744,G29232);
  nand GNAME30526(G30526,G30525,G30524);
  or GNAME30527(G30527,G34829,G29227);
  or GNAME30528(G30528,G34805,G29241);
  nand GNAME30529(G30529,G30528,G30527);
  or GNAME30530(G30530,G34748,G29226);
  or GNAME30531(G30531,G34799,G29240);
  nand GNAME30532(G30532,G30531,G30530);
  or GNAME30533(G30533,G34754,G29225);
  or GNAME30534(G30534,G34745,G29239);
  nand GNAME30535(G30535,G30534,G30533);
  or GNAME30536(G30536,G34779,G29172);
  or GNAME30537(G30537,G34761,G29210);
  nand GNAME30538(G30538,G30537,G30536);
  or GNAME30539(G30539,G29201,G34764);
  or GNAME30540(G30540,G34758,G29246);
  nand GNAME30541(G30541,G30540,G30539);
  or GNAME30542(G30542,G34779,G29210);
  or GNAME30543(G30543,G34761,G29217);
  nand GNAME30544(G30544,G30543,G30542);
  or GNAME30545(G30545,G29246,G34764);
  or GNAME30546(G30546,G34758,G29247);
  nand GNAME30547(G30547,G30546,G30545);
  or GNAME30548(G30548,G34780,G29193);
  or GNAME30549(G30549,G34762,G29224);
  nand GNAME30550(G30550,G30549,G30548);
  or GNAME30551(G30551,G29202,G34765);
  or GNAME30552(G30552,G34759,G29248);
  nand GNAME30553(G30553,G30552,G30551);
  or GNAME30554(G30554,G34781,G29200);
  or GNAME30555(G30555,G34763,G29231);
  nand GNAME30556(G30556,G30555,G30554);
  or GNAME30557(G30557,G29203,G34766);
  or GNAME30558(G30558,G34760,G29249);
  nand GNAME30559(G30559,G30558,G30557);
  or GNAME30560(G30560,G34780,G29224);
  or GNAME30561(G30561,G34762,G29238);
  nand GNAME30562(G30562,G30561,G30560);
  or GNAME30563(G30563,G29248,G34765);
  or GNAME30564(G30564,G34759,G29250);
  nand GNAME30565(G30565,G30564,G30563);
  or GNAME30566(G30566,G34781,G29231);
  or GNAME30567(G30567,G34763,G29245);
  nand GNAME30568(G30568,G30567,G30566);
  or GNAME30569(G30569,G29249,G34766);
  or GNAME30570(G30570,G34760,G29251);
  nand GNAME30571(G30571,G30570,G30569);
  or GNAME30572(G30572,G34824,G29171);
  or GNAME30573(G30573,G34806,G29209);
  nand GNAME30574(G30574,G30573,G30572);
  or GNAME30575(G30575,G34731,G29170);
  or GNAME30576(G30576,G34788,G29208);
  nand GNAME30577(G30577,G30576,G30575);
  or GNAME30578(G30578,G34737,G29169);
  or GNAME30579(G30579,G34789,G29207);
  nand GNAME30580(G30580,G30579,G30578);
  or GNAME30581(G30581,G34824,G29209);
  or GNAME30582(G30582,G34806,G29216);
  nand GNAME30583(G30583,G30582,G30581);
  or GNAME30584(G30584,G34731,G29208);
  or GNAME30585(G30585,G34788,G29215);
  nand GNAME30586(G30586,G30585,G30584);
  or GNAME30587(G30587,G34737,G29207);
  or GNAME30588(G30588,G34789,G29214);
  nand GNAME30589(G30589,G30588,G30587);
  or GNAME30590(G30590,G34825,G29192);
  or GNAME30591(G30591,G34807,G29223);
  nand GNAME30592(G30592,G30591,G30590);
  or GNAME30593(G30593,G34732,G29191);
  or GNAME30594(G30594,G34790,G29222);
  nand GNAME30595(G30595,G30594,G30593);
  or GNAME30596(G30596,G34738,G29190);
  or GNAME30597(G30597,G34792,G29221);
  nand GNAME30598(G30598,G30597,G30596);
  or GNAME30599(G30599,G34826,G29199);
  or GNAME30600(G30600,G34808,G29230);
  nand GNAME30601(G30601,G30600,G30599);
  or GNAME30602(G30602,G34733,G29198);
  or GNAME30603(G30603,G34791,G29229);
  nand GNAME30604(G30604,G30603,G30602);
  or GNAME30605(G30605,G34739,G29197);
  or GNAME30606(G30606,G34793,G29228);
  nand GNAME30607(G30607,G30606,G30605);
  or GNAME30608(G30608,G34825,G29223);
  or GNAME30609(G30609,G34807,G29237);
  nand GNAME30610(G30610,G30609,G30608);
  or GNAME30611(G30611,G34732,G29222);
  or GNAME30612(G30612,G34790,G29236);
  nand GNAME30613(G30613,G30612,G30611);
  or GNAME30614(G30614,G34738,G29221);
  or GNAME30615(G30615,G34792,G29235);
  nand GNAME30616(G30616,G30615,G30614);
  or GNAME30617(G30617,G34826,G29230);
  or GNAME30618(G30618,G34808,G29244);
  nand GNAME30619(G30619,G30618,G30617);
  or GNAME30620(G30620,G34733,G29229);
  or GNAME30621(G30621,G34791,G29243);
  nand GNAME30622(G30622,G30621,G30620);
  or GNAME30623(G30623,G34739,G29228);
  or GNAME30624(G30624,G34793,G29242);
  nand GNAME30625(G30625,G30624,G30623);
  or GNAME30626(G30626,G34827,G29213);
  or GNAME30627(G30627,G34803,G29254);
  nand GNAME30628(G30628,G30627,G30626);
  or GNAME30629(G30629,G34746,G29212);
  or GNAME30630(G30630,G34797,G29253);
  nand GNAME30631(G30631,G30630,G30629);
  or GNAME30632(G30632,G34750,G29211);
  or GNAME30633(G30633,G34815,G29252);
  nand GNAME30634(G30634,G30633,G30632);
  or GNAME30635(G30635,G34827,G29254);
  or GNAME30636(G30636,G34803,G29261);
  nand GNAME30637(G30637,G30636,G30635);
  or GNAME30638(G30638,G34746,G29253);
  or GNAME30639(G30639,G34797,G29260);
  nand GNAME30640(G30640,G30639,G30638);
  or GNAME30641(G30641,G34809,G29252);
  or GNAME30642(G30642,G34815,G29259);
  nand GNAME30643(G30643,G30642,G30641);
  or GNAME30644(G30644,G34828,G29234);
  or GNAME30645(G30645,G34804,G29268);
  nand GNAME30646(G30646,G30645,G30644);
  or GNAME30647(G30647,G34747,G29233);
  or GNAME30648(G30648,G34798,G29267);
  nand GNAME30649(G30649,G30648,G30647);
  or GNAME30650(G30650,G34753,G29232);
  or GNAME30651(G30651,G34816,G29266);
  nand GNAME30652(G30652,G30651,G30650);
  or GNAME30653(G30653,G34829,G29241);
  or GNAME30654(G30654,G34805,G29275);
  nand GNAME30655(G30655,G30654,G30653);
  or GNAME30656(G30656,G34748,G29240);
  or GNAME30657(G30657,G34799,G29274);
  nand GNAME30658(G30658,G30657,G30656);
  or GNAME30659(G30659,G34754,G29239);
  or GNAME30660(G30660,G34817,G29273);
  nand GNAME30661(G30661,G30660,G30659);
  or GNAME30662(G30662,G34828,G29268);
  or GNAME30663(G30663,G34804,G29282);
  nand GNAME30664(G30664,G30663,G30662);
  or GNAME30665(G30665,G34747,G29267);
  or GNAME30666(G30666,G34798,G29281);
  nand GNAME30667(G30667,G30666,G30665);
  or GNAME30668(G30668,G34810,G29266);
  or GNAME30669(G30669,G34816,G29280);
  nand GNAME30670(G30670,G30669,G30668);
  or GNAME30671(G30671,G34829,G29275);
  or GNAME30672(G30672,G34805,G29289);
  nand GNAME30673(G30673,G30672,G30671);
  or GNAME30674(G30674,G34748,G29274);
  or GNAME30675(G30675,G34799,G29288);
  nand GNAME30676(G30676,G30675,G30674);
  or GNAME30677(G30677,G34811,G29273);
  or GNAME30678(G30678,G34817,G29287);
  nand GNAME30679(G30679,G30678,G30677);
  or GNAME30680(G30680,G34779,G29217);
  or GNAME30681(G30681,G34761,G29258);
  nand GNAME30682(G30682,G30681,G30680);
  or GNAME30683(G30683,G29247,G34764);
  or GNAME30684(G30684,G34758,G29294);
  nand GNAME30685(G30685,G30684,G30683);
  or GNAME30686(G30686,G34779,G29258);
  or GNAME30687(G30687,G34761,G29265);
  nand GNAME30688(G30688,G30687,G30686);
  or GNAME30689(G30689,G29294,G34764);
  or GNAME30690(G30690,G34758,G29295);
  nand GNAME30691(G30691,G30690,G30689);
  or GNAME30692(G30692,G34780,G29238);
  or GNAME30693(G30693,G34762,G29272);
  nand GNAME30694(G30694,G30693,G30692);
  or GNAME30695(G30695,G29250,G34765);
  or GNAME30696(G30696,G34759,G29296);
  nand GNAME30697(G30697,G30696,G30695);
  or GNAME30698(G30698,G34781,G29245);
  or GNAME30699(G30699,G34763,G29279);
  nand GNAME30700(G30700,G30699,G30698);
  or GNAME30701(G30701,G29251,G34766);
  or GNAME30702(G30702,G34760,G29297);
  nand GNAME30703(G30703,G30702,G30701);
  or GNAME30704(G30704,G34780,G29272);
  or GNAME30705(G30705,G34762,G29286);
  nand GNAME30706(G30706,G30705,G30704);
  or GNAME30707(G30707,G29296,G34765);
  or GNAME30708(G30708,G34759,G29298);
  nand GNAME30709(G30709,G30708,G30707);
  or GNAME30710(G30710,G34781,G29279);
  or GNAME30711(G30711,G34763,G29293);
  nand GNAME30712(G30712,G30711,G30710);
  or GNAME30713(G30713,G29297,G34766);
  or GNAME30714(G30714,G34760,G29299);
  nand GNAME30715(G30715,G30714,G30713);
  or GNAME30716(G30716,G34824,G29216);
  or GNAME30717(G30717,G34806,G29257);
  nand GNAME30718(G30718,G30717,G30716);
  or GNAME30719(G30719,G34731,G29215);
  or GNAME30720(G30720,G34788,G29256);
  nand GNAME30721(G30721,G30720,G30719);
  or GNAME30722(G30722,G34737,G29214);
  or GNAME30723(G30723,G34789,G29255);
  nand GNAME30724(G30724,G30723,G30722);
  or GNAME30725(G30725,G34824,G29257);
  or GNAME30726(G30726,G34806,G29264);
  nand GNAME30727(G30727,G30726,G30725);
  or GNAME30728(G30728,G34731,G29256);
  or GNAME30729(G30729,G34788,G29263);
  nand GNAME30730(G30730,G30729,G30728);
  or GNAME30731(G30731,G34737,G29255);
  or GNAME30732(G30732,G34789,G29262);
  nand GNAME30733(G30733,G30732,G30731);
  or GNAME30734(G30734,G34825,G29237);
  or GNAME30735(G30735,G34807,G29271);
  nand GNAME30736(G30736,G30735,G30734);
  or GNAME30737(G30737,G34732,G29236);
  or GNAME30738(G30738,G34790,G29270);
  nand GNAME30739(G30739,G30738,G30737);
  or GNAME30740(G30740,G34738,G29235);
  or GNAME30741(G30741,G34792,G29269);
  nand GNAME30742(G30742,G30741,G30740);
  or GNAME30743(G30743,G34826,G29244);
  or GNAME30744(G30744,G34808,G29278);
  nand GNAME30745(G30745,G30744,G30743);
  or GNAME30746(G30746,G34733,G29243);
  or GNAME30747(G30747,G34791,G29277);
  nand GNAME30748(G30748,G30747,G30746);
  or GNAME30749(G30749,G34739,G29242);
  or GNAME30750(G30750,G34793,G29276);
  nand GNAME30751(G30751,G30750,G30749);
  or GNAME30752(G30752,G34825,G29271);
  or GNAME30753(G30753,G34807,G29285);
  nand GNAME30754(G30754,G30753,G30752);
  or GNAME30755(G30755,G34732,G29270);
  or GNAME30756(G30756,G34790,G29284);
  nand GNAME30757(G30757,G30756,G30755);
  or GNAME30758(G30758,G34738,G29269);
  or GNAME30759(G30759,G34792,G29283);
  nand GNAME30760(G30760,G30759,G30758);
  or GNAME30761(G30761,G34826,G29278);
  or GNAME30762(G30762,G34808,G29292);
  nand GNAME30763(G30763,G30762,G30761);
  or GNAME30764(G30764,G34733,G29277);
  or GNAME30765(G30765,G34791,G29291);
  nand GNAME30766(G30766,G30765,G30764);
  or GNAME30767(G30767,G34739,G29276);
  or GNAME30768(G30768,G34793,G29290);
  nand GNAME30769(G30769,G30768,G30767);
  or GNAME30770(G30770,G34827,G29261);
  or GNAME30771(G30771,G34821,G29302);
  nand GNAME30772(G30772,G30771,G30770);
  or GNAME30773(G30773,G34746,G29260);
  or GNAME30774(G30774,G34797,G29301);
  nand GNAME30775(G30775,G30774,G30773);
  or GNAME30776(G30776,G34809,G29259);
  or GNAME30777(G30777,G34815,G29300);
  nand GNAME30778(G30778,G30777,G30776);
  or GNAME30779(G30779,G34812,G29302);
  or GNAME30780(G30780,G34821,G29309);
  nand GNAME30781(G30781,G30780,G30779);
  or GNAME30782(G30782,G34746,G29301);
  or GNAME30783(G30783,G34797,G29308);
  nand GNAME30784(G30784,G30783,G30782);
  or GNAME30785(G30785,G34809,G29300);
  or GNAME30786(G30786,G34815,G29307);
  nand GNAME30787(G30787,G30786,G30785);
  or GNAME30788(G30788,G34828,G29282);
  or GNAME30789(G30789,G34822,G29316);
  nand GNAME30790(G30790,G30789,G30788);
  or GNAME30791(G30791,G34747,G29281);
  or GNAME30792(G30792,G34798,G29315);
  nand GNAME30793(G30793,G30792,G30791);
  or GNAME30794(G30794,G34810,G29280);
  or GNAME30795(G30795,G34816,G29314);
  nand GNAME30796(G30796,G30795,G30794);
  or GNAME30797(G30797,G34829,G29289);
  or GNAME30798(G30798,G34823,G29323);
  nand GNAME30799(G30799,G30798,G30797);
  or GNAME30800(G30800,G34748,G29288);
  or GNAME30801(G30801,G34799,G29322);
  nand GNAME30802(G30802,G30801,G30800);
  or GNAME30803(G30803,G34811,G29287);
  or GNAME30804(G30804,G34817,G29321);
  nand GNAME30805(G30805,G30804,G30803);
  or GNAME30806(G30806,G34813,G29316);
  or GNAME30807(G30807,G34822,G29330);
  nand GNAME30808(G30808,G30807,G30806);
  or GNAME30809(G30809,G34747,G29315);
  or GNAME30810(G30810,G34798,G29329);
  nand GNAME30811(G30811,G30810,G30809);
  or GNAME30812(G30812,G34810,G29314);
  or GNAME30813(G30813,G34816,G29328);
  nand GNAME30814(G30814,G30813,G30812);
  or GNAME30815(G30815,G34814,G29323);
  or GNAME30816(G30816,G34823,G29337);
  nand GNAME30817(G30817,G30816,G30815);
  or GNAME30818(G30818,G34748,G29322);
  or GNAME30819(G30819,G34799,G29336);
  nand GNAME30820(G30820,G30819,G30818);
  or GNAME30821(G30821,G34811,G29321);
  or GNAME30822(G30822,G34817,G29335);
  nand GNAME30823(G30823,G30822,G30821);
  or GNAME30824(G30824,G34779,G29265);
  or GNAME30825(G30825,G34761,G29306);
  nand GNAME30826(G30826,G30825,G30824);
  or GNAME30827(G30827,G29295,G34764);
  or GNAME30828(G30828,G34758,G29342);
  nand GNAME30829(G30829,G30828,G30827);
  or GNAME30830(G30830,G34779,G29306);
  or GNAME30831(G30831,G34761,G29313);
  nand GNAME30832(G30832,G30831,G30830);
  or GNAME30833(G30833,G29342,G34764);
  or GNAME30834(G30834,G34758,G29343);
  nand GNAME30835(G30835,G30834,G30833);
  or GNAME30836(G30836,G34780,G29286);
  or GNAME30837(G30837,G34762,G29320);
  nand GNAME30838(G30838,G30837,G30836);
  or GNAME30839(G30839,G29298,G34765);
  or GNAME30840(G30840,G34759,G29344);
  nand GNAME30841(G30841,G30840,G30839);
  or GNAME30842(G30842,G34781,G29293);
  or GNAME30843(G30843,G34763,G29327);
  nand GNAME30844(G30844,G30843,G30842);
  or GNAME30845(G30845,G29299,G34766);
  or GNAME30846(G30846,G34760,G29345);
  nand GNAME30847(G30847,G30846,G30845);
  or GNAME30848(G30848,G34780,G29320);
  or GNAME30849(G30849,G34762,G29334);
  nand GNAME30850(G30850,G30849,G30848);
  or GNAME30851(G30851,G29344,G34765);
  or GNAME30852(G30852,G34759,G29346);
  nand GNAME30853(G30853,G30852,G30851);
  or GNAME30854(G30854,G34781,G29327);
  or GNAME30855(G30855,G34763,G29341);
  nand GNAME30856(G30856,G30855,G30854);
  or GNAME30857(G30857,G29345,G34766);
  or GNAME30858(G30858,G34760,G29347);
  nand GNAME30859(G30859,G30858,G30857);
  or GNAME30860(G30860,G34824,G29264);
  or GNAME30861(G30861,G34806,G29305);
  nand GNAME30862(G30862,G30861,G30860);
  or GNAME30863(G30863,G34731,G29263);
  or GNAME30864(G30864,G34788,G29304);
  nand GNAME30865(G30865,G30864,G30863);
  or GNAME30866(G30866,G34737,G29262);
  or GNAME30867(G30867,G34789,G29303);
  nand GNAME30868(G30868,G30867,G30866);
  or GNAME30869(G30869,G34824,G29305);
  or GNAME30870(G30870,G34806,G29312);
  nand GNAME30871(G30871,G30870,G30869);
  or GNAME30872(G30872,G34731,G29304);
  or GNAME30873(G30873,G34788,G29311);
  nand GNAME30874(G30874,G30873,G30872);
  or GNAME30875(G30875,G34737,G29303);
  or GNAME30876(G30876,G34789,G29310);
  nand GNAME30877(G30877,G30876,G30875);
  or GNAME30878(G30878,G34825,G29285);
  or GNAME30879(G30879,G34807,G29319);
  nand GNAME30880(G30880,G30879,G30878);
  or GNAME30881(G30881,G34732,G29284);
  or GNAME30882(G30882,G34790,G29318);
  nand GNAME30883(G30883,G30882,G30881);
  or GNAME30884(G30884,G34738,G29283);
  or GNAME30885(G30885,G34792,G29317);
  nand GNAME30886(G30886,G30885,G30884);
  or GNAME30887(G30887,G34826,G29292);
  or GNAME30888(G30888,G34808,G29326);
  nand GNAME30889(G30889,G30888,G30887);
  or GNAME30890(G30890,G34733,G29291);
  or GNAME30891(G30891,G34791,G29325);
  nand GNAME30892(G30892,G30891,G30890);
  or GNAME30893(G30893,G34739,G29290);
  or GNAME30894(G30894,G34793,G29324);
  nand GNAME30895(G30895,G30894,G30893);
  or GNAME30896(G30896,G34825,G29319);
  or GNAME30897(G30897,G34807,G29333);
  nand GNAME30898(G30898,G30897,G30896);
  or GNAME30899(G30899,G34732,G29318);
  or GNAME30900(G30900,G34790,G29332);
  nand GNAME30901(G30901,G30900,G30899);
  or GNAME30902(G30902,G34738,G29317);
  or GNAME30903(G30903,G34792,G29331);
  nand GNAME30904(G30904,G30903,G30902);
  or GNAME30905(G30905,G34826,G29326);
  or GNAME30906(G30906,G34808,G29340);
  nand GNAME30907(G30907,G30906,G30905);
  or GNAME30908(G30908,G34733,G29325);
  or GNAME30909(G30909,G34791,G29339);
  nand GNAME30910(G30910,G30909,G30908);
  or GNAME30911(G30911,G34739,G29324);
  or GNAME30912(G30912,G34793,G29338);
  nand GNAME30913(G30913,G30912,G30911);
  or GNAME30914(G30914,G34812,G29309);
  or GNAME30915(G30915,G34821,G29353);
  nand GNAME30916(G30916,G30915,G30914);
  or GNAME30917(G30917,G34746,G29308);
  or GNAME30918(G30918,G34797,G29352);
  nand GNAME30919(G30919,G30918,G30917);
  or GNAME30920(G30920,G34809,G29307);
  or GNAME30921(G30921,G34815,G29351);
  nand GNAME30922(G30922,G30921,G30920);
  or GNAME30923(G30923,G34812,G29353);
  or GNAME30924(G30924,G34821,G29360);
  nand GNAME30925(G30925,G30924,G30923);
  or GNAME30926(G30926,G34746,G29352);
  or GNAME30927(G30927,G34797,G29359);
  nand GNAME30928(G30928,G30927,G30926);
  or GNAME30929(G30929,G34809,G29351);
  or GNAME30930(G30930,G34815,G29358);
  nand GNAME30931(G30931,G30930,G30929);
  or GNAME30932(G30932,G34813,G29330);
  or GNAME30933(G30933,G34822,G29365);
  nand GNAME30934(G30934,G30933,G30932);
  or GNAME30935(G30935,G34747,G29329);
  or GNAME30936(G30936,G34798,G29364);
  nand GNAME30937(G30937,G30936,G30935);
  or GNAME30938(G30938,G34810,G29328);
  or GNAME30939(G30939,G34816,G29363);
  nand GNAME30940(G30940,G30939,G30938);
  or GNAME30941(G30941,G34814,G29337);
  or GNAME30942(G30942,G34823,G29372);
  nand GNAME30943(G30943,G30942,G30941);
  or GNAME30944(G30944,G34748,G29336);
  or GNAME30945(G30945,G34799,G29371);
  nand GNAME30946(G30946,G30945,G30944);
  or GNAME30947(G30947,G34811,G29335);
  or GNAME30948(G30948,G34817,G29370);
  nand GNAME30949(G30949,G30948,G30947);
  or GNAME30950(G30950,G34813,G29365);
  or GNAME30951(G30951,G34822,G29379);
  nand GNAME30952(G30952,G30951,G30950);
  or GNAME30953(G30953,G34747,G29364);
  or GNAME30954(G30954,G34798,G29378);
  nand GNAME30955(G30955,G30954,G30953);
  or GNAME30956(G30956,G34810,G29363);
  or GNAME30957(G30957,G34816,G29377);
  nand GNAME30958(G30958,G30957,G30956);
  or GNAME30959(G30959,G34814,G29372);
  or GNAME30960(G30960,G34823,G29384);
  nand GNAME30961(G30961,G30960,G30959);
  or GNAME30962(G30962,G34748,G29371);
  or GNAME30963(G30963,G34799,G29383);
  nand GNAME30964(G30964,G30963,G30962);
  or GNAME30965(G30965,G34811,G29370);
  or GNAME30966(G30966,G34817,G29382);
  nand GNAME30967(G30967,G30966,G30965);
  or GNAME30968(G30968,G34779,G29313);
  or GNAME30969(G30969,G34761,G29357);
  nand GNAME30970(G30970,G30969,G30968);
  or GNAME30971(G30971,G29343,G34764);
  or GNAME30972(G30972,G34758,G29387);
  nand GNAME30973(G30973,G30972,G30971);
  or GNAME30974(G30974,G34780,G29334);
  or GNAME30975(G30975,G34762,G29369);
  nand GNAME30976(G30976,G30975,G30974);
  or GNAME30977(G30977,G29346,G34765);
  or GNAME30978(G30978,G34759,G29388);
  nand GNAME30979(G30979,G30978,G30977);
  or GNAME30980(G30980,G34781,G29341);
  or GNAME30981(G30981,G34763,G29376);
  nand GNAME30982(G30982,G30981,G30980);
  or GNAME30983(G30983,G29347,G34766);
  or GNAME30984(G30984,G34760,G29389);
  nand GNAME30985(G30985,G30984,G30983);
  or GNAME30986(G30986,G34824,G29312);
  or GNAME30987(G30987,G34818,G29356);
  nand GNAME30988(G30988,G30987,G30986);
  or GNAME30989(G30989,G34731,G29311);
  or GNAME30990(G30990,G34788,G29355);
  nand GNAME30991(G30991,G30990,G30989);
  or GNAME30992(G30992,G34737,G29310);
  or GNAME30993(G30993,G34789,G29354);
  nand GNAME30994(G30994,G30993,G30992);
  or GNAME30995(G30995,G34773,G29356);
  or GNAME30996(G30996,G34818,G29348);
  nand GNAME30997(G30997,G30996,G30995);
  or GNAME30998(G30998,G34731,G29355);
  or GNAME30999(G30999,G34788,G29399);
  nand GNAME31000(G31000,G30999,G30998);
  or GNAME31001(G31001,G34737,G29354);
  or GNAME31002(G31002,G34789,G29361);
  nand GNAME31003(G31003,G31002,G31001);
  or GNAME31004(G31004,G34825,G29333);
  or GNAME31005(G31005,G34819,G29368);
  nand GNAME31006(G31006,G31005,G31004);
  or GNAME31007(G31007,G34732,G29332);
  or GNAME31008(G31008,G34790,G29367);
  nand GNAME31009(G31009,G31008,G31007);
  or GNAME31010(G31010,G34738,G29331);
  or GNAME31011(G31011,G34792,G29366);
  nand GNAME31012(G31012,G31011,G31010);
  or GNAME31013(G31013,G34826,G29340);
  or GNAME31014(G31014,G34820,G29375);
  nand GNAME31015(G31015,G31014,G31013);
  or GNAME31016(G31016,G34733,G29339);
  or GNAME31017(G31017,G34791,G29374);
  nand GNAME31018(G31018,G31017,G31016);
  or GNAME31019(G31019,G34739,G29338);
  or GNAME31020(G31020,G34793,G29373);
  nand GNAME31021(G31021,G31020,G31019);
  or GNAME31022(G31022,G34775,G29368);
  or GNAME31023(G31023,G34819,G29349);
  nand GNAME31024(G31024,G31023,G31022);
  or GNAME31025(G31025,G34732,G29367);
  or GNAME31026(G31026,G34790,G29412);
  nand GNAME31027(G31027,G31026,G31025);
  or GNAME31028(G31028,G34738,G29366);
  or GNAME31029(G31029,G34792,G29380);
  nand GNAME31030(G31030,G31029,G31028);
  or GNAME31031(G31031,G34777,G29375);
  or GNAME31032(G31032,G34820,G29350);
  nand GNAME31033(G31033,G31032,G31031);
  or GNAME31034(G31034,G34733,G29374);
  or GNAME31035(G31035,G34791,G29418);
  nand GNAME31036(G31036,G31035,G31034);
  or GNAME31037(G31037,G34739,G29373);
  or GNAME31038(G31038,G34793,G29385);
  nand GNAME31039(G31039,G31038,G31037);
  or GNAME31040(G31040,G34746,G29359);
  or GNAME31041(G31041,G34797,G29402);
  nand GNAME31042(G31042,G31041,G31040);
  or GNAME31043(G31043,G34779,G29362);
  or GNAME31044(G31044,G34770,G29401);
  nand GNAME31045(G31045,G31044,G31043);
  or GNAME31046(G31046,G34812,G29360);
  or GNAME31047(G31047,G34821,G29400);
  nand GNAME31048(G31048,G31047,G31046);
  or GNAME31049(G31049,G34747,G29378);
  or GNAME31050(G31050,G34798,G29415);
  nand GNAME31051(G31051,G31050,G31049);
  or GNAME31052(G31052,G34780,G29381);
  or GNAME31053(G31053,G34771,G29414);
  nand GNAME31054(G31054,G31053,G31052);
  or GNAME31055(G31055,G34813,G29379);
  or GNAME31056(G31056,G34822,G29413);
  nand GNAME31057(G31057,G31056,G31055);
  or GNAME31058(G31058,G34748,G29383);
  or GNAME31059(G31059,G34799,G29421);
  nand GNAME31060(G31060,G31059,G31058);
  or GNAME31061(G31061,G34781,G29386);
  or GNAME31062(G31062,G34772,G29420);
  nand GNAME31063(G31063,G31062,G31061);
  or GNAME31064(G31064,G34814,G29384);
  or GNAME31065(G31065,G34823,G29419);
  nand GNAME31066(G31066,G31065,G31064);
  or GNAME31067(G31067,G34812,G29400);
  or GNAME31068(G31068,G34821,G29411);
  nand GNAME31069(G31069,G31068,G31067);
  or GNAME31070(G31070,G34809,G29404);
  or GNAME31071(G31071,G34815,G29410);
  nand GNAME31072(G31072,G31071,G31070);
  or GNAME31073(G31073,G34813,G29413);
  or GNAME31074(G31074,G34822,G29430);
  nand GNAME31075(G31075,G31074,G31073);
  or GNAME31076(G31076,G34810,G29417);
  or GNAME31077(G31077,G34816,G29429);
  nand GNAME31078(G31078,G31077,G31076);
  or GNAME31079(G31079,G34814,G29419);
  or GNAME31080(G31080,G34823,G29437);
  nand GNAME31081(G31081,G31080,G31079);
  or GNAME31082(G31082,G34811,G29423);
  or GNAME31083(G31083,G34817,G29436);
  nand GNAME31084(G31084,G31083,G31082);
  or GNAME31085(G31085,G34773,G29348);
  or GNAME31086(G31086,G34818,G29408);
  nand GNAME31087(G31087,G31086,G31085);
  or GNAME31088(G31088,G34775,G29349);
  or GNAME31089(G31089,G34819,G29427);
  nand GNAME31090(G31090,G31089,G31088);
  or GNAME31091(G31091,G34777,G29350);
  or GNAME31092(G31092,G34820,G29434);
  nand GNAME31093(G31093,G31092,G31091);
  or GNAME31094(G31094,G34809,G29358);
  or GNAME31095(G31095,G34815,G29404);
  nand GNAME31096(G31096,G31095,G31094);
  or GNAME31097(G31097,G34737,G29361);
  or GNAME31098(G31098,G34789,G29403);
  nand GNAME31099(G31099,G31098,G31097);
  or GNAME31100(G31100,G34794,G27861);
  or GNAME31101(G31101,G34726,G31513);
  nand GNAME31102(G31102,G31101,G31100);
  or GNAME31103(G31103,G34773,G29408);
  or GNAME31104(G31104,G34818,G29409);
  nand GNAME31105(G31105,G31104,G31103);
  or GNAME31106(G31106,G34737,G29403);
  or GNAME31107(G31107,G34789,G29407);
  nand GNAME31108(G31108,G31107,G31106);
  or GNAME31109(G31109,G34746,G29402);
  or GNAME31110(G31110,G34797,G29406);
  nand GNAME31111(G31111,G31110,G31109);
  or GNAME31112(G31112,G34810,G29377);
  or GNAME31113(G31113,G34816,G29417);
  nand GNAME31114(G31114,G31113,G31112);
  or GNAME31115(G31115,G34738,G29380);
  or GNAME31116(G31116,G34792,G29416);
  nand GNAME31117(G31117,G31116,G31115);
  or GNAME31118(G31118,G34795,G27864);
  or GNAME31119(G31119,G34727,G31512);
  nand GNAME31120(G31120,G31119,G31118);
  or GNAME31121(G31121,G34811,G29382);
  or GNAME31122(G31122,G34817,G29423);
  nand GNAME31123(G31123,G31122,G31121);
  or GNAME31124(G31124,G34739,G29385);
  or GNAME31125(G31125,G34793,G29422);
  nand GNAME31126(G31126,G31125,G31124);
  or GNAME31127(G31127,G34796,G27867);
  or GNAME31128(G31128,G34728,G31514);
  nand GNAME31129(G31129,G31128,G31127);
  or GNAME31130(G31130,G34775,G29427);
  or GNAME31131(G31131,G34819,G29428);
  nand GNAME31132(G31132,G31131,G31130);
  or GNAME31133(G31133,G34738,G29416);
  or GNAME31134(G31134,G34792,G29426);
  nand GNAME31135(G31135,G31134,G31133);
  or GNAME31136(G31136,G34747,G29415);
  or GNAME31137(G31137,G34798,G29425);
  nand GNAME31138(G31138,G31137,G31136);
  or GNAME31139(G31139,G34777,G29434);
  or GNAME31140(G31140,G34820,G29435);
  nand GNAME31141(G31141,G31140,G31139);
  or GNAME31142(G31142,G34739,G29422);
  or GNAME31143(G31143,G34793,G29433);
  nand GNAME31144(G31144,G31143,G31142);
  or GNAME31145(G31145,G34748,G29421);
  or GNAME31146(G31146,G34799,G29432);
  nand GNAME31147(G31147,G31146,G31145);
  or GNAME31148(G31148,G34809,G29410);
  or GNAME31149(G31149,G34815,G29465);
  nand GNAME31150(G31150,G31149,G31148);
  or GNAME31151(G31151,G34774,G29405);
  or GNAME31152(G31152,G34770,G29464);
  nand GNAME31153(G31153,G31152,G31151);
  or GNAME31154(G31154,G34773,G29409);
  or GNAME31155(G31155,G34818,G29463);
  nand GNAME31156(G31156,G31155,G31154);
  or GNAME31157(G31157,G34773,G29463);
  or GNAME31158(G31158,G34818,G29449);
  nand GNAME31159(G31159,G31158,G31157);
  or GNAME31160(G31160,G34746,G29462);
  or GNAME31161(G31161,G34797,G29466);
  nand GNAME31162(G31162,G31161,G31160);
  or GNAME31163(G31163,G34809,G29465);
  or GNAME31164(G31164,G34815,G29447);
  nand GNAME31165(G31165,G31164,G31163);
  or GNAME31166(G31166,G34810,G29429);
  or GNAME31167(G31167,G34816,G29472);
  nand GNAME31168(G31168,G31167,G31166);
  or GNAME31169(G31169,G34776,G29424);
  or GNAME31170(G31170,G34771,G29471);
  nand GNAME31171(G31171,G31170,G31169);
  or GNAME31172(G31172,G34775,G29428);
  or GNAME31173(G31173,G34819,G29470);
  nand GNAME31174(G31174,G31173,G31172);
  or GNAME31175(G31175,G34811,G29436);
  or GNAME31176(G31176,G34817,G29476);
  nand GNAME31177(G31177,G31176,G31175);
  or GNAME31178(G31178,G34778,G29431);
  or GNAME31179(G31179,G34772,G29475);
  nand GNAME31180(G31180,G31179,G31178);
  or GNAME31181(G31181,G34777,G29435);
  or GNAME31182(G31182,G34820,G29474);
  nand GNAME31183(G31183,G31182,G31181);
  or GNAME31184(G31184,G34775,G29470);
  or GNAME31185(G31185,G34819,G29454);
  nand GNAME31186(G31186,G31185,G31184);
  or GNAME31187(G31187,G34747,G29469);
  or GNAME31188(G31188,G34798,G29477);
  nand GNAME31189(G31189,G31188,G31187);
  or GNAME31190(G31190,G34810,G29472);
  or GNAME31191(G31191,G34816,G29452);
  nand GNAME31192(G31192,G31191,G31190);
  or GNAME31193(G31193,G34777,G29474);
  or GNAME31194(G31194,G34820,G29459);
  nand GNAME31195(G31195,G31194,G31193);
  or GNAME31196(G31196,G34748,G29473);
  or GNAME31197(G31197,G34799,G29480);
  nand GNAME31198(G31198,G31197,G31196);
  or GNAME31199(G31199,G34811,G29476);
  or GNAME31200(G31200,G34817,G29457);
  nand GNAME31201(G31201,G31200,G31199);
  or GNAME31202(G31202,G34812,G29396);
  or GNAME31203(G31203,G34821,G29468);
  nand GNAME31204(G31204,G31203,G31202);
  or GNAME31205(G31205,G34773,G29449);
  or GNAME31206(G31206,G34818,G29450);
  nand GNAME31207(G31207,G31206,G31205);
  or GNAME31208(G31208,G34809,G29447);
  or GNAME31209(G31209,G34815,G29448);
  nand GNAME31210(G31210,G31209,G31208);
  or GNAME31211(G31211,G34813,G29397);
  or GNAME31212(G31212,G34822,G29479);
  nand GNAME31213(G31213,G31212,G31211);
  or GNAME31214(G31214,G34814,G29398);
  or GNAME31215(G31215,G34823,G29482);
  nand GNAME31216(G31216,G31215,G31214);
  or GNAME31217(G31217,G34775,G29454);
  or GNAME31218(G31218,G34819,G29455);
  nand GNAME31219(G31219,G31218,G31217);
  or GNAME31220(G31220,G34810,G29452);
  or GNAME31221(G31221,G34816,G29453);
  nand GNAME31222(G31222,G31221,G31220);
  or GNAME31223(G31223,G34777,G29459);
  or GNAME31224(G31224,G34820,G29460);
  nand GNAME31225(G31225,G31224,G31223);
  or GNAME31226(G31226,G34811,G29457);
  or GNAME31227(G31227,G34817,G29458);
  nand GNAME31228(G31228,G31227,G31226);
  or GNAME31229(G31229,G34812,G29411);
  or GNAME31230(G31230,G34821,G29396);
  nand GNAME31231(G31231,G31230,G31229);
  or GNAME31232(G31232,G34746,G29406);
  or GNAME31233(G31233,G34797,G29462);
  nand GNAME31234(G31234,G31233,G31232);
  or GNAME31235(G31235,G34800,G27870);
  or GNAME31236(G31236,G34734,G31515);
  nand GNAME31237(G31237,G31236,G31235);
  or GNAME31238(G31238,G34813,G29430);
  or GNAME31239(G31239,G34822,G29397);
  nand GNAME31240(G31240,G31239,G31238);
  or GNAME31241(G31241,G34747,G29425);
  or GNAME31242(G31242,G34798,G29469);
  nand GNAME31243(G31243,G31242,G31241);
  or GNAME31244(G31244,G34801,G27873);
  or GNAME31245(G31245,G34735,G31516);
  nand GNAME31246(G31246,G31245,G31244);
  or GNAME31247(G31247,G34814,G29437);
  or GNAME31248(G31248,G34823,G29398);
  nand GNAME31249(G31249,G31248,G31247);
  or GNAME31250(G31250,G34748,G29432);
  or GNAME31251(G31251,G34799,G29473);
  nand GNAME31252(G31252,G31251,G31250);
  or GNAME31253(G31253,G34802,G27876);
  or GNAME31254(G31254,G34736,G31517);
  nand GNAME31255(G31255,G31254,G31253);
  or GNAME31256(G31256,G34812,G29468);
  or GNAME31257(G31257,G34821,G29451);
  nand GNAME31258(G31258,G31257,G31256);
  or GNAME31259(G31259,G34774,G29467);
  or GNAME31260(G31260,G34770,G29507);
  nand GNAME31261(G31261,G31260,G31259);
  or GNAME31262(G31262,G34749,G27879);
  or GNAME31263(G31263,G34740,G31520);
  nand GNAME31264(G31264,G31263,G31262);
  or GNAME31265(G31265,G34813,G29479);
  or GNAME31266(G31266,G34822,G29456);
  nand GNAME31267(G31267,G31266,G31265);
  or GNAME31268(G31268,G34776,G29478);
  or GNAME31269(G31269,G34771,G29513);
  nand GNAME31270(G31270,G31269,G31268);
  or GNAME31271(G31271,G34751,G27882);
  or GNAME31272(G31272,G34742,G31522);
  nand GNAME31273(G31273,G31272,G31271);
  or GNAME31274(G31274,G34814,G29482);
  or GNAME31275(G31275,G34823,G29461);
  nand GNAME31276(G31276,G31275,G31274);
  or GNAME31277(G31277,G34778,G29481);
  or GNAME31278(G31278,G34772,G29517);
  nand GNAME31279(G31279,G31278,G31277);
  or GNAME31280(G31280,G34752,G27885);
  or GNAME31281(G31281,G34743,G31523);
  nand GNAME31282(G31282,G31281,G31280);
  or GNAME31283(G31283,G34812,G29504);
  or GNAME31284(G31284,G34821,G29496);
  nand GNAME31285(G31285,G31284,G31283);
  or GNAME31286(G31286,G34773,G29506);
  or GNAME31287(G31287,G34818,G29497);
  nand GNAME31288(G31288,G31287,G31286);
  or GNAME31289(G31289,G34750,G27888);
  or GNAME31290(G31290,G34741,G31521);
  nand GNAME31291(G31291,G31290,G31289);
  or GNAME31292(G31292,G34813,G29510);
  or GNAME31293(G31293,G34822,G29500);
  nand GNAME31294(G31294,G31293,G31292);
  or GNAME31295(G31295,G34775,G29512);
  or GNAME31296(G31296,G34819,G29501);
  nand GNAME31297(G31297,G31296,G31295);
  or GNAME31298(G31298,G34753,G27891);
  or GNAME31299(G31299,G34744,G31524);
  nand GNAME31300(G31300,G31299,G31298);
  or GNAME31301(G31301,G34814,G29514);
  or GNAME31302(G31302,G34823,G29502);
  nand GNAME31303(G31303,G31302,G31301);
  or GNAME31304(G31304,G34777,G29516);
  or GNAME31305(G31305,G34820,G29503);
  nand GNAME31306(G31306,G31305,G31304);
  or GNAME31307(G31307,G34754,G27894);
  or GNAME31308(G31308,G34745,G31525);
  nand GNAME31309(G31309,G31308,G31307);
  or GNAME31310(G31310,G34773,G29450);
  or GNAME31311(G31311,G34818,G29506);
  nand GNAME31312(G31312,G31311,G31310);
  or GNAME31313(G31313,G34809,G29448);
  or GNAME31314(G31314,G34815,G29505);
  nand GNAME31315(G31315,G31314,G31313);
  or GNAME31316(G31316,G34812,G29451);
  or GNAME31317(G31317,G34821,G29504);
  nand GNAME31318(G31318,G31317,G31316);
  or GNAME31319(G31319,G34775,G29455);
  or GNAME31320(G31320,G34819,G29512);
  nand GNAME31321(G31321,G31320,G31319);
  or GNAME31322(G31322,G34810,G29453);
  or GNAME31323(G31323,G34816,G29511);
  nand GNAME31324(G31324,G31323,G31322);
  or GNAME31325(G31325,G34813,G29456);
  or GNAME31326(G31326,G34822,G29510);
  nand GNAME31327(G31327,G31326,G31325);
  or GNAME31328(G31328,G34777,G29460);
  or GNAME31329(G31329,G34820,G29516);
  nand GNAME31330(G31330,G31329,G31328);
  or GNAME31331(G31331,G34811,G29458);
  or GNAME31332(G31332,G34817,G29515);
  nand GNAME31333(G31333,G31332,G31331);
  or GNAME31334(G31334,G34814,G29461);
  or GNAME31335(G31335,G34823,G29514);
  nand GNAME31336(G31336,G31335,G31334);
  or GNAME31337(G31337,G34774,G29542);
  or GNAME31338(G31338,G34770,G29543);
  nand GNAME31339(G31339,G31338,G31337);
  or GNAME31340(G31340,G34773,G29541);
  or GNAME31341(G31341,G34818,G29540);
  nand GNAME31342(G31342,G31341,G31340);
  or GNAME31343(G31343,G34827,G27897);
  or GNAME31344(G31344,G34803,G31526);
  nand GNAME31345(G31345,G31344,G31343);
  or GNAME31346(G31346,G34776,G29546);
  or GNAME31347(G31347,G34771,G29547);
  nand GNAME31348(G31348,G31347,G31346);
  or GNAME31349(G31349,G34775,G29544);
  or GNAME31350(G31350,G34819,G29545);
  nand GNAME31351(G31351,G31350,G31349);
  or GNAME31352(G31352,G34828,G27900);
  or GNAME31353(G31353,G34804,G31527);
  nand GNAME31354(G31354,G31353,G31352);
  or GNAME31355(G31355,G34778,G29550);
  or GNAME31356(G31356,G34772,G29551);
  nand GNAME31357(G31357,G31356,G31355);
  or GNAME31358(G31358,G34777,G29548);
  or GNAME31359(G31359,G34820,G29549);
  nand GNAME31360(G31360,G31359,G31358);
  or GNAME31361(G31361,G34829,G27903);
  or GNAME31362(G31362,G34805,G31528);
  nand GNAME31363(G31363,G31362,G31361);
  or GNAME31364(G31364,G34773,G29497);
  or GNAME31365(G31365,G34818,G29541);
  nand GNAME31366(G31366,G31365,G31364);
  or GNAME31367(G31367,G34812,G29496);
  or GNAME31368(G31368,G34821,G29509);
  nand GNAME31369(G31369,G31368,G31367);
  or GNAME31370(G31370,G34775,G29501);
  or GNAME31371(G31371,G34819,G29544);
  nand GNAME31372(G31372,G31371,G31370);
  or GNAME31373(G31373,G34813,G29500);
  or GNAME31374(G31374,G34822,G29520);
  nand GNAME31375(G31375,G31374,G31373);
  or GNAME31376(G31376,G34777,G29503);
  or GNAME31377(G31377,G34820,G29548);
  nand GNAME31378(G31378,G31377,G31376);
  or GNAME31379(G31379,G34814,G29502);
  or GNAME31380(G31380,G34823,G29521);
  nand GNAME31381(G31381,G31380,G31379);
  or GNAME31382(G31382,G34774,G29495);
  or GNAME31383(G31383,G34770,G29508);
  nand GNAME31384(G31384,G31383,G31382);
  or GNAME31385(G31385,G34776,G29498);
  or GNAME31386(G31386,G34771,G29518);
  nand GNAME31387(G31387,G31386,G31385);
  or GNAME31388(G31388,G34778,G29499);
  or GNAME31389(G31389,G34772,G29519);
  nand GNAME31390(G31390,G31389,G31388);
  or GNAME31391(G31391,G34773,G29540);
  or GNAME31392(G31392,G34818,G29553);
  nand GNAME31393(G31393,G31392,G31391);
  or GNAME31394(G31394,G34775,G29545);
  or GNAME31395(G31395,G34819,G29555);
  nand GNAME31396(G31396,G31395,G31394);
  or GNAME31397(G31397,G34777,G29549);
  or GNAME31398(G31398,G34820,G29557);
  nand GNAME31399(G31399,G31398,G31397);
  or GNAME31400(G31400,G34779,G27906);
  or GNAME31401(G31401,G34761,G31531);
  nand GNAME31402(G31402,G31401,G31400);
  or GNAME31403(G31403,G34780,G27909);
  or GNAME31404(G31404,G34762,G31533);
  nand GNAME31405(G31405,G31404,G31403);
  or GNAME31406(G31406,G34781,G27912);
  or GNAME31407(G31407,G34763,G31534);
  nand GNAME31408(G31408,G31407,G31406);
  or GNAME31409(G31409,G34774,G29552);
  or GNAME31410(G31410,G34770,G29564);
  nand GNAME31411(G31411,G31410,G31409);
  or GNAME31412(G31412,G29558,G34755);
  or GNAME31413(G31413,G34767,G29570);
  nand GNAME31414(G31414,G31413,G31412);
  or GNAME31415(G31415,G34776,G29554);
  or GNAME31416(G31416,G34771,G29566);
  nand GNAME31417(G31417,G31416,G31415);
  or GNAME31418(G31418,G29562,G34756);
  or GNAME31419(G31419,G34768,G29572);
  nand GNAME31420(G31420,G31419,G31418);
  or GNAME31421(G31421,G34778,G29556);
  or GNAME31422(G31422,G34772,G29568);
  nand GNAME31423(G31423,G31422,G31421);
  or GNAME31424(G31424,G29563,G34757);
  or GNAME31425(G31425,G34769,G29574);
  nand GNAME31426(G31426,G31425,G31424);
  or GNAME31427(G31427,G29571,G34755);
  or GNAME31428(G31428,G34767,G29576);
  nand GNAME31429(G31429,G31428,G31427);
  or GNAME31430(G31430,G29573,G34756);
  or GNAME31431(G31431,G34768,G29578);
  nand GNAME31432(G31432,G31431,G31430);
  or GNAME31433(G31433,G29575,G34757);
  or GNAME31434(G31434,G34769,G29580);
  nand GNAME31435(G31435,G31434,G31433);
  not GNAME31436(G31436,G32863);
  not GNAME31437(G31437,G31628);
  not GNAME31438(G31438,G31641);
  not GNAME31439(G31439,G2344);
  not GNAME31440(G31440,G1928);
  not GNAME31441(G31441,G1512);
  not GNAME31442(G31442,G34597);
  not GNAME31443(G31443,G34602);
  not GNAME31444(G31444,G34601);
  not GNAME31445(G31445,G34603);
  not GNAME31446(G31446,G34611);
  not GNAME31447(G31447,G34610);
  not GNAME31448(G31448,G34612);
  not GNAME31449(G31449,G34607);
  not GNAME31450(G31450,G34608);
  not GNAME31451(G31451,G34609);
  not GNAME31452(G31452,G34619);
  not GNAME31453(G31453,G34620);
  not GNAME31454(G31454,G34621);
  not GNAME31455(G31455,G34616);
  not GNAME31456(G31456,G34617);
  not GNAME31457(G31457,G34618);
  not GNAME31458(G31458,G34628);
  not GNAME31459(G31459,G34629);
  not GNAME31460(G31460,G34630);
  not GNAME31461(G31461,G34625);
  not GNAME31462(G31462,G34626);
  not GNAME31463(G31463,G34627);
  not GNAME31464(G31464,G34637);
  not GNAME31465(G31465,G34638);
  not GNAME31466(G31466,G34639);
  not GNAME31467(G31467,G34634);
  not GNAME31468(G31468,G34635);
  not GNAME31469(G31469,G34636);
  not GNAME31470(G31470,G34644);
  not GNAME31471(G31471,G34646);
  not GNAME31472(G31472,G34648);
  not GNAME31473(G31473,G34643);
  not GNAME31474(G31474,G34645);
  not GNAME31475(G31475,G34647);
  not GNAME31476(G31476,G34662);
  not GNAME31477(G31477,G34665);
  not GNAME31478(G31478,G34667);
  not GNAME31479(G31479,G34681);
  not GNAME31480(G31480,G34683);
  not GNAME31481(G31481,G34685);
  not GNAME31482(G31482,G34663);
  not GNAME31483(G31483,G34666);
  not GNAME31484(G31484,G34668);
  not GNAME31485(G31485,G34664);
  not GNAME31486(G31486,G34669);
  not GNAME31487(G31487,G34670);
  not GNAME31488(G31488,G34686);
  not GNAME31489(G31489,G34687);
  not GNAME31490(G31490,G34688);
  not GNAME31491(G31491,G34680);
  not GNAME31492(G31492,G34695);
  not GNAME31493(G31493,G34682);
  not GNAME31494(G31494,G34684);
  not GNAME31495(G31495,G34696);
  not GNAME31496(G31496,G34697);
  not GNAME31497(G31497,G34692);
  not GNAME31498(G31498,G34693);
  not GNAME31499(G31499,G34700);
  not GNAME31500(G31500,G34703);
  not GNAME31501(G31501,G34699);
  not GNAME31502(G31502,G34702);
  not GNAME31503(G31503,G34694);
  not GNAME31504(G31504,G34713);
  not GNAME31505(G31505,G34698);
  not GNAME31506(G31506,G34701);
  not GNAME31507(G31507,G34715);
  not GNAME31508(G31508,G34717);
  not GNAME31509(G31509,G34714);
  not GNAME31510(G31510,G34716);
  not GNAME31511(G31511,G34718);
  not GNAME31512(G31512,G34655);
  not GNAME31513(G31513,G34654);
  not GNAME31514(G31514,G34656);
  not GNAME31515(G31515,G34657);
  not GNAME31516(G31516,G34658);
  not GNAME31517(G31517,G34659);
  not GNAME31518(G31518,G34660);
  not GNAME31519(G31519,G34661);
  not GNAME31520(G31520,G34674);
  not GNAME31521(G31521,G34689);
  not GNAME31522(G31522,G34675);
  not GNAME31523(G31523,G34676);
  not GNAME31524(G31524,G34690);
  not GNAME31525(G31525,G34691);
  not GNAME31526(G31526,G34704);
  not GNAME31527(G31527,G34705);
  not GNAME31528(G31528,G34706);
  not GNAME31529(G31529,G34708);
  not GNAME31530(G31530,G34709);
  not GNAME31531(G31531,G34719);
  not GNAME31532(G31532,G34707);
  not GNAME31533(G31533,G34720);
  not GNAME31534(G31534,G34721);
  not GNAME31535(G31535,G34722);
  not GNAME31536(G31536,G34723);
  not GNAME31537(G31537,G34724);
  not GNAME31538(G31538,G28922);
  not GNAME31539(G31539,G28921);
  not GNAME31540(G31540,G28923);
  not GNAME31541(G31541,G28927);
  not GNAME31542(G31542,G28928);
  not GNAME31543(G31543,G28929);
  not GNAME31544(G31544,G28933);
  not GNAME31545(G31545,G28934);
  not GNAME31546(G31546,G28935);
  not GNAME31547(G31547,G28939);
  not GNAME31548(G31548,G28940);
  not GNAME31549(G31549,G28941);
  not GNAME31550(G31550,G28945);
  not GNAME31551(G31551,G28946);
  not GNAME31552(G31552,G28947);
  not GNAME31553(G31553,G28951);
  not GNAME31554(G31554,G28952);
  not GNAME31555(G31555,G28953);
  not GNAME31556(G31556,G28960);
  not GNAME31557(G31557,G28961);
  not GNAME31558(G31558,G28962);
  nand GNAME31559(G31559,G28991,G31588);
  nand GNAME31560(G31560,G28992,G31589);
  nand GNAME31561(G31561,G28993,G31590);
  nand GNAME31562(G31562,G28994,G31591);
  nand GNAME31563(G31563,G28995,G31592);
  nand GNAME31564(G31564,G28996,G31593);
  nand GNAME31565(G31565,G28997,G31594);
  nand GNAME31566(G31566,G28998,G31595);
  nand GNAME31567(G31567,G28999,G31596);
  nand GNAME31568(G31568,G29000,G31597);
  nand GNAME31569(G31569,G29001,G31598);
  nand GNAME31570(G31570,G29002,G31599);
  nand GNAME31571(G31571,G29006,G31600);
  nand GNAME31572(G31572,G29003,G31601);
  nand GNAME31573(G31573,G29004,G31602);
  nand GNAME31574(G31574,G29005,G31603);
  nand GNAME31575(G31575,G29007,G31604);
  nand GNAME31576(G31576,G29008,G31605);
  nand GNAME31577(G31577,G31606,G31439);
  nand GNAME31578(G31578,G31607,G31440);
  nand GNAME31579(G31579,G31608,G31441);
  nand GNAME31580(G31580,G29009,G31609);
  nand GNAME31581(G31581,G29010,G31610);
  nand GNAME31582(G31582,G29011,G31611);
  xor GNAME31583(G31583,G31706,G31680);
  xor GNAME31584(G31584,G28601,G34345);
  xor GNAME31585(G31585,G28583,G34332);
  xor GNAME31586(G31586,G28589,G34358);
  xor GNAME31587(G31587,G34592,G26201);
  xor GNAME31588(G31588,G2678,G2699);
  xor GNAME31589(G31589,G2262,G2283);
  xor GNAME31590(G31590,G1846,G1867);
  xor GNAME31591(G31591,G2636,G2657);
  xor GNAME31592(G31592,G2220,G2241);
  xor GNAME31593(G31593,G1804,G1825);
  xor GNAME31594(G31594,G2552,G2573);
  xor GNAME31595(G31595,G2136,G2157);
  xor GNAME31596(G31596,G1720,G1741);
  xor GNAME31597(G31597,G2594,G2615);
  xor GNAME31598(G31598,G2178,G2199);
  xor GNAME31599(G31599,G1762,G1783);
  xor GNAME31600(G31600,G2428,G2449);
  xor GNAME31601(G31601,G2470,G2491);
  xor GNAME31602(G31602,G2054,G2075);
  xor GNAME31603(G31603,G1638,G1659);
  xor GNAME31604(G31604,G2012,G2033);
  xor GNAME31605(G31605,G1596,G1617);
  xor GNAME31606(G31606,G2344,G2365);
  xor GNAME31607(G31607,G1928,G1949);
  xor GNAME31608(G31608,G1512,G1533);
  xor GNAME31609(G31609,G2386,G2407);
  xor GNAME31610(G31610,G1970,G1991);
  xor GNAME31611(G31611,G1554,G1575);
  xor GNAME31612(G31612,G27857,G27860);
  xor GNAME31613(G31613,G17921,G27933);
  xor GNAME31614(G31614,G24176,G31613);
  xor GNAME31615(G31615,G17906,G27935);
  xor GNAME31616(G31616,G24161,G31615);
  xor GNAME31617(G31617,G17936,G27937);
  xor GNAME31618(G31618,G24191,G31617);
  dff DFF_31627(CK,G31626,G24141);
  and GNAME31628(G31628,G31626,G31629);
  nand GNAME31629(G31629,G80,G31631);
  buf GNAME31630(G31630,G31626);
  buf GNAME31631(G31631,G31621);
  dff DFF_31640(CK,G31639,G24126);
  and GNAME31641(G31641,G31639,G31642);
  nand GNAME31642(G31642,G80,G31644);
  buf GNAME31643(G31643,G31639);
  buf GNAME31644(G31644,G31634);
  dff DFF_31653(CK,G31652,G21846);
  and GNAME31654(G31654,G31652,G31655);
  nand GNAME31655(G31655,G80,G31657);
  buf GNAME31656(G31656,G31652);
  buf GNAME31657(G31657,G31647);
  dff DFF_31666(CK,G31665,G21816);
  and GNAME31667(G31667,G31665,G31668);
  nand GNAME31668(G31668,G80,G31670);
  buf GNAME31669(G31669,G31665);
  buf GNAME31670(G31670,G31660);
  dff DFF_31679(CK,G31678,G27587);
  and GNAME31680(G31680,G31678,G31681);
  nand GNAME31681(G31681,G80,G31683);
  buf GNAME31682(G31682,G31678);
  buf GNAME31683(G31683,G31673);
  dff DFF_31692(CK,G31691,G31583);
  and GNAME31693(G31693,G31691,G31694);
  nand GNAME31694(G31694,G80,G31696);
  buf GNAME31695(G31695,G31691);
  buf GNAME31696(G31696,G31686);
  dff DFF_31705(CK,G31704,G31612);
  and GNAME31706(G31706,G31704,G31707);
  nand GNAME31707(G31707,G80,G31709);
  buf GNAME31708(G31708,G31704);
  buf GNAME31709(G31709,G31699);
  dff DFF_31718(CK,G31717,G24111);
  and GNAME31719(G31719,G31717,G31720);
  nand GNAME31720(G31720,G80,G31722);
  buf GNAME31721(G31721,G31717);
  buf GNAME31722(G31722,G31712);
  dff DFF_31731(CK,G31730,G25806);
  and GNAME31732(G31732,G31730,G31733);
  nand GNAME31733(G31733,G80,G31735);
  buf GNAME31734(G31734,G31730);
  buf GNAME31735(G31735,G31725);
  dff DFF_31744(CK,G31743,G24096);
  and GNAME31745(G31745,G31743,G31746);
  nand GNAME31746(G31746,G80,G31748);
  buf GNAME31747(G31747,G31743);
  buf GNAME31748(G31748,G31738);
  dff DFF_31757(CK,G31756,G25791);
  and GNAME31758(G31758,G31756,G31759);
  nand GNAME31759(G31759,G80,G31761);
  buf GNAME31760(G31760,G31756);
  buf GNAME31761(G31761,G31751);
  dff DFF_31770(CK,G31769,G26226);
  and GNAME31771(G31771,G31769,G31772);
  nand GNAME31772(G31772,G80,G31774);
  buf GNAME31773(G31773,G31769);
  buf GNAME31774(G31774,G31764);
  dff DFF_31783(CK,G31782,G26691);
  and GNAME31784(G31784,G31782,G31785);
  nand GNAME31785(G31785,G80,G31787);
  buf GNAME31786(G31786,G31782);
  buf GNAME31787(G31787,G31777);
  dff DFF_31796(CK,G31795,G26241);
  and GNAME31797(G31797,G31795,G31798);
  nand GNAME31798(G31798,G80,G31800);
  buf GNAME31799(G31799,G31795);
  buf GNAME31800(G31800,G31790);
  dff DFF_31809(CK,G31808,G27584);
  and GNAME31810(G31810,G31808,G31811);
  nand GNAME31811(G31811,G80,G31813);
  buf GNAME31812(G31812,G31808);
  buf GNAME31813(G31813,G31803);
  dff DFF_31822(CK,G31821,G25776);
  and GNAME31823(G31823,G31821,G31824);
  nand GNAME31824(G31824,G80,G31826);
  buf GNAME31825(G31825,G31821);
  buf GNAME31826(G31826,G31816);
  dff DFF_31835(CK,G31834,G25761);
  and GNAME31836(G31836,G31834,G31837);
  nand GNAME31837(G31837,G80,G31839);
  buf GNAME31838(G31838,G31834);
  buf GNAME31839(G31839,G31829);
  dff DFF_31848(CK,G31847,G25746);
  and GNAME31849(G31849,G31847,G31850);
  nand GNAME31850(G31850,G80,G31852);
  buf GNAME31851(G31851,G31847);
  buf GNAME31852(G31852,G31842);
  dff DFF_31861(CK,G31860,G25731);
  and GNAME31862(G31862,G31860,G31863);
  nand GNAME31863(G31863,G80,G31865);
  buf GNAME31864(G31864,G31860);
  buf GNAME31865(G31865,G31855);
  dff DFF_31874(CK,G31873,G26706);
  and GNAME31875(G31875,G31873,G31876);
  nand GNAME31876(G31876,G80,G31878);
  buf GNAME31877(G31877,G31873);
  buf GNAME31878(G31878,G31868);
  dff DFF_31887(CK,G31886,G26721);
  and GNAME31888(G31888,G31886,G31889);
  nand GNAME31889(G31889,G80,G31891);
  buf GNAME31890(G31890,G31886);
  buf GNAME31891(G31891,G31881);
  dff DFF_31900(CK,G31899,G26736);
  and GNAME31901(G31901,G31899,G31902);
  nand GNAME31902(G31902,G80,G31904);
  buf GNAME31903(G31903,G31899);
  buf GNAME31904(G31904,G31894);
  dff DFF_31913(CK,G31912,G26781);
  and GNAME31914(G31914,G31912,G31915);
  nand GNAME31915(G31915,G80,G31917);
  buf GNAME31916(G31916,G31912);
  buf GNAME31917(G31917,G31907);
  dff DFF_31926(CK,G31925,G27581);
  and GNAME31927(G31927,G31925,G31928);
  nand GNAME31928(G31928,G80,G31930);
  buf GNAME31929(G31929,G31925);
  buf GNAME31930(G31930,G31920);
  dff DFF_31939(CK,G31938,G27578);
  and GNAME31940(G31940,G31938,G31941);
  nand GNAME31941(G31941,G80,G31943);
  buf GNAME31942(G31942,G31938);
  buf GNAME31943(G31943,G31933);
  dff DFF_31952(CK,G31951,G25716);
  and GNAME31953(G31953,G31951,G31954);
  nand GNAME31954(G31954,G80,G31956);
  buf GNAME31955(G31955,G31951);
  buf GNAME31956(G31956,G31946);
  dff DFF_31965(CK,G31964,G25701);
  and GNAME31966(G31966,G31964,G31967);
  nand GNAME31967(G31967,G80,G31969);
  buf GNAME31968(G31968,G31964);
  buf GNAME31969(G31969,G31959);
  dff DFF_31978(CK,G31977,G25686);
  and GNAME31979(G31979,G31977,G31980);
  nand GNAME31980(G31980,G80,G31982);
  buf GNAME31981(G31981,G31977);
  buf GNAME31982(G31982,G31972);
  dff DFF_31991(CK,G31990,G25671);
  and GNAME31992(G31992,G31990,G31993);
  nand GNAME31993(G31993,G80,G31995);
  buf GNAME31994(G31994,G31990);
  buf GNAME31995(G31995,G31985);
  dff DFF_32004(CK,G32003,G26751);
  and GNAME32005(G32005,G32003,G32006);
  nand GNAME32006(G32006,G80,G32008);
  buf GNAME32007(G32007,G32003);
  buf GNAME32008(G32008,G31998);
  dff DFF_32017(CK,G32016,G26766);
  and GNAME32018(G32018,G32016,G32019);
  nand GNAME32019(G32019,G80,G32021);
  buf GNAME32020(G32020,G32016);
  buf GNAME32021(G32021,G32011);
  dff DFF_32030(CK,G32029,G26796);
  and GNAME32031(G32031,G32029,G32032);
  nand GNAME32032(G32032,G80,G32034);
  buf GNAME32033(G32033,G32029);
  buf GNAME32034(G32034,G32024);
  dff DFF_32043(CK,G32042,G26841);
  and GNAME32044(G32044,G32042,G32045);
  nand GNAME32045(G32045,G80,G32047);
  buf GNAME32046(G32046,G32042);
  buf GNAME32047(G32047,G32037);
  dff DFF_32056(CK,G32055,G27575);
  and GNAME32057(G32057,G32055,G32058);
  nand GNAME32058(G32058,G80,G32060);
  buf GNAME32059(G32059,G32055);
  buf GNAME32060(G32060,G32050);
  dff DFF_32069(CK,G32068,G27596);
  and GNAME32070(G32070,G32068,G32071);
  nand GNAME32071(G32071,G80,G32073);
  buf GNAME32072(G32072,G32068);
  buf GNAME32073(G32073,G32063);
  dff DFF_32082(CK,G32081,G25656);
  and GNAME32083(G32083,G32081,G32084);
  nand GNAME32084(G32084,G80,G32086);
  buf GNAME32085(G32085,G32081);
  buf GNAME32086(G32086,G32076);
  dff DFF_32095(CK,G32094,G25641);
  and GNAME32096(G32096,G32094,G32097);
  nand GNAME32097(G32097,G80,G32099);
  buf GNAME32098(G32098,G32094);
  buf GNAME32099(G32099,G32089);
  dff DFF_32108(CK,G32107,G25626);
  and GNAME32109(G32109,G32107,G32110);
  nand GNAME32110(G32110,G80,G32112);
  buf GNAME32111(G32111,G32107);
  buf GNAME32112(G32112,G32102);
  dff DFF_32121(CK,G32120,G25611);
  and GNAME32122(G32122,G32120,G32123);
  nand GNAME32123(G32123,G80,G32125);
  buf GNAME32124(G32124,G32120);
  buf GNAME32125(G32125,G32115);
  dff DFF_32134(CK,G32133,G26811);
  and GNAME32135(G32135,G32133,G32136);
  nand GNAME32136(G32136,G80,G32138);
  buf GNAME32137(G32137,G32133);
  buf GNAME32138(G32138,G32128);
  dff DFF_32147(CK,G32146,G26826);
  and GNAME32148(G32148,G32146,G32149);
  nand GNAME32149(G32149,G80,G32151);
  buf GNAME32150(G32150,G32146);
  buf GNAME32151(G32151,G32141);
  dff DFF_32160(CK,G32159,G26856);
  and GNAME32161(G32161,G32159,G32162);
  nand GNAME32162(G32162,G80,G32164);
  buf GNAME32163(G32163,G32159);
  buf GNAME32164(G32164,G32154);
  dff DFF_32173(CK,G32172,G26901);
  and GNAME32174(G32174,G32172,G32175);
  nand GNAME32175(G32175,G80,G32177);
  buf GNAME32176(G32176,G32172);
  buf GNAME32177(G32177,G32167);
  dff DFF_32186(CK,G32185,G27593);
  and GNAME32187(G32187,G32185,G32188);
  nand GNAME32188(G32188,G80,G32190);
  buf GNAME32189(G32189,G32185);
  buf GNAME32190(G32190,G32180);
  dff DFF_32199(CK,G32198,G27590);
  and GNAME32200(G32200,G32198,G32201);
  nand GNAME32201(G32201,G80,G32203);
  buf GNAME32202(G32202,G32198);
  buf GNAME32203(G32203,G32193);
  dff DFF_32212(CK,G32211,G25596);
  and GNAME32213(G32213,G32211,G32214);
  nand GNAME32214(G32214,G80,G32216);
  buf GNAME32215(G32215,G32211);
  buf GNAME32216(G32216,G32206);
  dff DFF_32225(CK,G32224,G26166);
  and GNAME32226(G32226,G32224,G32227);
  nand GNAME32227(G32227,G80,G32229);
  buf GNAME32228(G32228,G32224);
  buf GNAME32229(G32229,G32219);
  dff DFF_32238(CK,G32237,G25581);
  and GNAME32239(G32239,G32237,G32240);
  nand GNAME32240(G32240,G80,G32242);
  buf GNAME32241(G32241,G32237);
  buf GNAME32242(G32242,G32232);
  dff DFF_32251(CK,G32250,G26151);
  and GNAME32252(G32252,G32250,G32253);
  nand GNAME32253(G32253,G80,G32255);
  buf GNAME32254(G32254,G32250);
  buf GNAME32255(G32255,G32245);
  dff DFF_32264(CK,G32263,G26871);
  and GNAME32265(G32265,G32263,G32266);
  nand GNAME32266(G32266,G80,G32268);
  buf GNAME32267(G32267,G32263);
  buf GNAME32268(G32268,G32258);
  dff DFF_32277(CK,G32276,G26886);
  and GNAME32278(G32278,G32276,G32279);
  nand GNAME32279(G32279,G80,G32281);
  buf GNAME32280(G32280,G32276);
  buf GNAME32281(G32281,G32271);
  dff DFF_32290(CK,G32289,G26916);
  and GNAME32291(G32291,G32289,G32292);
  nand GNAME32292(G32292,G80,G32294);
  buf GNAME32293(G32293,G32289);
  buf GNAME32294(G32294,G32284);
  dff DFF_32303(CK,G32302,G26931);
  and GNAME32304(G32304,G32302,G32305);
  nand GNAME32305(G32305,G80,G32307);
  buf GNAME32306(G32306,G32302);
  buf GNAME32307(G32307,G32297);
  dff DFF_32316(CK,G32315,G27599);
  and GNAME32317(G32317,G32315,G32318);
  nand GNAME32318(G32318,G80,G32320);
  buf GNAME32319(G32319,G32315);
  buf GNAME32320(G32320,G32310);
  dff DFF_32329(CK,G32328,G27602);
  and GNAME32330(G32330,G32328,G32331);
  nand GNAME32331(G32331,G80,G32333);
  buf GNAME32332(G32332,G32328);
  buf GNAME32333(G32333,G32323);
  dff DFF_32342(CK,G32341,G26136);
  and GNAME32343(G32343,G32341,G32344);
  nand GNAME32344(G32344,G80,G32346);
  buf GNAME32345(G32345,G32341);
  buf GNAME32346(G32346,G32336);
  dff DFF_32355(CK,G32354,G26121);
  and GNAME32356(G32356,G32354,G32357);
  nand GNAME32357(G32357,G80,G32359);
  buf GNAME32358(G32358,G32354);
  buf GNAME32359(G32359,G32349);
  dff DFF_32368(CK,G32367,G26106);
  and GNAME32369(G32369,G32367,G32370);
  nand GNAME32370(G32370,G80,G32372);
  buf GNAME32371(G32371,G32367);
  buf GNAME32372(G32372,G32362);
  dff DFF_32381(CK,G32380,G26091);
  and GNAME32382(G32382,G32380,G32383);
  nand GNAME32383(G32383,G80,G32385);
  buf GNAME32384(G32384,G32380);
  buf GNAME32385(G32385,G32375);
  dff DFF_32394(CK,G32393,G26946);
  and GNAME32395(G32395,G32393,G32396);
  nand GNAME32396(G32396,G80,G32398);
  buf GNAME32397(G32397,G32393);
  buf GNAME32398(G32398,G32388);
  dff DFF_32407(CK,G32406,G26961);
  and GNAME32408(G32408,G32406,G32409);
  nand GNAME32409(G32409,G80,G32411);
  buf GNAME32410(G32410,G32406);
  buf GNAME32411(G32411,G32401);
  dff DFF_32420(CK,G32419,G26976);
  and GNAME32421(G32421,G32419,G32422);
  nand GNAME32422(G32422,G80,G32424);
  buf GNAME32423(G32423,G32419);
  buf GNAME32424(G32424,G32414);
  dff DFF_32433(CK,G32432,G26991);
  and GNAME32434(G32434,G32432,G32435);
  nand GNAME32435(G32435,G80,G32437);
  buf GNAME32436(G32436,G32432);
  buf GNAME32437(G32437,G32427);
  dff DFF_32446(CK,G32445,G27614);
  and GNAME32447(G32447,G32445,G32448);
  nand GNAME32448(G32448,G80,G32450);
  buf GNAME32449(G32449,G32445);
  buf GNAME32450(G32450,G32440);
  dff DFF_32459(CK,G32458,G27611);
  and GNAME32460(G32460,G32458,G32461);
  nand GNAME32461(G32461,G80,G32463);
  buf GNAME32462(G32462,G32458);
  buf GNAME32463(G32463,G32453);
  dff DFF_32472(CK,G32471,G26076);
  and GNAME32473(G32473,G32471,G32474);
  nand GNAME32474(G32474,G80,G32476);
  buf GNAME32475(G32475,G32471);
  buf GNAME32476(G32476,G32466);
  dff DFF_32485(CK,G32484,G26061);
  and GNAME32486(G32486,G32484,G32487);
  nand GNAME32487(G32487,G80,G32489);
  buf GNAME32488(G32488,G32484);
  buf GNAME32489(G32489,G32479);
  dff DFF_32498(CK,G32497,G26046);
  and GNAME32499(G32499,G32497,G32500);
  nand GNAME32500(G32500,G80,G32502);
  buf GNAME32501(G32501,G32497);
  buf GNAME32502(G32502,G32492);
  dff DFF_32511(CK,G32510,G26031);
  and GNAME32512(G32512,G32510,G32513);
  nand GNAME32513(G32513,G80,G32515);
  buf GNAME32514(G32514,G32510);
  buf GNAME32515(G32515,G32505);
  dff DFF_32524(CK,G32523,G27006);
  and GNAME32525(G32525,G32523,G32526);
  nand GNAME32526(G32526,G80,G32528);
  buf GNAME32527(G32527,G32523);
  buf GNAME32528(G32528,G32518);
  dff DFF_32537(CK,G32536,G27021);
  and GNAME32538(G32538,G32536,G32539);
  nand GNAME32539(G32539,G80,G32541);
  buf GNAME32540(G32540,G32536);
  buf GNAME32541(G32541,G32531);
  dff DFF_32550(CK,G32549,G27036);
  and GNAME32551(G32551,G32549,G32552);
  nand GNAME32552(G32552,G80,G32554);
  buf GNAME32553(G32553,G32549);
  buf GNAME32554(G32554,G32544);
  dff DFF_32563(CK,G32562,G27051);
  and GNAME32564(G32564,G32562,G32565);
  nand GNAME32565(G32565,G80,G32567);
  buf GNAME32566(G32566,G32562);
  buf GNAME32567(G32567,G32557);
  dff DFF_32576(CK,G32575,G27608);
  and GNAME32577(G32577,G32575,G32578);
  nand GNAME32578(G32578,G80,G32580);
  buf GNAME32579(G32579,G32575);
  buf GNAME32580(G32580,G32570);
  dff DFF_32589(CK,G32588,G27605);
  and GNAME32590(G32590,G32588,G32591);
  nand GNAME32591(G32591,G80,G32593);
  buf GNAME32592(G32592,G32588);
  buf GNAME32593(G32593,G32583);
  dff DFF_32602(CK,G32601,G26016);
  and GNAME32603(G32603,G32601,G32604);
  nand GNAME32604(G32604,G80,G32606);
  buf GNAME32605(G32605,G32601);
  buf GNAME32606(G32606,G32596);
  dff DFF_32615(CK,G32614,G26001);
  and GNAME32616(G32616,G32614,G32617);
  nand GNAME32617(G32617,G80,G32619);
  buf GNAME32618(G32618,G32614);
  buf GNAME32619(G32619,G32609);
  dff DFF_32628(CK,G32627,G25986);
  and GNAME32629(G32629,G32627,G32630);
  nand GNAME32630(G32630,G80,G32632);
  buf GNAME32631(G32631,G32627);
  buf GNAME32632(G32632,G32622);
  dff DFF_32641(CK,G32640,G25971);
  and GNAME32642(G32642,G32640,G32643);
  nand GNAME32643(G32643,G80,G32645);
  buf GNAME32644(G32644,G32640);
  buf GNAME32645(G32645,G32635);
  dff DFF_32654(CK,G32653,G27066);
  and GNAME32655(G32655,G32653,G32656);
  nand GNAME32656(G32656,G80,G32658);
  buf GNAME32657(G32657,G32653);
  buf GNAME32658(G32658,G32648);
  dff DFF_32667(CK,G32666,G27081);
  and GNAME32668(G32668,G32666,G32669);
  nand GNAME32669(G32669,G80,G32671);
  buf GNAME32670(G32670,G32666);
  buf GNAME32671(G32671,G32661);
  dff DFF_32680(CK,G32679,G27096);
  and GNAME32681(G32681,G32679,G32682);
  nand GNAME32682(G32682,G80,G32684);
  buf GNAME32683(G32683,G32679);
  buf GNAME32684(G32684,G32674);
  dff DFF_32693(CK,G32692,G27111);
  and GNAME32694(G32694,G32692,G32695);
  nand GNAME32695(G32695,G80,G32697);
  buf GNAME32696(G32696,G32692);
  buf GNAME32697(G32697,G32687);
  dff DFF_32706(CK,G32705,G27629);
  and GNAME32707(G32707,G32705,G32708);
  nand GNAME32708(G32708,G80,G32710);
  buf GNAME32709(G32709,G32705);
  buf GNAME32710(G32710,G32700);
  dff DFF_32719(CK,G32718,G27626);
  and GNAME32720(G32720,G32718,G32721);
  nand GNAME32721(G32721,G80,G32723);
  buf GNAME32722(G32722,G32718);
  buf GNAME32723(G32723,G32713);
  dff DFF_32732(CK,G32731,G25956);
  and GNAME32733(G32733,G32731,G32734);
  nand GNAME32734(G32734,G80,G32736);
  buf GNAME32735(G32735,G32731);
  buf GNAME32736(G32736,G32726);
  dff DFF_32745(CK,G32744,G25566);
  and GNAME32746(G32746,G32744,G32747);
  nand GNAME32747(G32747,G80,G32749);
  buf GNAME32748(G32748,G32744);
  buf GNAME32749(G32749,G32739);
  dff DFF_32758(CK,G32757,G25941);
  and GNAME32759(G32759,G32757,G32760);
  nand GNAME32760(G32760,G80,G32762);
  buf GNAME32761(G32761,G32757);
  buf GNAME32762(G32762,G32752);
  dff DFF_32771(CK,G32770,G25551);
  and GNAME32772(G32772,G32770,G32773);
  nand GNAME32773(G32773,G80,G32775);
  buf GNAME32774(G32774,G32770);
  buf GNAME32775(G32775,G32765);
  dff DFF_32784(CK,G32783,G27126);
  and GNAME32785(G32785,G32783,G32786);
  nand GNAME32786(G32786,G80,G32788);
  buf GNAME32787(G32787,G32783);
  buf GNAME32788(G32788,G32778);
  dff DFF_32797(CK,G32796,G27141);
  and GNAME32798(G32798,G32796,G32799);
  nand GNAME32799(G32799,G80,G32801);
  buf GNAME32800(G32800,G32796);
  buf GNAME32801(G32801,G32791);
  dff DFF_32810(CK,G32809,G27156);
  and GNAME32811(G32811,G32809,G32812);
  nand GNAME32812(G32812,G80,G32814);
  buf GNAME32813(G32813,G32809);
  buf GNAME32814(G32814,G32804);
  dff DFF_32823(CK,G32822,G27171);
  and GNAME32824(G32824,G32822,G32825);
  nand GNAME32825(G32825,G80,G32827);
  buf GNAME32826(G32826,G32822);
  buf GNAME32827(G32827,G32817);
  dff DFF_32836(CK,G32835,G27623);
  and GNAME32837(G32837,G32835,G32838);
  nand GNAME32838(G32838,G80,G32840);
  buf GNAME32839(G32839,G32835);
  buf GNAME32840(G32840,G32830);
  dff DFF_32849(CK,G32848,G27620);
  and GNAME32850(G32850,G32848,G32851);
  nand GNAME32851(G32851,G80,G32853);
  buf GNAME32852(G32852,G32848);
  buf GNAME32853(G32853,G32843);
  dff DFF_32862(CK,G32861,G24081);
  and GNAME32863(G32863,G32861,G32864);
  nand GNAME32864(G32864,G80,G32866);
  buf GNAME32865(G32865,G32861);
  buf GNAME32866(G32866,G32856);
  dff DFF_32875(CK,G32874,G25536);
  and GNAME32876(G32876,G32874,G32877);
  nand GNAME32877(G32877,G80,G32879);
  buf GNAME32878(G32878,G32874);
  buf GNAME32879(G32879,G32869);
  dff DFF_32888(CK,G32887,G25521);
  and GNAME32889(G32889,G32887,G32890);
  nand GNAME32890(G32890,G80,G32892);
  buf GNAME32891(G32891,G32887);
  buf GNAME32892(G32892,G32882);
  dff DFF_32901(CK,G32900,G24066);
  and GNAME32902(G32902,G32900,G32903);
  nand GNAME32903(G32903,G80,G32905);
  buf GNAME32904(G32904,G32900);
  buf GNAME32905(G32905,G32895);
  dff DFF_32914(CK,G32913,G25506);
  and GNAME32915(G32915,G32913,G32916);
  nand GNAME32916(G32916,G80,G32918);
  buf GNAME32917(G32917,G32913);
  buf GNAME32918(G32918,G32908);
  dff DFF_32927(CK,G32926,G25491);
  and GNAME32928(G32928,G32926,G32929);
  nand GNAME32929(G32929,G80,G32931);
  buf GNAME32930(G32930,G32926);
  buf GNAME32931(G32931,G32921);
  dff DFF_32940(CK,G32939,G25476);
  and GNAME32941(G32941,G32939,G32942);
  nand GNAME32942(G32942,G80,G32944);
  buf GNAME32943(G32943,G32939);
  buf GNAME32944(G32944,G32934);
  dff DFF_32953(CK,G32952,G25461);
  and GNAME32954(G32954,G32952,G32955);
  nand GNAME32955(G32955,G80,G32957);
  buf GNAME32956(G32956,G32952);
  buf GNAME32957(G32957,G32947);
  dff DFF_32966(CK,G32965,G25446);
  and GNAME32967(G32967,G32965,G32968);
  nand GNAME32968(G32968,G80,G32970);
  buf GNAME32969(G32969,G32965);
  buf GNAME32970(G32970,G32960);
  dff DFF_32979(CK,G32978,G27186);
  and GNAME32980(G32980,G32978,G32981);
  nand GNAME32981(G32981,G80,G32983);
  buf GNAME32982(G32982,G32978);
  buf GNAME32983(G32983,G32973);
  dff DFF_32992(CK,G32991,G27201);
  and GNAME32993(G32993,G32991,G32994);
  nand GNAME32994(G32994,G80,G32996);
  buf GNAME32995(G32995,G32991);
  buf GNAME32996(G32996,G32986);
  dff DFF_33005(CK,G33004,G27231);
  and GNAME33006(G33006,G33004,G33007);
  nand GNAME33007(G33007,G80,G33009);
  buf GNAME33008(G33008,G33004);
  buf GNAME33009(G33009,G32999);
  dff DFF_33018(CK,G33017,G27246);
  and GNAME33019(G33019,G33017,G33020);
  nand GNAME33020(G33020,G80,G33022);
  buf GNAME33021(G33021,G33017);
  buf GNAME33022(G33022,G33012);
  dff DFF_33031(CK,G33030,G27617);
  and GNAME33032(G33032,G33030,G33033);
  nand GNAME33033(G33033,G80,G33035);
  buf GNAME33034(G33034,G33030);
  buf GNAME33035(G33035,G33025);
  dff DFF_33044(CK,G33043,G27641);
  and GNAME33045(G33045,G33043,G33046);
  nand GNAME33046(G33046,G80,G33048);
  buf GNAME33047(G33047,G33043);
  buf GNAME33048(G33048,G33038);
  dff DFF_33057(CK,G33056,G25431);
  and GNAME33058(G33058,G33056,G33059);
  nand GNAME33059(G33059,G80,G33061);
  buf GNAME33060(G33060,G33056);
  buf GNAME33061(G33061,G33051);
  dff DFF_33070(CK,G33069,G25416);
  and GNAME33071(G33071,G33069,G33072);
  nand GNAME33072(G33072,G80,G33074);
  buf GNAME33073(G33073,G33069);
  buf GNAME33074(G33074,G33064);
  dff DFF_33083(CK,G33082,G25401);
  and GNAME33084(G33084,G33082,G33085);
  nand GNAME33085(G33085,G80,G33087);
  buf GNAME33086(G33086,G33082);
  buf GNAME33087(G33087,G33077);
  dff DFF_33096(CK,G33095,G25386);
  and GNAME33097(G33097,G33095,G33098);
  nand GNAME33098(G33098,G80,G33100);
  buf GNAME33099(G33099,G33095);
  buf GNAME33100(G33100,G33090);
  dff DFF_33109(CK,G33108,G25371);
  and GNAME33110(G33110,G33108,G33111);
  nand GNAME33111(G33111,G80,G33113);
  buf GNAME33112(G33112,G33108);
  buf GNAME33113(G33113,G33103);
  dff DFF_33122(CK,G33121,G25356);
  and GNAME33123(G33123,G33121,G33124);
  nand GNAME33124(G33124,G80,G33126);
  buf GNAME33125(G33125,G33121);
  buf GNAME33126(G33126,G33116);
  dff DFF_33135(CK,G33134,G25341);
  and GNAME33136(G33136,G33134,G33137);
  nand GNAME33137(G33137,G80,G33139);
  buf GNAME33138(G33138,G33134);
  buf GNAME33139(G33139,G33129);
  dff DFF_33148(CK,G33147,G25326);
  and GNAME33149(G33149,G33147,G33150);
  nand GNAME33150(G33150,G80,G33152);
  buf GNAME33151(G33151,G33147);
  buf GNAME33152(G33152,G33142);
  dff DFF_33161(CK,G33160,G27216);
  and GNAME33162(G33162,G33160,G33163);
  nand GNAME33163(G33163,G80,G33165);
  buf GNAME33164(G33164,G33160);
  buf GNAME33165(G33165,G33155);
  dff DFF_33174(CK,G33173,G27261);
  and GNAME33175(G33175,G33173,G33176);
  nand GNAME33176(G33176,G80,G33178);
  buf GNAME33177(G33177,G33173);
  buf GNAME33178(G33178,G33168);
  dff DFF_33187(CK,G33186,G27276);
  and GNAME33188(G33188,G33186,G33189);
  nand GNAME33189(G33189,G80,G33191);
  buf GNAME33190(G33190,G33186);
  buf GNAME33191(G33191,G33181);
  dff DFF_33200(CK,G33199,G27291);
  and GNAME33201(G33201,G33199,G33202);
  nand GNAME33202(G33202,G80,G33204);
  buf GNAME33203(G33203,G33199);
  buf GNAME33204(G33204,G33194);
  dff DFF_33213(CK,G33212,G27306);
  and GNAME33214(G33214,G33212,G33215);
  nand GNAME33215(G33215,G80,G33217);
  buf GNAME33216(G33216,G33212);
  buf GNAME33217(G33217,G33207);
  dff DFF_33226(CK,G33225,G27638);
  and GNAME33227(G33227,G33225,G33228);
  nand GNAME33228(G33228,G80,G33230);
  buf GNAME33229(G33229,G33225);
  buf GNAME33230(G33230,G33220);
  dff DFF_33239(CK,G33238,G27635);
  and GNAME33240(G33240,G33238,G33241);
  nand GNAME33241(G33241,G80,G33243);
  buf GNAME33242(G33242,G33238);
  buf GNAME33243(G33243,G33233);
  dff DFF_33252(CK,G33251,G25311);
  and GNAME33253(G33253,G33251,G33254);
  nand GNAME33254(G33254,G80,G33256);
  buf GNAME33255(G33255,G33251);
  buf GNAME33256(G33256,G33246);
  dff DFF_33265(CK,G33264,G25296);
  and GNAME33266(G33266,G33264,G33267);
  nand GNAME33267(G33267,G80,G33269);
  buf GNAME33268(G33268,G33264);
  buf GNAME33269(G33269,G33259);
  dff DFF_33278(CK,G33277,G25281);
  and GNAME33279(G33279,G33277,G33280);
  nand GNAME33280(G33280,G80,G33282);
  buf GNAME33281(G33281,G33277);
  buf GNAME33282(G33282,G33272);
  dff DFF_33291(CK,G33290,G25926);
  and GNAME33292(G33292,G33290,G33293);
  nand GNAME33293(G33293,G80,G33295);
  buf GNAME33294(G33294,G33290);
  buf GNAME33295(G33295,G33285);
  dff DFF_33304(CK,G33303,G25911);
  and GNAME33305(G33305,G33303,G33306);
  nand GNAME33306(G33306,G80,G33308);
  buf GNAME33307(G33307,G33303);
  buf GNAME33308(G33308,G33298);
  dff DFF_33317(CK,G33316,G25896);
  and GNAME33318(G33318,G33316,G33319);
  nand GNAME33319(G33319,G80,G33321);
  buf GNAME33320(G33320,G33316);
  buf GNAME33321(G33321,G33311);
  dff DFF_33330(CK,G33329,G25881);
  and GNAME33331(G33331,G33329,G33332);
  nand GNAME33332(G33332,G80,G33334);
  buf GNAME33333(G33333,G33329);
  buf GNAME33334(G33334,G33324);
  dff DFF_33343(CK,G33342,G25266);
  and GNAME33344(G33344,G33342,G33345);
  nand GNAME33345(G33345,G80,G33347);
  buf GNAME33346(G33346,G33342);
  buf GNAME33347(G33347,G33337);
  dff DFF_33356(CK,G33355,G25251);
  and GNAME33357(G33357,G33355,G33358);
  nand GNAME33358(G33358,G80,G33360);
  buf GNAME33359(G33359,G33355);
  buf GNAME33360(G33360,G33350);
  dff DFF_33369(CK,G33368,G27321);
  and GNAME33370(G33370,G33368,G33371);
  nand GNAME33371(G33371,G80,G33373);
  buf GNAME33372(G33372,G33368);
  buf GNAME33373(G33373,G33363);
  dff DFF_33382(CK,G33381,G27336);
  and GNAME33383(G33383,G33381,G33384);
  nand GNAME33384(G33384,G80,G33386);
  buf GNAME33385(G33385,G33381);
  buf GNAME33386(G33386,G33376);
  dff DFF_33395(CK,G33394,G27351);
  and GNAME33396(G33396,G33394,G33397);
  nand GNAME33397(G33397,G80,G33399);
  buf GNAME33398(G33398,G33394);
  buf GNAME33399(G33399,G33389);
  dff DFF_33408(CK,G33407,G27366);
  and GNAME33409(G33409,G33407,G33410);
  nand GNAME33410(G33410,G80,G33412);
  buf GNAME33411(G33411,G33407);
  buf GNAME33412(G33412,G33402);
  dff DFF_33421(CK,G33420,G27632);
  and GNAME33422(G33422,G33420,G33423);
  nand GNAME33423(G33423,G80,G33425);
  buf GNAME33424(G33424,G33420);
  buf GNAME33425(G33425,G33415);
  dff DFF_33434(CK,G33433,G27656);
  and GNAME33435(G33435,G33433,G33436);
  nand GNAME33436(G33436,G80,G33438);
  buf GNAME33437(G33437,G33433);
  buf GNAME33438(G33438,G33428);
  dff DFF_33447(CK,G33446,G25236);
  and GNAME33448(G33448,G33446,G33449);
  nand GNAME33449(G33449,G80,G33451);
  buf GNAME33450(G33450,G33446);
  buf GNAME33451(G33451,G33441);
  dff DFF_33460(CK,G33459,G25221);
  and GNAME33461(G33461,G33459,G33462);
  nand GNAME33462(G33462,G80,G33464);
  buf GNAME33463(G33463,G33459);
  buf GNAME33464(G33464,G33454);
  dff DFF_33473(CK,G33472,G25866);
  and GNAME33474(G33474,G33472,G33475);
  nand GNAME33475(G33475,G80,G33477);
  buf GNAME33476(G33476,G33472);
  buf GNAME33477(G33477,G33467);
  dff DFF_33486(CK,G33485,G25851);
  and GNAME33487(G33487,G33485,G33488);
  nand GNAME33488(G33488,G80,G33490);
  buf GNAME33489(G33489,G33485);
  buf GNAME33490(G33490,G33480);
  dff DFF_33499(CK,G33498,G25836);
  and GNAME33500(G33500,G33498,G33501);
  nand GNAME33501(G33501,G80,G33503);
  buf GNAME33502(G33502,G33498);
  buf GNAME33503(G33503,G33493);
  dff DFF_33512(CK,G33511,G25821);
  and GNAME33513(G33513,G33511,G33514);
  nand GNAME33514(G33514,G80,G33516);
  buf GNAME33515(G33515,G33511);
  buf GNAME33516(G33516,G33506);
  dff DFF_33525(CK,G33524,G25206);
  and GNAME33526(G33526,G33524,G33527);
  nand GNAME33527(G33527,G80,G33529);
  buf GNAME33528(G33528,G33524);
  buf GNAME33529(G33529,G33519);
  dff DFF_33538(CK,G33537,G25191);
  and GNAME33539(G33539,G33537,G33540);
  nand GNAME33540(G33540,G80,G33542);
  buf GNAME33541(G33541,G33537);
  buf GNAME33542(G33542,G33532);
  dff DFF_33551(CK,G33550,G27381);
  and GNAME33552(G33552,G33550,G33553);
  nand GNAME33553(G33553,G80,G33555);
  buf GNAME33554(G33554,G33550);
  buf GNAME33555(G33555,G33545);
  dff DFF_33564(CK,G33563,G27396);
  and GNAME33565(G33565,G33563,G33566);
  nand GNAME33566(G33566,G80,G33568);
  buf GNAME33567(G33567,G33563);
  buf GNAME33568(G33568,G33558);
  dff DFF_33577(CK,G33576,G27411);
  and GNAME33578(G33578,G33576,G33579);
  nand GNAME33579(G33579,G80,G33581);
  buf GNAME33580(G33580,G33576);
  buf GNAME33581(G33581,G33571);
  dff DFF_33590(CK,G33589,G27426);
  and GNAME33591(G33591,G33589,G33592);
  nand GNAME33592(G33592,G80,G33594);
  buf GNAME33593(G33593,G33589);
  buf GNAME33594(G33594,G33584);
  dff DFF_33603(CK,G33602,G27653);
  and GNAME33604(G33604,G33602,G33605);
  nand GNAME33605(G33605,G80,G33607);
  buf GNAME33606(G33606,G33602);
  buf GNAME33607(G33607,G33597);
  dff DFF_33616(CK,G33615,G27650);
  and GNAME33617(G33617,G33615,G33618);
  nand GNAME33618(G33618,G80,G33620);
  buf GNAME33619(G33619,G33615);
  buf GNAME33620(G33620,G33610);
  dff DFF_33629(CK,G33628,G24051);
  and GNAME33630(G33630,G33628,G33631);
  nand GNAME33631(G33631,G80,G33633);
  buf GNAME33632(G33632,G33628);
  buf GNAME33633(G33633,G33623);
  dff DFF_33642(CK,G33641,G24036);
  and GNAME33643(G33643,G33641,G33644);
  nand GNAME33644(G33644,G80,G33646);
  buf GNAME33645(G33645,G33641);
  buf GNAME33646(G33646,G33636);
  dff DFF_33655(CK,G33654,G25176);
  and GNAME33656(G33656,G33654,G33657);
  nand GNAME33657(G33657,G80,G33659);
  buf GNAME33658(G33658,G33654);
  buf GNAME33659(G33659,G33649);
  dff DFF_33668(CK,G33667,G25161);
  and GNAME33669(G33669,G33667,G33670);
  nand GNAME33670(G33670,G80,G33672);
  buf GNAME33671(G33671,G33667);
  buf GNAME33672(G33672,G33662);
  dff DFF_33681(CK,G33680,G25146);
  and GNAME33682(G33682,G33680,G33683);
  nand GNAME33683(G33683,G80,G33685);
  buf GNAME33684(G33684,G33680);
  buf GNAME33685(G33685,G33675);
  dff DFF_33694(CK,G33693,G25131);
  and GNAME33695(G33695,G33693,G33696);
  nand GNAME33696(G33696,G80,G33698);
  buf GNAME33697(G33697,G33693);
  buf GNAME33698(G33698,G33688);
  dff DFF_33707(CK,G33706,G25116);
  and GNAME33708(G33708,G33706,G33709);
  nand GNAME33709(G33709,G80,G33711);
  buf GNAME33710(G33710,G33706);
  buf GNAME33711(G33711,G33701);
  dff DFF_33720(CK,G33719,G24021);
  and GNAME33721(G33721,G33719,G33722);
  nand GNAME33722(G33722,G80,G33724);
  buf GNAME33723(G33723,G33719);
  buf GNAME33724(G33724,G33714);
  dff DFF_33733(CK,G33732,G24006);
  and GNAME33734(G33734,G33732,G33735);
  nand GNAME33735(G33735,G80,G33737);
  buf GNAME33736(G33736,G33732);
  buf GNAME33737(G33737,G33727);
  dff DFF_33746(CK,G33745,G27441);
  and GNAME33747(G33747,G33745,G33748);
  nand GNAME33748(G33748,G80,G33750);
  buf GNAME33749(G33749,G33745);
  buf GNAME33750(G33750,G33740);
  dff DFF_33759(CK,G33758,G27456);
  and GNAME33760(G33760,G33758,G33761);
  nand GNAME33761(G33761,G80,G33763);
  buf GNAME33762(G33762,G33758);
  buf GNAME33763(G33763,G33753);
  dff DFF_33772(CK,G33771,G27471);
  and GNAME33773(G33773,G33771,G33774);
  nand GNAME33774(G33774,G80,G33776);
  buf GNAME33775(G33775,G33771);
  buf GNAME33776(G33776,G33766);
  dff DFF_33785(CK,G33784,G27486);
  and GNAME33786(G33786,G33784,G33787);
  nand GNAME33787(G33787,G80,G33789);
  buf GNAME33788(G33788,G33784);
  buf GNAME33789(G33789,G33779);
  dff DFF_33798(CK,G33797,G27647);
  and GNAME33799(G33799,G33797,G33800);
  nand GNAME33800(G33800,G80,G33802);
  buf GNAME33801(G33801,G33797);
  buf GNAME33802(G33802,G33792);
  dff DFF_33811(CK,G33810,G27644);
  and GNAME33812(G33812,G33810,G33813);
  nand GNAME33813(G33813,G80,G33815);
  buf GNAME33814(G33814,G33810);
  buf GNAME33815(G33815,G33805);
  dff DFF_33824(CK,G33823,G23991);
  and GNAME33825(G33825,G33823,G33826);
  nand GNAME33826(G33826,G80,G33828);
  buf GNAME33827(G33827,G33823);
  buf GNAME33828(G33828,G33818);
  dff DFF_33837(CK,G33836,G24186);
  and GNAME33838(G33838,G33836,G33839);
  nand GNAME33839(G33839,G80,G33841);
  buf GNAME33840(G33840,G33836);
  buf GNAME33841(G33841,G33831);
  dff DFF_33850(CK,G33849,G25101);
  and GNAME33851(G33851,G33849,G33852);
  nand GNAME33852(G33852,G80,G33854);
  buf GNAME33853(G33853,G33849);
  buf GNAME33854(G33854,G33844);
  dff DFF_33863(CK,G33862,G25086);
  and GNAME33864(G33864,G33862,G33865);
  nand GNAME33865(G33865,G80,G33867);
  buf GNAME33866(G33866,G33862);
  buf GNAME33867(G33867,G33857);
  dff DFF_33876(CK,G33875,G25071);
  and GNAME33877(G33877,G33875,G33878);
  nand GNAME33878(G33878,G80,G33880);
  buf GNAME33879(G33879,G33875);
  buf GNAME33880(G33880,G33870);
  dff DFF_33889(CK,G33888,G25056);
  and GNAME33890(G33890,G33888,G33891);
  nand GNAME33891(G33891,G80,G33893);
  buf GNAME33892(G33892,G33888);
  buf GNAME33893(G33893,G33883);
  dff DFF_33902(CK,G33901,G23976);
  and GNAME33903(G33903,G33901,G33904);
  nand GNAME33904(G33904,G80,G33906);
  buf GNAME33905(G33905,G33901);
  buf GNAME33906(G33906,G33896);
  dff DFF_33915(CK,G33914,G24171);
  and GNAME33916(G33916,G33914,G33917);
  nand GNAME33917(G33917,G80,G33919);
  buf GNAME33918(G33918,G33914);
  buf GNAME33919(G33919,G33909);
  dff DFF_33928(CK,G33927,G27501);
  and GNAME33929(G33929,G33927,G33930);
  nand GNAME33930(G33930,G80,G33932);
  buf GNAME33931(G33931,G33927);
  buf GNAME33932(G33932,G33922);
  dff DFF_33941(CK,G33940,G26196);
  and GNAME33942(G33942,G33940,G33943);
  nand GNAME33943(G33943,G80,G33945);
  buf GNAME33944(G33944,G33940);
  buf GNAME33945(G33945,G33935);
  dff DFF_33954(CK,G33953,G27516);
  and GNAME33955(G33955,G33953,G33956);
  nand GNAME33956(G33956,G80,G33958);
  buf GNAME33957(G33957,G33953);
  buf GNAME33958(G33958,G33948);
  dff DFF_33967(CK,G33966,G27531);
  and GNAME33968(G33968,G33966,G33969);
  nand GNAME33969(G33969,G80,G33971);
  buf GNAME33970(G33970,G33966);
  buf GNAME33971(G33971,G33961);
  dff DFF_33980(CK,G33979,G27668);
  and GNAME33981(G33981,G33979,G33982);
  nand GNAME33982(G33982,G80,G33984);
  buf GNAME33983(G33983,G33979);
  buf GNAME33984(G33984,G33974);
  dff DFF_33993(CK,G33992,G27665);
  and GNAME33994(G33994,G33992,G33995);
  nand GNAME33995(G33995,G80,G33997);
  buf GNAME33996(G33996,G33992);
  buf GNAME33997(G33997,G33987);
  dff DFF_34006(CK,G34005,G21786);
  and GNAME34007(G34007,G34005,G34008);
  nand GNAME34008(G34008,G80,G34010);
  buf GNAME34009(G34009,G34005);
  buf GNAME34010(G34010,G34000);
  dff DFF_34019(CK,G34018,G28920);
  and GNAME34020(G34020,G34018,G34021);
  nand GNAME34021(G34021,G80,G34023);
  buf GNAME34022(G34022,G34018);
  buf GNAME34023(G34023,G34013);
  dff DFF_34032(CK,G34031,G28025);
  and GNAME34033(G34033,G34031,G34034);
  nand GNAME34034(G34034,G80,G34036);
  buf GNAME34035(G34035,G34031);
  buf GNAME34036(G34036,G34026);
  dff DFF_34045(CK,G34044,G28022);
  and GNAME34046(G34046,G34044,G34047);
  nand GNAME34047(G34047,G80,G34049);
  buf GNAME34048(G34048,G34044);
  buf GNAME34049(G34049,G34039);
  dff DFF_34058(CK,G34057,G28019);
  and GNAME34059(G34059,G34057,G34060);
  nand GNAME34060(G34060,G80,G34062);
  buf GNAME34061(G34061,G34057);
  buf GNAME34062(G34062,G34052);
  dff DFF_34071(CK,G34070,G28016);
  and GNAME34072(G34072,G34070,G34073);
  nand GNAME34073(G34073,G80,G34075);
  buf GNAME34074(G34074,G34070);
  buf GNAME34075(G34075,G34065);
  dff DFF_34084(CK,G34083,G28013);
  and GNAME34085(G34085,G34083,G34086);
  nand GNAME34086(G34086,G80,G34088);
  buf GNAME34087(G34087,G34083);
  buf GNAME34088(G34088,G34078);
  dff DFF_34097(CK,G34096,G28007);
  and GNAME34098(G34098,G34096,G34099);
  nand GNAME34099(G34099,G80,G34101);
  buf GNAME34100(G34100,G34096);
  buf GNAME34101(G34101,G34091);
  dff DFF_34110(CK,G34109,G28010);
  and GNAME34111(G34111,G34109,G34112);
  nand GNAME34112(G34112,G80,G34114);
  buf GNAME34113(G34113,G34109);
  buf GNAME34114(G34114,G34104);
  dff DFF_34123(CK,G34122,G27980);
  and GNAME34124(G34124,G34122,G34125);
  nand GNAME34125(G34125,G80,G34127);
  buf GNAME34126(G34126,G34122);
  buf GNAME34127(G34127,G34117);
  dff DFF_34136(CK,G34135,G27977);
  and GNAME34137(G34137,G34135,G34138);
  nand GNAME34138(G34138,G80,G34140);
  buf GNAME34139(G34139,G34135);
  buf GNAME34140(G34140,G34130);
  dff DFF_34149(CK,G34148,G27974);
  and GNAME34150(G34150,G34148,G34151);
  nand GNAME34151(G34151,G80,G34153);
  buf GNAME34152(G34152,G34148);
  buf GNAME34153(G34153,G34143);
  dff DFF_34162(CK,G34161,G27971);
  and GNAME34163(G34163,G34161,G34164);
  nand GNAME34164(G34164,G80,G34166);
  buf GNAME34165(G34165,G34161);
  buf GNAME34166(G34166,G34156);
  dff DFF_34175(CK,G34174,G27968);
  and GNAME34176(G34176,G34174,G34177);
  nand GNAME34177(G34177,G80,G34179);
  buf GNAME34178(G34178,G34174);
  buf GNAME34179(G34179,G34169);
  dff DFF_34188(CK,G34187,G27965);
  and GNAME34189(G34189,G34187,G34190);
  nand GNAME34190(G34190,G80,G34192);
  buf GNAME34191(G34191,G34187);
  buf GNAME34192(G34192,G34182);
  dff DFF_34201(CK,G34200,G27962);
  and GNAME34202(G34202,G34200,G34203);
  nand GNAME34203(G34203,G80,G34205);
  buf GNAME34204(G34204,G34200);
  buf GNAME34205(G34205,G34195);
  dff DFF_34214(CK,G34213,G27959);
  and GNAME34215(G34215,G34213,G34216);
  nand GNAME34216(G34216,G80,G34218);
  buf GNAME34217(G34217,G34213);
  buf GNAME34218(G34218,G34208);
  dff DFF_34227(CK,G34226,G28004);
  and GNAME34228(G34228,G34226,G34229);
  nand GNAME34229(G34229,G80,G34231);
  buf GNAME34230(G34230,G34226);
  buf GNAME34231(G34231,G34221);
  dff DFF_34240(CK,G34239,G28001);
  and GNAME34241(G34241,G34239,G34242);
  nand GNAME34242(G34242,G80,G34244);
  buf GNAME34243(G34243,G34239);
  buf GNAME34244(G34244,G34234);
  dff DFF_34253(CK,G34252,G27998);
  and GNAME34254(G34254,G34252,G34255);
  nand GNAME34255(G34255,G80,G34257);
  buf GNAME34256(G34256,G34252);
  buf GNAME34257(G34257,G34247);
  dff DFF_34266(CK,G34265,G27995);
  and GNAME34267(G34267,G34265,G34268);
  nand GNAME34268(G34268,G80,G34270);
  buf GNAME34269(G34269,G34265);
  buf GNAME34270(G34270,G34260);
  dff DFF_34279(CK,G34278,G27992);
  and GNAME34280(G34280,G34278,G34281);
  nand GNAME34281(G34281,G80,G34283);
  buf GNAME34282(G34282,G34278);
  buf GNAME34283(G34283,G34273);
  dff DFF_34292(CK,G34291,G27989);
  and GNAME34293(G34293,G34291,G34294);
  nand GNAME34294(G34294,G80,G34296);
  buf GNAME34295(G34295,G34291);
  buf GNAME34296(G34296,G34286);
  dff DFF_34305(CK,G34304,G27986);
  and GNAME34306(G34306,G34304,G34307);
  nand GNAME34307(G34307,G80,G34309);
  buf GNAME34308(G34308,G34304);
  buf GNAME34309(G34309,G34299);
  dff DFF_34318(CK,G34317,G27983);
  and GNAME34319(G34319,G34317,G34320);
  nand GNAME34320(G34320,G80,G34322);
  buf GNAME34321(G34321,G34317);
  buf GNAME34322(G34322,G34312);
  dff DFF_34331(CK,G34330,G31618);
  and GNAME34332(G34332,G34330,G34333);
  nand GNAME34333(G34333,G80,G34335);
  buf GNAME34334(G34334,G34330);
  buf GNAME34335(G34335,G34325);
  dff DFF_34344(CK,G34343,G31616);
  and GNAME34345(G34345,G34343,G34346);
  nand GNAME34346(G34346,G80,G34348);
  buf GNAME34347(G34347,G34343);
  buf GNAME34348(G34348,G34338);
  dff DFF_34357(CK,G34356,G31614);
  and GNAME34358(G34358,G34356,G34359);
  nand GNAME34359(G34359,G80,G34361);
  buf GNAME34360(G34360,G34356);
  buf GNAME34361(G34361,G34351);
  dff DFF_34370(CK,G34369,G23961);
  and GNAME34371(G34371,G34369,G34372);
  nand GNAME34372(G34372,G80,G34374);
  buf GNAME34373(G34373,G34369);
  buf GNAME34374(G34374,G34364);
  dff DFF_34383(CK,G34382,G23946);
  and GNAME34384(G34384,G34382,G34385);
  nand GNAME34385(G34385,G80,G34387);
  buf GNAME34386(G34386,G34382);
  buf GNAME34387(G34387,G34377);
  dff DFF_34396(CK,G34395,G23931);
  and GNAME34397(G34397,G34395,G34398);
  nand GNAME34398(G34398,G80,G34400);
  buf GNAME34399(G34399,G34395);
  buf GNAME34400(G34400,G34390);
  dff DFF_34409(CK,G34408,G24156);
  and GNAME34410(G34410,G34408,G34411);
  nand GNAME34411(G34411,G80,G34413);
  buf GNAME34412(G34412,G34408);
  buf GNAME34413(G34413,G34403);
  dff DFF_34422(CK,G34421,G27546);
  and GNAME34423(G34423,G34421,G34424);
  nand GNAME34424(G34424,G80,G34426);
  buf GNAME34425(G34425,G34421);
  buf GNAME34426(G34426,G34416);
  dff DFF_34435(CK,G34434,G27561);
  and GNAME34436(G34436,G34434,G34437);
  nand GNAME34437(G34437,G80,G34439);
  buf GNAME34438(G34438,G34434);
  buf GNAME34439(G34439,G34429);
  dff DFF_34448(CK,G34447,G27662);
  and GNAME34449(G34449,G34447,G34450);
  nand GNAME34450(G34450,G80,G34452);
  buf GNAME34451(G34451,G34447);
  buf GNAME34452(G34452,G34442);
  dff DFF_34461(CK,G34460,G27659);
  and GNAME34462(G34462,G34460,G34463);
  nand GNAME34463(G34463,G80,G34465);
  buf GNAME34464(G34464,G34460);
  buf GNAME34465(G34465,G34455);
  dff DFF_34474(CK,G34473,G31587);
  and GNAME34475(G34475,G34473,G34476);
  nand GNAME34476(G34476,G80,G34478);
  buf GNAME34477(G34477,G34473);
  buf GNAME34478(G34478,G34468);
  dff DFF_34487(CK,G34486,G28046);
  and GNAME34488(G34488,G34486,G34489);
  nand GNAME34489(G34489,G80,G34491);
  buf GNAME34490(G34490,G34486);
  buf GNAME34491(G34491,G34481);
  dff DFF_34500(CK,G34499,G28043);
  and GNAME34501(G34501,G34499,G34502);
  nand GNAME34502(G34502,G80,G34504);
  buf GNAME34503(G34503,G34499);
  buf GNAME34504(G34504,G34494);
  dff DFF_34513(CK,G34512,G28040);
  and GNAME34514(G34514,G34512,G34515);
  nand GNAME34515(G34515,G80,G34517);
  buf GNAME34516(G34516,G34512);
  buf GNAME34517(G34517,G34507);
  dff DFF_34526(CK,G34525,G28037);
  and GNAME34527(G34527,G34525,G34528);
  nand GNAME34528(G34528,G80,G34530);
  buf GNAME34529(G34529,G34525);
  buf GNAME34530(G34530,G34520);
  dff DFF_34539(CK,G34538,G28034);
  and GNAME34540(G34540,G34538,G34541);
  nand GNAME34541(G34541,G80,G34543);
  buf GNAME34542(G34542,G34538);
  buf GNAME34543(G34543,G34533);
  dff DFF_34552(CK,G34551,G28031);
  and GNAME34553(G34553,G34551,G34554);
  nand GNAME34554(G34554,G80,G34556);
  buf GNAME34555(G34555,G34551);
  buf GNAME34556(G34556,G34546);
  dff DFF_34565(CK,G34564,G28028);
  and GNAME34566(G34566,G34564,G34567);
  nand GNAME34567(G34567,G80,G34569);
  buf GNAME34568(G34568,G34564);
  buf GNAME34569(G34569,G34559);
  dff DFF_34578(CK,G34577,G34725);
  and GNAME34579(G34579,G34577,G34580);
  nand GNAME34580(G34580,G80,G34582);
  buf GNAME34581(G34581,G34577);
  buf GNAME34582(G34582,G34572);
  dff DFF_34591(CK,G34590,G27566);
  and GNAME34592(G34592,G34590,G34593);
  nand GNAME34593(G34593,G80,G34595);
  buf GNAME34594(G34594,G34590);
  buf GNAME34595(G34595,G34585);
  buf GNAME34596(G34596,G34007);
  buf GNAME34597(G34597,G34007);
  buf GNAME34598(G34598,G2699);
  buf GNAME34599(G34599,G2283);
  buf GNAME34600(G34600,G1867);
  buf GNAME34601(G34601,G9626);
  buf GNAME34602(G34602,G7754);
  buf GNAME34603(G34603,G5882);
  buf GNAME34604(G34604,G2657);
  buf GNAME34605(G34605,G2241);
  buf GNAME34606(G34606,G1825);
  buf GNAME34607(G34607,G9584);
  buf GNAME34608(G34608,G7712);
  buf GNAME34609(G34609,G5840);
  buf GNAME34610(G34610,G9605);
  buf GNAME34611(G34611,G7733);
  buf GNAME34612(G34612,G5861);
  buf GNAME34613(G34613,G2615);
  buf GNAME34614(G34614,G2199);
  buf GNAME34615(G34615,G1783);
  buf GNAME34616(G34616,G9542);
  buf GNAME34617(G34617,G7670);
  buf GNAME34618(G34618,G5798);
  buf GNAME34619(G34619,G9563);
  buf GNAME34620(G34620,G7691);
  buf GNAME34621(G34621,G5819);
  buf GNAME34622(G34622,G2573);
  buf GNAME34623(G34623,G2157);
  buf GNAME34624(G34624,G1741);
  buf GNAME34625(G34625,G9500);
  buf GNAME34626(G34626,G7628);
  buf GNAME34627(G34627,G5756);
  buf GNAME34628(G34628,G9521);
  buf GNAME34629(G34629,G7649);
  buf GNAME34630(G34630,G5777);
  buf GNAME34631(G34631,G2491);
  buf GNAME34632(G34632,G2075);
  buf GNAME34633(G34633,G1659);
  buf GNAME34634(G34634,G9418);
  buf GNAME34635(G34635,G7546);
  buf GNAME34636(G34636,G5674);
  buf GNAME34637(G34637,G9479);
  buf GNAME34638(G34638,G7607);
  buf GNAME34639(G34639,G5735);
  buf GNAME34640(G34640,G2449);
  buf GNAME34641(G34641,G2033);
  buf GNAME34642(G34642,G1617);
  buf GNAME34643(G34643,G9376);
  buf GNAME34644(G34644,G9397);
  buf GNAME34645(G34645,G7504);
  buf GNAME34646(G34646,G7525);
  buf GNAME34647(G34647,G5632);
  buf GNAME34648(G34648,G5653);
  buf GNAME34649(G34649,G2407);
  buf GNAME34650(G34650,G1991);
  buf GNAME34651(G34651,G1575);
  buf GNAME34652(G34652,G31667);
  buf GNAME34653(G34653,G31654);
  buf GNAME34654(G34654,G2699);
  buf GNAME34655(G34655,G2283);
  buf GNAME34656(G34656,G1867);
  buf GNAME34657(G34657,G2657);
  buf GNAME34658(G34658,G2241);
  buf GNAME34659(G34659,G1825);
  buf GNAME34660(G34660,G31667);
  buf GNAME34661(G34661,G31654);
  buf GNAME34662(G34662,G9355);
  buf GNAME34663(G34663,G9334);
  buf GNAME34664(G34664,G9313);
  buf GNAME34665(G34665,G7483);
  buf GNAME34666(G34666,G7462);
  buf GNAME34667(G34667,G5611);
  buf GNAME34668(G34668,G5590);
  buf GNAME34669(G34669,G7441);
  buf GNAME34670(G34670,G5569);
  buf GNAME34671(G34671,G2365);
  buf GNAME34672(G34672,G1949);
  buf GNAME34673(G34673,G1533);
  buf GNAME34674(G34674,G2615);
  buf GNAME34675(G34675,G2199);
  buf GNAME34676(G34676,G1783);
  buf GNAME34677(G34677,G9063);
  buf GNAME34678(G34678,G7191);
  buf GNAME34679(G34679,G5319);
  buf GNAME34680(G34680,G9210);
  buf GNAME34681(G34681,G9271);
  buf GNAME34682(G34682,G7338);
  buf GNAME34683(G34683,G7399);
  buf GNAME34684(G34684,G5466);
  buf GNAME34685(G34685,G5527);
  buf GNAME34686(G34686,G9292);
  buf GNAME34687(G34687,G7420);
  buf GNAME34688(G34688,G5548);
  buf GNAME34689(G34689,G2573);
  buf GNAME34690(G34690,G2157);
  buf GNAME34691(G34691,G1741);
  buf GNAME34692(G34692,G9168);
  buf GNAME34693(G34693,G9147);
  buf GNAME34694(G34694,G9126);
  buf GNAME34695(G34695,G9189);
  buf GNAME34696(G34696,G7317);
  buf GNAME34697(G34697,G5445);
  buf GNAME34698(G34698,G7254);
  buf GNAME34699(G34699,G7275);
  buf GNAME34700(G34700,G7296);
  buf GNAME34701(G34701,G5382);
  buf GNAME34702(G34702,G5403);
  buf GNAME34703(G34703,G5424);
  buf GNAME34704(G34704,G2491);
  buf GNAME34705(G34705,G2075);
  buf GNAME34706(G34706,G1659);
  buf GNAME34707(G34707,G2449);
  buf GNAME34708(G34708,G2033);
  buf GNAME34709(G34709,G1617);
  buf GNAME34710(G34710,G9063);
  buf GNAME34711(G34711,G7191);
  buf GNAME34712(G34712,G5319);
  buf GNAME34713(G34713,G9105);
  buf GNAME34714(G34714,G9084);
  buf GNAME34715(G34715,G7233);
  buf GNAME34716(G34716,G7212);
  buf GNAME34717(G34717,G5361);
  buf GNAME34718(G34718,G5340);
  buf GNAME34719(G34719,G2407);
  buf GNAME34720(G34720,G1991);
  buf GNAME34721(G34721,G1575);
  buf GNAME34722(G34722,G2365);
  buf GNAME34723(G34723,G1949);
  buf GNAME34724(G34724,G1533);
  buf GNAME34725(G34725,G28103);
  buf GNAME34726(G34726,G31559);
  buf GNAME34727(G34727,G31560);
  buf GNAME34728(G34728,G31561);
  buf GNAME34729(G34729,G28103);
  buf GNAME34730(G34730,G28103);
  buf GNAME34731(G34731,G28991);
  buf GNAME34732(G34732,G28992);
  buf GNAME34733(G34733,G28993);
  buf GNAME34734(G34734,G31562);
  buf GNAME34735(G34735,G31563);
  buf GNAME34736(G34736,G31564);
  buf GNAME34737(G34737,G28994);
  buf GNAME34738(G34738,G28995);
  buf GNAME34739(G34739,G28996);
  buf GNAME34740(G34740,G31568);
  buf GNAME34741(G34741,G31565);
  buf GNAME34742(G34742,G31569);
  buf GNAME34743(G34743,G31570);
  buf GNAME34744(G34744,G31566);
  buf GNAME34745(G34745,G31567);
  buf GNAME34746(G34746,G29000);
  buf GNAME34747(G34747,G29001);
  buf GNAME34748(G34748,G29002);
  buf GNAME34749(G34749,G29000);
  buf GNAME34750(G34750,G28997);
  buf GNAME34751(G34751,G29001);
  buf GNAME34752(G34752,G29002);
  buf GNAME34753(G34753,G28998);
  buf GNAME34754(G34754,G28999);
  buf GNAME34755(G34755,G31439);
  buf GNAME34756(G34756,G31440);
  buf GNAME34757(G34757,G31441);
  buf GNAME34758(G34758,G31577);
  buf GNAME34759(G34759,G31578);
  buf GNAME34760(G34760,G31579);
  buf GNAME34761(G34761,G31580);
  buf GNAME34762(G34762,G31581);
  buf GNAME34763(G34763,G31582);
  buf GNAME34764(G34764,G31439);
  buf GNAME34765(G34765,G31440);
  buf GNAME34766(G34766,G31441);
  buf GNAME34767(G34767,G31577);
  buf GNAME34768(G34768,G31578);
  buf GNAME34769(G34769,G31579);
  buf GNAME34770(G34770,G31580);
  buf GNAME34771(G34771,G31581);
  buf GNAME34772(G34772,G31582);
  buf GNAME34773(G34773,G29006);
  buf GNAME34774(G34774,G29009);
  buf GNAME34775(G34775,G29007);
  buf GNAME34776(G34776,G29010);
  buf GNAME34777(G34777,G29008);
  buf GNAME34778(G34778,G29011);
  buf GNAME34779(G34779,G29009);
  buf GNAME34780(G34780,G29010);
  buf GNAME34781(G34781,G29011);
  buf GNAME34782(G34782,G31512);
  buf GNAME34783(G34783,G31513);
  buf GNAME34784(G34784,G31514);
  buf GNAME34785(G34785,G31513);
  buf GNAME34786(G34786,G31512);
  buf GNAME34787(G34787,G31514);
  buf GNAME34788(G34788,G31559);
  buf GNAME34789(G34789,G31562);
  buf GNAME34790(G34790,G31560);
  buf GNAME34791(G34791,G31561);
  buf GNAME34792(G34792,G31563);
  buf GNAME34793(G34793,G31564);
  buf GNAME34794(G34794,G28991);
  buf GNAME34795(G34795,G28992);
  buf GNAME34796(G34796,G28993);
  buf GNAME34797(G34797,G31568);
  buf GNAME34798(G34798,G31569);
  buf GNAME34799(G34799,G31570);
  buf GNAME34800(G34800,G28994);
  buf GNAME34801(G34801,G28995);
  buf GNAME34802(G34802,G28996);
  buf GNAME34803(G34803,G31572);
  buf GNAME34804(G34804,G31573);
  buf GNAME34805(G34805,G31574);
  buf GNAME34806(G34806,G31571);
  buf GNAME34807(G34807,G31575);
  buf GNAME34808(G34808,G31576);
  buf GNAME34809(G34809,G28997);
  buf GNAME34810(G34810,G28998);
  buf GNAME34811(G34811,G28999);
  buf GNAME34812(G34812,G29003);
  buf GNAME34813(G34813,G29004);
  buf GNAME34814(G34814,G29005);
  buf GNAME34815(G34815,G31565);
  buf GNAME34816(G34816,G31566);
  buf GNAME34817(G34817,G31567);
  buf GNAME34818(G34818,G31571);
  buf GNAME34819(G34819,G31575);
  buf GNAME34820(G34820,G31576);
  buf GNAME34821(G34821,G31572);
  buf GNAME34822(G34822,G31573);
  buf GNAME34823(G34823,G31574);
  buf GNAME34824(G34824,G29006);
  buf GNAME34825(G34825,G29007);
  buf GNAME34826(G34826,G29008);
  buf GNAME34827(G34827,G29003);
  buf GNAME34828(G34828,G29004);
  buf GNAME34829(G34829,G29005);
  xor GNAME40353(G40353,G40354,G52765);
  xor GNAME40354(G40354,G52054,G52051);
  and GNAME40355(G40355,G52054,G52765);
  and GNAME40356(G40356,G52051,G52765);
  and GNAME40357(G40357,G52054,G52051);
  or GNAME40358(G40358,G40357,G40356,G40355);
  xor GNAME40368(G40368,G40369,G52768);
  xor GNAME40369(G40369,G52055,G52052);
  and GNAME40370(G40370,G52055,G52768);
  and GNAME40371(G40371,G52052,G52768);
  and GNAME40372(G40372,G52055,G52052);
  or GNAME40373(G40373,G40372,G40371,G40370);
  xor GNAME40383(G40383,G40384,G52771);
  xor GNAME40384(G40384,G52056,G52053);
  and GNAME40385(G40385,G52056,G52771);
  and GNAME40386(G40386,G52053,G52771);
  and GNAME40387(G40387,G52056,G52053);
  or GNAME40388(G40388,G40387,G40386,G40385);
  xor GNAME40398(G40398,G40399,G52774);
  xor GNAME40399(G40399,G52060,G52057);
  and GNAME40400(G40400,G52060,G52774);
  and GNAME40401(G40401,G52057,G52774);
  and GNAME40402(G40402,G52060,G52057);
  or GNAME40403(G40403,G40402,G40401,G40400);
  xor GNAME40413(G40413,G40414,G52777);
  xor GNAME40414(G40414,G52061,G52058);
  and GNAME40415(G40415,G52061,G52777);
  and GNAME40416(G40416,G52058,G52777);
  and GNAME40417(G40417,G52061,G52058);
  or GNAME40418(G40418,G40417,G40416,G40415);
  xor GNAME40428(G40428,G40429,G52780);
  xor GNAME40429(G40429,G52062,G52059);
  and GNAME40430(G40430,G52062,G52780);
  and GNAME40431(G40431,G52059,G52780);
  and GNAME40432(G40432,G52062,G52059);
  or GNAME40433(G40433,G40432,G40431,G40430);
  xor GNAME40443(G40443,G40444,G52783);
  xor GNAME40444(G40444,G52066,G52063);
  and GNAME40445(G40445,G52066,G52783);
  and GNAME40446(G40446,G52063,G52783);
  and GNAME40447(G40447,G52066,G52063);
  or GNAME40448(G40448,G40447,G40446,G40445);
  xor GNAME40458(G40458,G40459,G52786);
  xor GNAME40459(G40459,G52067,G52064);
  and GNAME40460(G40460,G52067,G52786);
  and GNAME40461(G40461,G52064,G52786);
  and GNAME40462(G40462,G52067,G52064);
  or GNAME40463(G40463,G40462,G40461,G40460);
  xor GNAME40473(G40473,G40474,G52789);
  xor GNAME40474(G40474,G52068,G52065);
  and GNAME40475(G40475,G52068,G52789);
  and GNAME40476(G40476,G52065,G52789);
  and GNAME40477(G40477,G52068,G52065);
  or GNAME40478(G40478,G40477,G40476,G40475);
  xor GNAME40488(G40488,G40489,G52792);
  xor GNAME40489(G40489,G52072,G52069);
  and GNAME40490(G40490,G52072,G52792);
  and GNAME40491(G40491,G52069,G52792);
  and GNAME40492(G40492,G52072,G52069);
  or GNAME40493(G40493,G40492,G40491,G40490);
  xor GNAME40503(G40503,G40504,G52795);
  xor GNAME40504(G40504,G52073,G52070);
  and GNAME40505(G40505,G52073,G52795);
  and GNAME40506(G40506,G52070,G52795);
  and GNAME40507(G40507,G52073,G52070);
  or GNAME40508(G40508,G40507,G40506,G40505);
  xor GNAME40518(G40518,G40519,G52798);
  xor GNAME40519(G40519,G52074,G52071);
  and GNAME40520(G40520,G52074,G52798);
  and GNAME40521(G40521,G52071,G52798);
  and GNAME40522(G40522,G52074,G52071);
  or GNAME40523(G40523,G40522,G40521,G40520);
  xor GNAME40533(G40533,G40534,G52801);
  xor GNAME40534(G40534,G52078,G52075);
  and GNAME40535(G40535,G52078,G52801);
  and GNAME40536(G40536,G52075,G52801);
  and GNAME40537(G40537,G52078,G52075);
  or GNAME40538(G40538,G40537,G40536,G40535);
  xor GNAME40548(G40548,G40549,G52804);
  xor GNAME40549(G40549,G52079,G52076);
  and GNAME40550(G40550,G52079,G52804);
  and GNAME40551(G40551,G52076,G52804);
  and GNAME40552(G40552,G52079,G52076);
  or GNAME40553(G40553,G40552,G40551,G40550);
  xor GNAME40563(G40563,G40564,G52807);
  xor GNAME40564(G40564,G52080,G52077);
  and GNAME40565(G40565,G52080,G52807);
  and GNAME40566(G40566,G52077,G52807);
  and GNAME40567(G40567,G52080,G52077);
  or GNAME40568(G40568,G40567,G40566,G40565);
  xor GNAME40578(G40578,G40579,G52810);
  xor GNAME40579(G40579,G52087,G52081);
  and GNAME40580(G40580,G52087,G52810);
  and GNAME40581(G40581,G52081,G52810);
  and GNAME40582(G40582,G52087,G52081);
  or GNAME40583(G40583,G40582,G40581,G40580);
  xor GNAME40593(G40593,G40594,G52813);
  xor GNAME40594(G40594,G52088,G52082);
  and GNAME40595(G40595,G52088,G52813);
  and GNAME40596(G40596,G52082,G52813);
  and GNAME40597(G40597,G52088,G52082);
  or GNAME40598(G40598,G40597,G40596,G40595);
  xor GNAME40608(G40608,G40609,G52816);
  xor GNAME40609(G40609,G52089,G52083);
  and GNAME40610(G40610,G52089,G52816);
  and GNAME40611(G40611,G52083,G52816);
  and GNAME40612(G40612,G52089,G52083);
  or GNAME40613(G40613,G40612,G40611,G40610);
  xor GNAME40623(G40623,G40624,G52819);
  xor GNAME40624(G40624,G52084,G54683);
  and GNAME40625(G40625,G52084,G52819);
  and GNAME40626(G40626,G54683,G52819);
  and GNAME40627(G40627,G52084,G54683);
  or GNAME40628(G40628,G40627,G40626,G40625);
  xor GNAME40638(G40638,G40639,G52822);
  xor GNAME40639(G40639,G52085,G54684);
  and GNAME40640(G40640,G52085,G52822);
  and GNAME40641(G40641,G54684,G52822);
  and GNAME40642(G40642,G52085,G54684);
  or GNAME40643(G40643,G40642,G40641,G40640);
  xor GNAME40653(G40653,G40654,G52825);
  xor GNAME40654(G40654,G52086,G54685);
  and GNAME40655(G40655,G52086,G52825);
  and GNAME40656(G40656,G54685,G52825);
  and GNAME40657(G40657,G52086,G54685);
  or GNAME40658(G40658,G40657,G40656,G40655);
  xor GNAME40668(G40668,G40669,G52828);
  xor GNAME40669(G40669,G51068,G52831);
  and GNAME40670(G40670,G51068,G52828);
  and GNAME40671(G40671,G52831,G52828);
  and GNAME40672(G40672,G51068,G52831);
  or GNAME40673(G40673,G40672,G40671,G40670);
  xor GNAME40683(G40683,G40684,G52834);
  xor GNAME40684(G40684,G51071,G52837);
  and GNAME40685(G40685,G51071,G52834);
  and GNAME40686(G40686,G52837,G52834);
  and GNAME40687(G40687,G51071,G52837);
  or GNAME40688(G40688,G40687,G40686,G40685);
  xor GNAME40698(G40698,G40699,G52840);
  xor GNAME40699(G40699,G51074,G52843);
  and GNAME40700(G40700,G51074,G52840);
  and GNAME40701(G40701,G52843,G52840);
  and GNAME40702(G40702,G51074,G52843);
  or GNAME40703(G40703,G40702,G40701,G40700);
  xor GNAME40713(G40713,G40714,G52846);
  xor GNAME40714(G40714,G51077,G52849);
  and GNAME40715(G40715,G51077,G52846);
  and GNAME40716(G40716,G52849,G52846);
  and GNAME40717(G40717,G51077,G52849);
  or GNAME40718(G40718,G40717,G40716,G40715);
  xor GNAME40728(G40728,G40729,G52852);
  xor GNAME40729(G40729,G51080,G52855);
  and GNAME40730(G40730,G51080,G52852);
  and GNAME40731(G40731,G52855,G52852);
  and GNAME40732(G40732,G51080,G52855);
  or GNAME40733(G40733,G40732,G40731,G40730);
  xor GNAME40743(G40743,G40744,G52858);
  xor GNAME40744(G40744,G51083,G52861);
  and GNAME40745(G40745,G51083,G52858);
  and GNAME40746(G40746,G52861,G52858);
  and GNAME40747(G40747,G51083,G52861);
  or GNAME40748(G40748,G40747,G40746,G40745);
  xor GNAME40758(G40758,G40759,G52900);
  xor GNAME40759(G40759,G51176,G52903);
  and GNAME40760(G40760,G51176,G52900);
  and GNAME40761(G40761,G52903,G52900);
  and GNAME40762(G40762,G51176,G52903);
  or GNAME40763(G40763,G40762,G40761,G40760);
  xor GNAME40773(G40773,G40774,G52906);
  xor GNAME40774(G40774,G51179,G52909);
  and GNAME40775(G40775,G51179,G52906);
  and GNAME40776(G40776,G52909,G52906);
  and GNAME40777(G40777,G51179,G52909);
  or GNAME40778(G40778,G40777,G40776,G40775);
  xor GNAME40788(G40788,G40789,G52912);
  xor GNAME40789(G40789,G51182,G52915);
  and GNAME40790(G40790,G51182,G52912);
  and GNAME40791(G40791,G52915,G52912);
  and GNAME40792(G40792,G51182,G52915);
  or GNAME40793(G40793,G40792,G40791,G40790);
  xor GNAME40803(G40803,G40804,G52936);
  xor GNAME40804(G40804,G51185,G52939);
  and GNAME40805(G40805,G51185,G52936);
  and GNAME40806(G40806,G52939,G52936);
  and GNAME40807(G40807,G51185,G52939);
  or GNAME40808(G40808,G40807,G40806,G40805);
  xor GNAME40818(G40818,G40819,G52942);
  xor GNAME40819(G40819,G51188,G52945);
  and GNAME40820(G40820,G51188,G52942);
  and GNAME40821(G40821,G52945,G52942);
  and GNAME40822(G40822,G51188,G52945);
  or GNAME40823(G40823,G40822,G40821,G40820);
  xor GNAME40833(G40833,G40834,G52948);
  xor GNAME40834(G40834,G51191,G52951);
  and GNAME40835(G40835,G51191,G52948);
  and GNAME40836(G40836,G52951,G52948);
  and GNAME40837(G40837,G51191,G52951);
  or GNAME40838(G40838,G40837,G40836,G40835);
  xor GNAME40848(G40848,G40849,G52972);
  xor GNAME40849(G40849,G51194,G52975);
  and GNAME40850(G40850,G51194,G52972);
  and GNAME40851(G40851,G52975,G52972);
  and GNAME40852(G40852,G51194,G52975);
  or GNAME40853(G40853,G40852,G40851,G40850);
  xor GNAME40863(G40863,G40864,G52978);
  xor GNAME40864(G40864,G51197,G52981);
  and GNAME40865(G40865,G51197,G52978);
  and GNAME40866(G40866,G52981,G52978);
  and GNAME40867(G40867,G51197,G52981);
  or GNAME40868(G40868,G40867,G40866,G40865);
  xor GNAME40878(G40878,G40879,G52984);
  xor GNAME40879(G40879,G51200,G52987);
  and GNAME40880(G40880,G51200,G52984);
  and GNAME40881(G40881,G52987,G52984);
  and GNAME40882(G40882,G51200,G52987);
  or GNAME40883(G40883,G40882,G40881,G40880);
  xor GNAME40893(G40893,G40894,G53008);
  xor GNAME40894(G40894,G51203,G53011);
  and GNAME40895(G40895,G51203,G53008);
  and GNAME40896(G40896,G53011,G53008);
  and GNAME40897(G40897,G51203,G53011);
  or GNAME40898(G40898,G40897,G40896,G40895);
  xor GNAME40908(G40908,G40909,G53014);
  xor GNAME40909(G40909,G51206,G53017);
  and GNAME40910(G40910,G51206,G53014);
  and GNAME40911(G40911,G53017,G53014);
  and GNAME40912(G40912,G51206,G53017);
  or GNAME40913(G40913,G40912,G40911,G40910);
  xor GNAME40923(G40923,G40924,G53020);
  xor GNAME40924(G40924,G51209,G53023);
  and GNAME40925(G40925,G51209,G53020);
  and GNAME40926(G40926,G53023,G53020);
  and GNAME40927(G40927,G51209,G53023);
  or GNAME40928(G40928,G40927,G40926,G40925);
  xor GNAME40938(G40938,G40939,G51343);
  xor GNAME40939(G40939,G53026,G53029);
  and GNAME40940(G40940,G53026,G51343);
  and GNAME40941(G40941,G53029,G51343);
  and GNAME40942(G40942,G53026,G53029);
  or GNAME40943(G40943,G40942,G40941,G40940);
  xor GNAME40953(G40953,G40954,G51349);
  xor GNAME40954(G40954,G53032,G53035);
  and GNAME40955(G40955,G53032,G51349);
  and GNAME40956(G40956,G53035,G51349);
  and GNAME40957(G40957,G53032,G53035);
  or GNAME40958(G40958,G40957,G40956,G40955);
  xor GNAME40968(G40968,G40969,G51355);
  xor GNAME40969(G40969,G53038,G53041);
  and GNAME40970(G40970,G53038,G51355);
  and GNAME40971(G40971,G53041,G51355);
  and GNAME40972(G40972,G53038,G53041);
  or GNAME40973(G40973,G40972,G40971,G40970);
  xor GNAME40983(G40983,G40984,G53044);
  xor GNAME40984(G40984,G51212,G53047);
  and GNAME40985(G40985,G51212,G53044);
  and GNAME40986(G40986,G53047,G53044);
  and GNAME40987(G40987,G51212,G53047);
  or GNAME40988(G40988,G40987,G40986,G40985);
  xor GNAME40998(G40998,G40999,G53050);
  xor GNAME40999(G40999,G51215,G53053);
  and GNAME41000(G41000,G51215,G53050);
  and GNAME41001(G41001,G53053,G53050);
  and GNAME41002(G41002,G51215,G53053);
  or GNAME41003(G41003,G41002,G41001,G41000);
  xor GNAME41013(G41013,G41014,G53056);
  xor GNAME41014(G41014,G51218,G53059);
  and GNAME41015(G41015,G51218,G53056);
  and GNAME41016(G41016,G53059,G53056);
  and GNAME41017(G41017,G51218,G53059);
  or GNAME41018(G41018,G41017,G41016,G41015);
  xor GNAME41028(G41028,G41029,G40358);
  xor GNAME41029(G41029,G54665,G53098);
  and GNAME41030(G41030,G54665,G40358);
  and GNAME41031(G41031,G53098,G40358);
  and GNAME41032(G41032,G54665,G53098);
  or GNAME41033(G41033,G41032,G41031,G41030);
  xor GNAME41043(G41043,G41044,G40373);
  xor GNAME41044(G41044,G54666,G53101);
  and GNAME41045(G41045,G54666,G40373);
  and GNAME41046(G41046,G53101,G40373);
  and GNAME41047(G41047,G54666,G53101);
  or GNAME41048(G41048,G41047,G41046,G41045);
  xor GNAME41058(G41058,G41059,G40388);
  xor GNAME41059(G41059,G54667,G53104);
  and GNAME41060(G41060,G54667,G40388);
  and GNAME41061(G41061,G53104,G40388);
  and GNAME41062(G41062,G54667,G53104);
  or GNAME41063(G41063,G41062,G41061,G41060);
  xor GNAME41073(G41073,G41074,G40353);
  xor GNAME41074(G41074,G52722,G41168);
  and GNAME41075(G41075,G52722,G40353);
  and GNAME41076(G41076,G41168,G40353);
  and GNAME41077(G41077,G52722,G41168);
  or GNAME41078(G41078,G41077,G41076,G41075);
  xor GNAME41088(G41088,G41089,G40368);
  xor GNAME41089(G41089,G52724,G41183);
  and GNAME41090(G41090,G52724,G40368);
  and GNAME41091(G41091,G41183,G40368);
  and GNAME41092(G41092,G52724,G41183);
  or GNAME41093(G41093,G41092,G41091,G41090);
  xor GNAME41103(G41103,G41104,G40383);
  xor GNAME41104(G41104,G52726,G41198);
  and GNAME41105(G41105,G52726,G40383);
  and GNAME41106(G41106,G41198,G40383);
  and GNAME41107(G41107,G52726,G41198);
  or GNAME41108(G41108,G41107,G41106,G41105);
  xor GNAME41118(G41118,G41119,G41213);
  xor GNAME41119(G41119,G40403,G41163);
  and GNAME41120(G41120,G40403,G41213);
  and GNAME41121(G41121,G41163,G41213);
  and GNAME41122(G41122,G40403,G41163);
  or GNAME41123(G41123,G41122,G41121,G41120);
  xor GNAME41133(G41133,G41134,G41228);
  xor GNAME41134(G41134,G40418,G41178);
  and GNAME41135(G41135,G40418,G41228);
  and GNAME41136(G41136,G41178,G41228);
  and GNAME41137(G41137,G40418,G41178);
  or GNAME41138(G41138,G41137,G41136,G41135);
  xor GNAME41148(G41148,G41149,G41243);
  xor GNAME41149(G41149,G40433,G41193);
  and GNAME41150(G41150,G40433,G41243);
  and GNAME41151(G41151,G41193,G41243);
  and GNAME41152(G41152,G40433,G41193);
  or GNAME41153(G41153,G41152,G41151,G41150);
  xor GNAME41163(G41163,G41164,G53110);
  xor GNAME41164(G41164,G54668,G53107);
  and GNAME41165(G41165,G54668,G53110);
  and GNAME41166(G41166,G53107,G53110);
  and GNAME41167(G41167,G54668,G53107);
  or GNAME41168(G41168,G41167,G41166,G41165);
  xor GNAME41178(G41178,G41179,G53116);
  xor GNAME41179(G41179,G54669,G53113);
  and GNAME41180(G41180,G54669,G53116);
  and GNAME41181(G41181,G53113,G53116);
  and GNAME41182(G41182,G54669,G53113);
  or GNAME41183(G41183,G41182,G41181,G41180);
  xor GNAME41193(G41193,G41194,G53122);
  xor GNAME41194(G41194,G54670,G53119);
  and GNAME41195(G41195,G54670,G53122);
  and GNAME41196(G41196,G53119,G53122);
  and GNAME41197(G41197,G54670,G53119);
  or GNAME41198(G41198,G41197,G41196,G41195);
  xor GNAME41208(G41208,G41209,G41348);
  xor GNAME41209(G41209,G53125,G52728);
  and GNAME41210(G41210,G53125,G41348);
  and GNAME41211(G41211,G52728,G41348);
  and GNAME41212(G41212,G53125,G52728);
  or GNAME41213(G41213,G41212,G41211,G41210);
  xor GNAME41223(G41223,G41224,G41363);
  xor GNAME41224(G41224,G53128,G52730);
  and GNAME41225(G41225,G53128,G41363);
  and GNAME41226(G41226,G52730,G41363);
  and GNAME41227(G41227,G53128,G52730);
  or GNAME41228(G41228,G41227,G41226,G41225);
  xor GNAME41238(G41238,G41239,G41378);
  xor GNAME41239(G41239,G53131,G52732);
  and GNAME41240(G41240,G53131,G41378);
  and GNAME41241(G41241,G52732,G41378);
  and GNAME41242(G41242,G53131,G52732);
  or GNAME41243(G41243,G41242,G41241,G41240);
  xor GNAME41253(G41253,G41254,G41208);
  xor GNAME41254(G41254,G40398,G41303);
  and GNAME41255(G41255,G40398,G41208);
  and GNAME41256(G41256,G41303,G41208);
  and GNAME41257(G41257,G40398,G41303);
  or GNAME41258(G41258,G41257,G41256,G41255);
  xor GNAME41268(G41268,G41269,G41223);
  xor GNAME41269(G41269,G40413,G41318);
  and GNAME41270(G41270,G40413,G41223);
  and GNAME41271(G41271,G41318,G41223);
  and GNAME41272(G41272,G40413,G41318);
  or GNAME41273(G41273,G41272,G41271,G41270);
  xor GNAME41283(G41283,G41284,G41238);
  xor GNAME41284(G41284,G40428,G41333);
  and GNAME41285(G41285,G40428,G41238);
  and GNAME41286(G41286,G41333,G41238);
  and GNAME41287(G41287,G40428,G41333);
  or GNAME41288(G41288,G41287,G41286,G41285);
  xor GNAME41298(G41298,G41299,G41393);
  xor GNAME41299(G41299,G53134,G40448);
  and GNAME41300(G41300,G53134,G41393);
  and GNAME41301(G41301,G40448,G41393);
  and GNAME41302(G41302,G53134,G40448);
  or GNAME41303(G41303,G41302,G41301,G41300);
  xor GNAME41313(G41313,G41314,G41408);
  xor GNAME41314(G41314,G53137,G40463);
  and GNAME41315(G41315,G53137,G41408);
  and GNAME41316(G41316,G40463,G41408);
  and GNAME41317(G41317,G53137,G40463);
  or GNAME41318(G41318,G41317,G41316,G41315);
  xor GNAME41328(G41328,G41329,G41423);
  xor GNAME41329(G41329,G53140,G40478);
  and GNAME41330(G41330,G53140,G41423);
  and GNAME41331(G41331,G40478,G41423);
  and GNAME41332(G41332,G53140,G40478);
  or GNAME41333(G41333,G41332,G41331,G41330);
  xor GNAME41343(G41343,G41344,G53146);
  xor GNAME41344(G41344,G54671,G53143);
  and GNAME41345(G41345,G54671,G53146);
  and GNAME41346(G41346,G53143,G53146);
  and GNAME41347(G41347,G54671,G53143);
  or GNAME41348(G41348,G41347,G41346,G41345);
  xor GNAME41358(G41358,G41359,G53152);
  xor GNAME41359(G41359,G54672,G53149);
  and GNAME41360(G41360,G54672,G53152);
  and GNAME41361(G41361,G53149,G53152);
  and GNAME41362(G41362,G54672,G53149);
  or GNAME41363(G41363,G41362,G41361,G41360);
  xor GNAME41373(G41373,G41374,G53158);
  xor GNAME41374(G41374,G54673,G53155);
  and GNAME41375(G41375,G54673,G53158);
  and GNAME41376(G41376,G53155,G53158);
  and GNAME41377(G41377,G54673,G53155);
  or GNAME41378(G41378,G41377,G41376,G41375);
  xor GNAME41388(G41388,G41389,G52734);
  xor GNAME41389(G41389,G53161,G53164);
  and GNAME41390(G41390,G53161,G52734);
  and GNAME41391(G41391,G53164,G52734);
  and GNAME41392(G41392,G53161,G53164);
  or GNAME41393(G41393,G41392,G41391,G41390);
  xor GNAME41403(G41403,G41404,G52736);
  xor GNAME41404(G41404,G53167,G53170);
  and GNAME41405(G41405,G53167,G52736);
  and GNAME41406(G41406,G53170,G52736);
  and GNAME41407(G41407,G53167,G53170);
  or GNAME41408(G41408,G41407,G41406,G41405);
  xor GNAME41418(G41418,G41419,G52738);
  xor GNAME41419(G41419,G53173,G53176);
  and GNAME41420(G41420,G53173,G52738);
  and GNAME41421(G41421,G53176,G52738);
  and GNAME41422(G41422,G53173,G53176);
  or GNAME41423(G41423,G41422,G41421,G41420);
  xor GNAME41433(G41433,G41434,G41388);
  xor GNAME41434(G41434,G41483,G40443);
  and GNAME41435(G41435,G41483,G41388);
  and GNAME41436(G41436,G40443,G41388);
  and GNAME41437(G41437,G41483,G40443);
  or GNAME41438(G41438,G41437,G41436,G41435);
  xor GNAME41448(G41448,G41449,G41403);
  xor GNAME41449(G41449,G41498,G40458);
  and GNAME41450(G41450,G41498,G41403);
  and GNAME41451(G41451,G40458,G41403);
  and GNAME41452(G41452,G41498,G40458);
  or GNAME41453(G41453,G41452,G41451,G41450);
  xor GNAME41463(G41463,G41464,G41418);
  xor GNAME41464(G41464,G41513,G40473);
  and GNAME41465(G41465,G41513,G41418);
  and GNAME41466(G41466,G40473,G41418);
  and GNAME41467(G41467,G41513,G40473);
  or GNAME41468(G41468,G41467,G41466,G41465);
  xor GNAME41478(G41478,G41479,G53182);
  xor GNAME41479(G41479,G54674,G53179);
  and GNAME41480(G41480,G54674,G53182);
  and GNAME41481(G41481,G53179,G53182);
  and GNAME41482(G41482,G54674,G53179);
  or GNAME41483(G41483,G41482,G41481,G41480);
  xor GNAME41493(G41493,G41494,G53188);
  xor GNAME41494(G41494,G54675,G53185);
  and GNAME41495(G41495,G54675,G53188);
  and GNAME41496(G41496,G53185,G53188);
  and GNAME41497(G41497,G54675,G53185);
  or GNAME41498(G41498,G41497,G41496,G41495);
  xor GNAME41508(G41508,G41509,G53194);
  xor GNAME41509(G41509,G54676,G53191);
  and GNAME41510(G41510,G54676,G53194);
  and GNAME41511(G41511,G53191,G53194);
  and GNAME41512(G41512,G54676,G53191);
  or GNAME41513(G41513,G41512,G41511,G41510);
  xor GNAME41523(G41523,G41524,G40493);
  xor GNAME41524(G41524,G53197,G53200);
  and GNAME41525(G41525,G53197,G40493);
  and GNAME41526(G41526,G53200,G40493);
  and GNAME41527(G41527,G53197,G53200);
  or GNAME41528(G41528,G41527,G41526,G41525);
  xor GNAME41538(G41538,G41539,G40508);
  xor GNAME41539(G41539,G53203,G53206);
  and GNAME41540(G41540,G53203,G40508);
  and GNAME41541(G41541,G53206,G40508);
  and GNAME41542(G41542,G53203,G53206);
  or GNAME41543(G41543,G41542,G41541,G41540);
  xor GNAME41553(G41553,G41554,G40523);
  xor GNAME41554(G41554,G53209,G53212);
  and GNAME41555(G41555,G53209,G40523);
  and GNAME41556(G41556,G53212,G40523);
  and GNAME41557(G41557,G53209,G53212);
  or GNAME41558(G41558,G41557,G41556,G41555);
  xor GNAME41568(G41568,G41569,G41663);
  xor GNAME41569(G41569,G40488,G41793);
  and GNAME41570(G41570,G40488,G41663);
  and GNAME41571(G41571,G41793,G41663);
  and GNAME41572(G41572,G40488,G41793);
  or GNAME41573(G41573,G41572,G41571,G41570);
  xor GNAME41583(G41583,G41584,G41678);
  xor GNAME41584(G41584,G40503,G41808);
  and GNAME41585(G41585,G40503,G41678);
  and GNAME41586(G41586,G41808,G41678);
  and GNAME41587(G41587,G40503,G41808);
  or GNAME41588(G41588,G41587,G41586,G41585);
  xor GNAME41598(G41598,G41599,G41693);
  xor GNAME41599(G41599,G40518,G41823);
  and GNAME41600(G41600,G40518,G41693);
  and GNAME41601(G41601,G41823,G41693);
  and GNAME41602(G41602,G40518,G41823);
  or GNAME41603(G41603,G41602,G41601,G41600);
  xor GNAME41613(G41613,G41614,G53218);
  xor GNAME41614(G41614,G54677,G53215);
  and GNAME41615(G41615,G54677,G53218);
  and GNAME41616(G41616,G53215,G53218);
  and GNAME41617(G41617,G54677,G53215);
  or GNAME41618(G41618,G41617,G41616,G41615);
  xor GNAME41628(G41628,G41629,G53224);
  xor GNAME41629(G41629,G54678,G53221);
  and GNAME41630(G41630,G54678,G53224);
  and GNAME41631(G41631,G53221,G53224);
  and GNAME41632(G41632,G54678,G53221);
  or GNAME41633(G41633,G41632,G41631,G41630);
  xor GNAME41643(G41643,G41644,G53230);
  xor GNAME41644(G41644,G54679,G53227);
  and GNAME41645(G41645,G54679,G53230);
  and GNAME41646(G41646,G53227,G53230);
  and GNAME41647(G41647,G54679,G53227);
  or GNAME41648(G41648,G41647,G41646,G41645);
  xor GNAME41658(G41658,G41659,G41613);
  xor GNAME41659(G41659,G40538,G41843);
  and GNAME41660(G41660,G40538,G41613);
  and GNAME41661(G41661,G41843,G41613);
  and GNAME41662(G41662,G40538,G41843);
  or GNAME41663(G41663,G41662,G41661,G41660);
  xor GNAME41673(G41673,G41674,G41628);
  xor GNAME41674(G41674,G40553,G41858);
  and GNAME41675(G41675,G40553,G41628);
  and GNAME41676(G41676,G41858,G41628);
  and GNAME41677(G41677,G40553,G41858);
  or GNAME41678(G41678,G41677,G41676,G41675);
  xor GNAME41688(G41688,G41689,G41643);
  xor GNAME41689(G41689,G40568,G41873);
  and GNAME41690(G41690,G40568,G41643);
  and GNAME41691(G41691,G41873,G41643);
  and GNAME41692(G41692,G40568,G41873);
  or GNAME41693(G41693,G41692,G41691,G41690);
  xor GNAME41703(G41703,G41704,G41753);
  xor GNAME41704(G41704,G53233,G41618);
  and GNAME41705(G41705,G53233,G41753);
  and GNAME41706(G41706,G41618,G41753);
  and GNAME41707(G41707,G53233,G41618);
  or GNAME41708(G41708,G41707,G41706,G41705);
  xor GNAME41718(G41718,G41719,G41768);
  xor GNAME41719(G41719,G53236,G41633);
  and GNAME41720(G41720,G53236,G41768);
  and GNAME41721(G41721,G41633,G41768);
  and GNAME41722(G41722,G53236,G41633);
  or GNAME41723(G41723,G41722,G41721,G41720);
  xor GNAME41733(G41733,G41734,G41783);
  xor GNAME41734(G41734,G53239,G41648);
  and GNAME41735(G41735,G53239,G41783);
  and GNAME41736(G41736,G41648,G41783);
  and GNAME41737(G41737,G53239,G41648);
  or GNAME41738(G41738,G41737,G41736,G41735);
  xor GNAME41748(G41748,G41749,G53248);
  xor GNAME41749(G41749,G53242,G53245);
  and GNAME41750(G41750,G53242,G53248);
  and GNAME41751(G41751,G53245,G53248);
  and GNAME41752(G41752,G53242,G53245);
  or GNAME41753(G41753,G41752,G41751,G41750);
  xor GNAME41763(G41763,G41764,G53257);
  xor GNAME41764(G41764,G53251,G53254);
  and GNAME41765(G41765,G53251,G53257);
  and GNAME41766(G41766,G53254,G53257);
  and GNAME41767(G41767,G53251,G53254);
  or GNAME41768(G41768,G41767,G41766,G41765);
  xor GNAME41778(G41778,G41779,G53266);
  xor GNAME41779(G41779,G53260,G53263);
  and GNAME41780(G41780,G53260,G53266);
  and GNAME41781(G41781,G53263,G53266);
  and GNAME41782(G41782,G53260,G53263);
  or GNAME41783(G41783,G41782,G41781,G41780);
  xor GNAME41793(G41793,G41794,G52740);
  xor GNAME41794(G41794,G53269,G53272);
  and GNAME41795(G41795,G53269,G52740);
  and GNAME41796(G41796,G53272,G52740);
  and GNAME41797(G41797,G53269,G53272);
  or GNAME41798(G41798,G41797,G41796,G41795);
  xor GNAME41808(G41808,G41809,G52742);
  xor GNAME41809(G41809,G53275,G53278);
  and GNAME41810(G41810,G53275,G52742);
  and GNAME41811(G41811,G53278,G52742);
  and GNAME41812(G41812,G53275,G53278);
  or GNAME41813(G41813,G41812,G41811,G41810);
  xor GNAME41823(G41823,G41824,G52744);
  xor GNAME41824(G41824,G53281,G53284);
  and GNAME41825(G41825,G53281,G52744);
  and GNAME41826(G41826,G53284,G52744);
  and GNAME41827(G41827,G53281,G53284);
  or GNAME41828(G41828,G41827,G41826,G41825);
  xor GNAME41838(G41838,G41839,G52746);
  xor GNAME41839(G41839,G53287,G53290);
  and GNAME41840(G41840,G53287,G52746);
  and GNAME41841(G41841,G53290,G52746);
  and GNAME41842(G41842,G53287,G53290);
  or GNAME41843(G41843,G41842,G41841,G41840);
  xor GNAME41853(G41853,G41854,G52748);
  xor GNAME41854(G41854,G53293,G53296);
  and GNAME41855(G41855,G53293,G52748);
  and GNAME41856(G41856,G53296,G52748);
  and GNAME41857(G41857,G53293,G53296);
  or GNAME41858(G41858,G41857,G41856,G41855);
  xor GNAME41868(G41868,G41869,G52750);
  xor GNAME41869(G41869,G53299,G53302);
  and GNAME41870(G41870,G53299,G52750);
  and GNAME41871(G41871,G53302,G52750);
  and GNAME41872(G41872,G53299,G53302);
  or GNAME41873(G41873,G41872,G41871,G41870);
  xor GNAME41883(G41883,G41884,G41933);
  xor GNAME41884(G41884,G53305,G53308);
  and GNAME41885(G41885,G53305,G41933);
  and GNAME41886(G41886,G53308,G41933);
  and GNAME41887(G41887,G53305,G53308);
  or GNAME41888(G41888,G41887,G41886,G41885);
  xor GNAME41898(G41898,G41899,G41948);
  xor GNAME41899(G41899,G53311,G53314);
  and GNAME41900(G41900,G53311,G41948);
  and GNAME41901(G41901,G53314,G41948);
  and GNAME41902(G41902,G53311,G53314);
  or GNAME41903(G41903,G41902,G41901,G41900);
  xor GNAME41913(G41913,G41914,G41963);
  xor GNAME41914(G41914,G53317,G53320);
  and GNAME41915(G41915,G53317,G41963);
  and GNAME41916(G41916,G53320,G41963);
  and GNAME41917(G41917,G53317,G53320);
  or GNAME41918(G41918,G41917,G41916,G41915);
  xor GNAME41928(G41928,G41929,G53326);
  xor GNAME41929(G41929,G54680,G53323);
  and GNAME41930(G41930,G54680,G53326);
  and GNAME41931(G41931,G53323,G53326);
  and GNAME41932(G41932,G54680,G53323);
  or GNAME41933(G41933,G41932,G41931,G41930);
  xor GNAME41943(G41943,G41944,G53332);
  xor GNAME41944(G41944,G54681,G53329);
  and GNAME41945(G41945,G54681,G53332);
  and GNAME41946(G41946,G53329,G53332);
  and GNAME41947(G41947,G54681,G53329);
  or GNAME41948(G41948,G41947,G41946,G41945);
  xor GNAME41958(G41958,G41959,G53338);
  xor GNAME41959(G41959,G54682,G53335);
  and GNAME41960(G41960,G54682,G53338);
  and GNAME41961(G41961,G53335,G53338);
  and GNAME41962(G41962,G54682,G53335);
  or GNAME41963(G41963,G41962,G41961,G41960);
  xor GNAME41973(G41973,G41974,G41838);
  xor GNAME41974(G41974,G42023,G40533);
  and GNAME41975(G41975,G42023,G41838);
  and GNAME41976(G41976,G40533,G41838);
  and GNAME41977(G41977,G42023,G40533);
  or GNAME41978(G41978,G41977,G41976,G41975);
  xor GNAME41988(G41988,G41989,G41853);
  xor GNAME41989(G41989,G42038,G40548);
  and GNAME41990(G41990,G42038,G41853);
  and GNAME41991(G41991,G40548,G41853);
  and GNAME41992(G41992,G42038,G40548);
  or GNAME41993(G41993,G41992,G41991,G41990);
  xor GNAME42003(G42003,G42004,G41868);
  xor GNAME42004(G42004,G42053,G40563);
  and GNAME42005(G42005,G42053,G41868);
  and GNAME42006(G42006,G40563,G41868);
  and GNAME42007(G42007,G42053,G40563);
  or GNAME42008(G42008,G42007,G42006,G42005);
  xor GNAME42018(G42018,G42019,G53347);
  xor GNAME42019(G42019,G53341,G53344);
  and GNAME42020(G42020,G53341,G53347);
  and GNAME42021(G42021,G53344,G53347);
  and GNAME42022(G42022,G53341,G53344);
  or GNAME42023(G42023,G42022,G42021,G42020);
  xor GNAME42033(G42033,G42034,G53356);
  xor GNAME42034(G42034,G53350,G53353);
  and GNAME42035(G42035,G53350,G53356);
  and GNAME42036(G42036,G53353,G53356);
  and GNAME42037(G42037,G53350,G53353);
  or GNAME42038(G42038,G42037,G42036,G42035);
  xor GNAME42048(G42048,G42049,G53365);
  xor GNAME42049(G42049,G53359,G53362);
  and GNAME42050(G42050,G53359,G53365);
  and GNAME42051(G42051,G53362,G53365);
  and GNAME42052(G42052,G53359,G53362);
  or GNAME42053(G42053,G42052,G42051,G42050);
  xor GNAME42063(G42063,G42064,G52752);
  xor GNAME42064(G42064,G53368,G53371);
  and GNAME42065(G42065,G53368,G52752);
  and GNAME42066(G42066,G53371,G52752);
  and GNAME42067(G42067,G53368,G53371);
  or GNAME42068(G42068,G42067,G42066,G42065);
  xor GNAME42078(G42078,G42079,G52754);
  xor GNAME42079(G42079,G53374,G53377);
  and GNAME42080(G42080,G53374,G52754);
  and GNAME42081(G42081,G53377,G52754);
  and GNAME42082(G42082,G53374,G53377);
  or GNAME42083(G42083,G42082,G42081,G42080);
  xor GNAME42093(G42093,G42094,G52756);
  xor GNAME42094(G42094,G53380,G53383);
  and GNAME42095(G42095,G53380,G52756);
  and GNAME42096(G42096,G53383,G52756);
  and GNAME42097(G42097,G53380,G53383);
  or GNAME42098(G42098,G42097,G42096,G42095);
  xor GNAME42108(G42108,G42109,G42068);
  xor GNAME42109(G42109,G53386,G40583);
  and GNAME42110(G42110,G53386,G42068);
  and GNAME42111(G42111,G40583,G42068);
  and GNAME42112(G42112,G53386,G40583);
  or GNAME42113(G42113,G42112,G42111,G42110);
  xor GNAME42123(G42123,G42124,G42218);
  xor GNAME42124(G42124,G40628,G42383);
  and GNAME42125(G42125,G40628,G42218);
  and GNAME42126(G42126,G42383,G42218);
  and GNAME42127(G42127,G40628,G42383);
  or GNAME42128(G42128,G42127,G42126,G42125);
  xor GNAME42138(G42138,G42139,G42083);
  xor GNAME42139(G42139,G53389,G40598);
  and GNAME42140(G42140,G53389,G42083);
  and GNAME42141(G42141,G40598,G42083);
  and GNAME42142(G42142,G53389,G40598);
  or GNAME42143(G42143,G42142,G42141,G42140);
  xor GNAME42153(G42153,G42154,G42098);
  xor GNAME42154(G42154,G53392,G40613);
  and GNAME42155(G42155,G53392,G42098);
  and GNAME42156(G42156,G40613,G42098);
  and GNAME42157(G42157,G53392,G40613);
  or GNAME42158(G42158,G42157,G42156,G42155);
  xor GNAME42168(G42168,G42169,G42263);
  xor GNAME42169(G42169,G40643,G42398);
  and GNAME42170(G42170,G40643,G42263);
  and GNAME42171(G42171,G42398,G42263);
  and GNAME42172(G42172,G40643,G42398);
  or GNAME42173(G42173,G42172,G42171,G42170);
  xor GNAME42183(G42183,G42184,G42278);
  xor GNAME42184(G42184,G40658,G42413);
  and GNAME42185(G42185,G40658,G42278);
  and GNAME42186(G42186,G42413,G42278);
  and GNAME42187(G42187,G40658,G42413);
  or GNAME42188(G42188,G42187,G42186,G42185);
  xor GNAME42198(G42198,G42199,G53401);
  xor GNAME42199(G42199,G53395,G53398);
  and GNAME42200(G42200,G53395,G53401);
  and GNAME42201(G42201,G53398,G53401);
  and GNAME42202(G42202,G53395,G53398);
  or GNAME42203(G42203,G42202,G42201,G42200);
  xor GNAME42213(G42213,G42214,G53410);
  xor GNAME42214(G42214,G53404,G53407);
  and GNAME42215(G42215,G53404,G53410);
  and GNAME42216(G42216,G53407,G53410);
  and GNAME42217(G42217,G53404,G53407);
  or GNAME42218(G42218,G42217,G42216,G42215);
  xor GNAME42228(G42228,G42229,G53419);
  xor GNAME42229(G42229,G53413,G53416);
  and GNAME42230(G42230,G53413,G53419);
  and GNAME42231(G42231,G53416,G53419);
  and GNAME42232(G42232,G53413,G53416);
  or GNAME42233(G42233,G42232,G42231,G42230);
  xor GNAME42243(G42243,G42244,G53428);
  xor GNAME42244(G42244,G53422,G53425);
  and GNAME42245(G42245,G53422,G53428);
  and GNAME42246(G42246,G53425,G53428);
  and GNAME42247(G42247,G53422,G53425);
  or GNAME42248(G42248,G42247,G42246,G42245);
  xor GNAME42258(G42258,G42259,G53437);
  xor GNAME42259(G42259,G53431,G53434);
  and GNAME42260(G42260,G53431,G53437);
  and GNAME42261(G42261,G53434,G53437);
  and GNAME42262(G42262,G53431,G53434);
  or GNAME42263(G42263,G42262,G42261,G42260);
  xor GNAME42273(G42273,G42274,G53446);
  xor GNAME42274(G42274,G53440,G53443);
  and GNAME42275(G42275,G53440,G53446);
  and GNAME42276(G42276,G53443,G53446);
  and GNAME42277(G42277,G53440,G53443);
  or GNAME42278(G42278,G42277,G42276,G42275);
  xor GNAME42288(G42288,G42289,G42063);
  xor GNAME42289(G42289,G40578,G42198);
  and GNAME42290(G42290,G40578,G42063);
  and GNAME42291(G42291,G42198,G42063);
  and GNAME42292(G42292,G40578,G42198);
  or GNAME42293(G42293,G42292,G42291,G42290);
  xor GNAME42303(G42303,G42304,G42378);
  xor GNAME42304(G42304,G40623,G42213);
  and GNAME42305(G42305,G40623,G42378);
  and GNAME42306(G42306,G42213,G42378);
  and GNAME42307(G42307,G40623,G42213);
  or GNAME42308(G42308,G42307,G42306,G42305);
  xor GNAME42318(G42318,G42319,G42078);
  xor GNAME42319(G42319,G40593,G42228);
  and GNAME42320(G42320,G40593,G42078);
  and GNAME42321(G42321,G42228,G42078);
  and GNAME42322(G42322,G40593,G42228);
  or GNAME42323(G42323,G42322,G42321,G42320);
  xor GNAME42333(G42333,G42334,G42393);
  xor GNAME42334(G42334,G40638,G42258);
  and GNAME42335(G42335,G40638,G42393);
  and GNAME42336(G42336,G42258,G42393);
  and GNAME42337(G42337,G40638,G42258);
  or GNAME42338(G42338,G42337,G42336,G42335);
  xor GNAME42348(G42348,G42349,G42093);
  xor GNAME42349(G42349,G40608,G42243);
  and GNAME42350(G42350,G40608,G42093);
  and GNAME42351(G42351,G42243,G42093);
  and GNAME42352(G42352,G40608,G42243);
  or GNAME42353(G42353,G42352,G42351,G42350);
  xor GNAME42363(G42363,G42364,G42408);
  xor GNAME42364(G42364,G40653,G42273);
  and GNAME42365(G42365,G40653,G42408);
  and GNAME42366(G42366,G42273,G42408);
  and GNAME42367(G42367,G40653,G42273);
  or GNAME42368(G42368,G42367,G42366,G42365);
  xor GNAME42378(G42378,G42379,G53455);
  xor GNAME42379(G42379,G53449,G53452);
  and GNAME42380(G42380,G53449,G53455);
  and GNAME42381(G42381,G53452,G53455);
  and GNAME42382(G42382,G53449,G53452);
  or GNAME42383(G42383,G42382,G42381,G42380);
  xor GNAME42393(G42393,G42394,G53464);
  xor GNAME42394(G42394,G53458,G53461);
  and GNAME42395(G42395,G53458,G53464);
  and GNAME42396(G42396,G53461,G53464);
  and GNAME42397(G42397,G53458,G53461);
  or GNAME42398(G42398,G42397,G42396,G42395);
  xor GNAME42408(G42408,G42409,G53473);
  xor GNAME42409(G42409,G53467,G53470);
  and GNAME42410(G42410,G53467,G53473);
  and GNAME42411(G42411,G53470,G53473);
  and GNAME42412(G42412,G53467,G53470);
  or GNAME42413(G42413,G42412,G42411,G42410);
  xor GNAME42423(G42423,G42424,G52758);
  xor GNAME42424(G42424,G53476,G53479);
  and GNAME42425(G42425,G53476,G52758);
  and GNAME42426(G42426,G53479,G52758);
  and GNAME42427(G42427,G53476,G53479);
  or GNAME42428(G42428,G42427,G42426,G42425);
  xor GNAME42438(G42438,G42439,G52760);
  xor GNAME42439(G42439,G53482,G53485);
  and GNAME42440(G42440,G53482,G52760);
  and GNAME42441(G42441,G53485,G52760);
  and GNAME42442(G42442,G53482,G53485);
  or GNAME42443(G42443,G42442,G42441,G42440);
  xor GNAME42453(G42453,G42454,G52762);
  xor GNAME42454(G42454,G53488,G53491);
  and GNAME42455(G42455,G53488,G52762);
  and GNAME42456(G42456,G53491,G52762);
  and GNAME42457(G42457,G53488,G53491);
  or GNAME42458(G42458,G42457,G42456,G42455);
  xor GNAME42468(G42468,G42469,G53500);
  xor GNAME42469(G42469,G53494,G53497);
  and GNAME42470(G42470,G53494,G53500);
  and GNAME42471(G42471,G53497,G53500);
  and GNAME42472(G42472,G53494,G53497);
  or GNAME42473(G42473,G42472,G42471,G42470);
  xor GNAME42483(G42483,G42484,G53509);
  xor GNAME42484(G42484,G53503,G53506);
  and GNAME42485(G42485,G53503,G53509);
  and GNAME42486(G42486,G53506,G53509);
  and GNAME42487(G42487,G53503,G53506);
  or GNAME42488(G42488,G42487,G42486,G42485);
  xor GNAME42498(G42498,G42499,G53518);
  xor GNAME42499(G42499,G53512,G53515);
  and GNAME42500(G42500,G53512,G53518);
  and GNAME42501(G42501,G53515,G53518);
  and GNAME42502(G42502,G53512,G53515);
  or GNAME42503(G42503,G42502,G42501,G42500);
  xor GNAME42513(G42513,G42514,G53521);
  xor GNAME42514(G42514,G52090,G53524);
  and GNAME42515(G42515,G52090,G53521);
  and GNAME42516(G42516,G53524,G53521);
  and GNAME42517(G42517,G52090,G53524);
  or GNAME42518(G42518,G42517,G42516,G42515);
  xor GNAME42528(G42528,G42529,G53527);
  xor GNAME42529(G42529,G52091,G53530);
  and GNAME42530(G42530,G52091,G53527);
  and GNAME42531(G42531,G53530,G53527);
  and GNAME42532(G42532,G52091,G53530);
  or GNAME42533(G42533,G42532,G42531,G42530);
  xor GNAME42543(G42543,G42544,G53533);
  xor GNAME42544(G42544,G52092,G53536);
  and GNAME42545(G42545,G52092,G53533);
  and GNAME42546(G42546,G53536,G53533);
  and GNAME42547(G42547,G52092,G53536);
  or GNAME42548(G42548,G42547,G42546,G42545);
  xor GNAME42558(G42558,G42559,G53542);
  xor GNAME42559(G42559,G54683,G53539);
  and GNAME42560(G42560,G54683,G53542);
  and GNAME42561(G42561,G53539,G53542);
  and GNAME42562(G42562,G54683,G53539);
  or GNAME42563(G42563,G42562,G42561,G42560);
  xor GNAME42573(G42573,G42574,G53548);
  xor GNAME42574(G42574,G54684,G53545);
  and GNAME42575(G42575,G54684,G53548);
  and GNAME42576(G42576,G53545,G53548);
  and GNAME42577(G42577,G54684,G53545);
  or GNAME42578(G42578,G42577,G42576,G42575);
  xor GNAME42588(G42588,G42589,G53554);
  xor GNAME42589(G42589,G54685,G53551);
  and GNAME42590(G42590,G54685,G53554);
  and GNAME42591(G42591,G53551,G53554);
  and GNAME42592(G42592,G54685,G53551);
  or GNAME42593(G42593,G42592,G42591,G42590);
  xor GNAME42603(G42603,G42604,G53563);
  xor GNAME42604(G42604,G53557,G53560);
  and GNAME42605(G42605,G53557,G53563);
  and GNAME42606(G42606,G53560,G53563);
  and GNAME42607(G42607,G53557,G53560);
  or GNAME42608(G42608,G42607,G42606,G42605);
  xor GNAME42618(G42618,G42619,G53572);
  xor GNAME42619(G42619,G53566,G53569);
  and GNAME42620(G42620,G53566,G53572);
  and GNAME42621(G42621,G53569,G53572);
  and GNAME42622(G42622,G53566,G53569);
  or GNAME42623(G42623,G42622,G42621,G42620);
  xor GNAME42633(G42633,G42634,G53581);
  xor GNAME42634(G42634,G53575,G53578);
  and GNAME42635(G42635,G53575,G53581);
  and GNAME42636(G42636,G53578,G53581);
  and GNAME42637(G42637,G53575,G53578);
  or GNAME42638(G42638,G42637,G42636,G42635);
  xor GNAME42648(G42648,G42649,G53590);
  xor GNAME42649(G42649,G53584,G53587);
  and GNAME42650(G42650,G53584,G53590);
  and GNAME42651(G42651,G53587,G53590);
  and GNAME42652(G42652,G53584,G53587);
  or GNAME42653(G42653,G42652,G42651,G42650);
  xor GNAME42663(G42663,G42664,G53599);
  xor GNAME42664(G42664,G53593,G53596);
  and GNAME42665(G42665,G53593,G53599);
  and GNAME42666(G42666,G53596,G53599);
  and GNAME42667(G42667,G53593,G53596);
  or GNAME42668(G42668,G42667,G42666,G42665);
  xor GNAME42678(G42678,G42679,G53608);
  xor GNAME42679(G42679,G53602,G53605);
  and GNAME42680(G42680,G53602,G53608);
  and GNAME42681(G42681,G53605,G53608);
  and GNAME42682(G42682,G53602,G53605);
  or GNAME42683(G42683,G42682,G42681,G42680);
  xor GNAME42693(G42693,G42694,G53617);
  xor GNAME42694(G42694,G53611,G53614);
  and GNAME42695(G42695,G53611,G53617);
  and GNAME42696(G42696,G53614,G53617);
  and GNAME42697(G42697,G53611,G53614);
  or GNAME42698(G42698,G42697,G42696,G42695);
  xor GNAME42708(G42708,G42709,G53626);
  xor GNAME42709(G42709,G53620,G53623);
  and GNAME42710(G42710,G53620,G53626);
  and GNAME42711(G42711,G53623,G53626);
  and GNAME42712(G42712,G53620,G53623);
  or GNAME42713(G42713,G42712,G42711,G42710);
  xor GNAME42723(G42723,G42724,G53635);
  xor GNAME42724(G42724,G53629,G53632);
  and GNAME42725(G42725,G53629,G53635);
  and GNAME42726(G42726,G53632,G53635);
  and GNAME42727(G42727,G53629,G53632);
  or GNAME42728(G42728,G42727,G42726,G42725);
  xor GNAME42738(G42738,G42739,G53644);
  xor GNAME42739(G42739,G53638,G53641);
  and GNAME42740(G42740,G53638,G53644);
  and GNAME42741(G42741,G53641,G53644);
  and GNAME42742(G42742,G53638,G53641);
  or GNAME42743(G42743,G42742,G42741,G42740);
  xor GNAME42753(G42753,G42754,G53653);
  xor GNAME42754(G42754,G53647,G53650);
  and GNAME42755(G42755,G53647,G53653);
  and GNAME42756(G42756,G53650,G53653);
  and GNAME42757(G42757,G53647,G53650);
  or GNAME42758(G42758,G42757,G42756,G42755);
  xor GNAME42768(G42768,G42769,G53662);
  xor GNAME42769(G42769,G53656,G53659);
  and GNAME42770(G42770,G53656,G53662);
  and GNAME42771(G42771,G53659,G53662);
  and GNAME42772(G42772,G53656,G53659);
  or GNAME42773(G42773,G42772,G42771,G42770);
  xor GNAME42783(G42783,G42784,G53665);
  xor GNAME42784(G42784,G52093,G53668);
  and GNAME42785(G42785,G52093,G53665);
  and GNAME42786(G42786,G53668,G53665);
  and GNAME42787(G42787,G52093,G53668);
  or GNAME42788(G42788,G42787,G42786,G42785);
  xor GNAME42798(G42798,G42799,G53671);
  xor GNAME42799(G42799,G52094,G53674);
  and GNAME42800(G42800,G52094,G53671);
  and GNAME42801(G42801,G53674,G53671);
  and GNAME42802(G42802,G52094,G53674);
  or GNAME42803(G42803,G42802,G42801,G42800);
  xor GNAME42813(G42813,G42814,G53677);
  xor GNAME42814(G42814,G52095,G53680);
  and GNAME42815(G42815,G52095,G53677);
  and GNAME42816(G42816,G53680,G53677);
  and GNAME42817(G42817,G52095,G53680);
  or GNAME42818(G42818,G42817,G42816,G42815);
  xor GNAME42828(G42828,G42829,G53683);
  xor GNAME42829(G42829,G52096,G53686);
  and GNAME42830(G42830,G52096,G53683);
  and GNAME42831(G42831,G53686,G53683);
  and GNAME42832(G42832,G52096,G53686);
  or GNAME42833(G42833,G42832,G42831,G42830);
  xor GNAME42843(G42843,G42844,G53689);
  xor GNAME42844(G42844,G52097,G53692);
  and GNAME42845(G42845,G52097,G53689);
  and GNAME42846(G42846,G53692,G53689);
  and GNAME42847(G42847,G52097,G53692);
  or GNAME42848(G42848,G42847,G42846,G42845);
  xor GNAME42858(G42858,G42859,G53695);
  xor GNAME42859(G42859,G52098,G53698);
  and GNAME42860(G42860,G52098,G53695);
  and GNAME42861(G42861,G53698,G53695);
  and GNAME42862(G42862,G52098,G53698);
  or GNAME42863(G42863,G42862,G42861,G42860);
  xor GNAME42873(G42873,G42874,G53707);
  xor GNAME42874(G42874,G53701,G53704);
  and GNAME42875(G42875,G53701,G53707);
  and GNAME42876(G42876,G53704,G53707);
  and GNAME42877(G42877,G53701,G53704);
  or GNAME42878(G42878,G42877,G42876,G42875);
  xor GNAME42888(G42888,G42889,G53716);
  xor GNAME42889(G42889,G53710,G53713);
  and GNAME42890(G42890,G53710,G53716);
  and GNAME42891(G42891,G53713,G53716);
  and GNAME42892(G42892,G53710,G53713);
  or GNAME42893(G42893,G42892,G42891,G42890);
  xor GNAME42903(G42903,G42904,G53725);
  xor GNAME42904(G42904,G53719,G53722);
  and GNAME42905(G42905,G53719,G53725);
  and GNAME42906(G42906,G53722,G53725);
  and GNAME42907(G42907,G53719,G53722);
  or GNAME42908(G42908,G42907,G42906,G42905);
  xor GNAME42918(G42918,G42919,G53734);
  xor GNAME42919(G42919,G53728,G53731);
  and GNAME42920(G42920,G53728,G53734);
  and GNAME42921(G42921,G53731,G53734);
  and GNAME42922(G42922,G53728,G53731);
  or GNAME42923(G42923,G42922,G42921,G42920);
  xor GNAME42933(G42933,G42934,G53743);
  xor GNAME42934(G42934,G53737,G53740);
  and GNAME42935(G42935,G53737,G53743);
  and GNAME42936(G42936,G53740,G53743);
  and GNAME42937(G42937,G53737,G53740);
  or GNAME42938(G42938,G42937,G42936,G42935);
  xor GNAME42948(G42948,G42949,G53752);
  xor GNAME42949(G42949,G53746,G53749);
  and GNAME42950(G42950,G53746,G53752);
  and GNAME42951(G42951,G53749,G53752);
  and GNAME42952(G42952,G53746,G53749);
  or GNAME42953(G42953,G42952,G42951,G42950);
  xor GNAME42963(G42963,G42964,G53761);
  xor GNAME42964(G42964,G53755,G53758);
  and GNAME42965(G42965,G53755,G53761);
  and GNAME42966(G42966,G53758,G53761);
  and GNAME42967(G42967,G53755,G53758);
  or GNAME42968(G42968,G42967,G42966,G42965);
  xor GNAME42978(G42978,G42979,G53770);
  xor GNAME42979(G42979,G53764,G53767);
  and GNAME42980(G42980,G53764,G53770);
  and GNAME42981(G42981,G53767,G53770);
  and GNAME42982(G42982,G53764,G53767);
  or GNAME42983(G42983,G42982,G42981,G42980);
  xor GNAME42993(G42993,G42994,G53779);
  xor GNAME42994(G42994,G53773,G53776);
  and GNAME42995(G42995,G53773,G53779);
  and GNAME42996(G42996,G53776,G53779);
  and GNAME42997(G42997,G53773,G53776);
  or GNAME42998(G42998,G42997,G42996,G42995);
  xor GNAME43008(G43008,G43009,G53788);
  xor GNAME43009(G43009,G53782,G53785);
  and GNAME43010(G43010,G53782,G53788);
  and GNAME43011(G43011,G53785,G53788);
  and GNAME43012(G43012,G53782,G53785);
  or GNAME43013(G43013,G43012,G43011,G43010);
  xor GNAME43023(G43023,G43024,G53797);
  xor GNAME43024(G43024,G53791,G53794);
  and GNAME43025(G43025,G53791,G53797);
  and GNAME43026(G43026,G53794,G53797);
  and GNAME43027(G43027,G53791,G53794);
  or GNAME43028(G43028,G43027,G43026,G43025);
  xor GNAME43038(G43038,G43039,G53806);
  xor GNAME43039(G43039,G53800,G53803);
  and GNAME43040(G43040,G53800,G53806);
  and GNAME43041(G43041,G53803,G53806);
  and GNAME43042(G43042,G53800,G53803);
  or GNAME43043(G43043,G43042,G43041,G43040);
  xor GNAME43053(G43053,G43054,G53809);
  xor GNAME43054(G43054,G52099,G53812);
  and GNAME43055(G43055,G52099,G53809);
  and GNAME43056(G43056,G53812,G53809);
  and GNAME43057(G43057,G52099,G53812);
  or GNAME43058(G43058,G43057,G43056,G43055);
  xor GNAME43068(G43068,G43069,G53815);
  xor GNAME43069(G43069,G52100,G53818);
  and GNAME43070(G43070,G52100,G53815);
  and GNAME43071(G43071,G53818,G53815);
  and GNAME43072(G43072,G52100,G53818);
  or GNAME43073(G43073,G43072,G43071,G43070);
  xor GNAME43083(G43083,G43084,G53821);
  xor GNAME43084(G43084,G52101,G53824);
  and GNAME43085(G43085,G52101,G53821);
  and GNAME43086(G43086,G53824,G53821);
  and GNAME43087(G43087,G52101,G53824);
  or GNAME43088(G43088,G43087,G43086,G43085);
  xor GNAME43098(G43098,G43099,G53827);
  xor GNAME43099(G43099,G52102,G53830);
  and GNAME43100(G43100,G52102,G53827);
  and GNAME43101(G43101,G53830,G53827);
  and GNAME43102(G43102,G52102,G53830);
  or GNAME43103(G43103,G43102,G43101,G43100);
  xor GNAME43113(G43113,G43114,G53833);
  xor GNAME43114(G43114,G52103,G53836);
  and GNAME43115(G43115,G52103,G53833);
  and GNAME43116(G43116,G53836,G53833);
  and GNAME43117(G43117,G52103,G53836);
  or GNAME43118(G43118,G43117,G43116,G43115);
  xor GNAME43128(G43128,G43129,G53839);
  xor GNAME43129(G43129,G52104,G53842);
  and GNAME43130(G43130,G52104,G53839);
  and GNAME43131(G43131,G53842,G53839);
  and GNAME43132(G43132,G52104,G53842);
  or GNAME43133(G43133,G43132,G43131,G43130);
  xor GNAME43143(G43143,G43144,G53851);
  xor GNAME43144(G43144,G53845,G53848);
  and GNAME43145(G43145,G53845,G53851);
  and GNAME43146(G43146,G53848,G53851);
  and GNAME43147(G43147,G53845,G53848);
  or GNAME43148(G43148,G43147,G43146,G43145);
  xor GNAME43158(G43158,G43159,G53860);
  xor GNAME43159(G43159,G53854,G53857);
  and GNAME43160(G43160,G53854,G53860);
  and GNAME43161(G43161,G53857,G53860);
  and GNAME43162(G43162,G53854,G53857);
  or GNAME43163(G43163,G43162,G43161,G43160);
  xor GNAME43173(G43173,G43174,G53869);
  xor GNAME43174(G43174,G53863,G53866);
  and GNAME43175(G43175,G53863,G53869);
  and GNAME43176(G43176,G53866,G53869);
  and GNAME43177(G43177,G53863,G53866);
  or GNAME43178(G43178,G43177,G43176,G43175);
  xor GNAME43188(G43188,G43189,G53878);
  xor GNAME43189(G43189,G53872,G53875);
  and GNAME43190(G43190,G53872,G53878);
  and GNAME43191(G43191,G53875,G53878);
  and GNAME43192(G43192,G53872,G53875);
  or GNAME43193(G43193,G43192,G43191,G43190);
  xor GNAME43203(G43203,G43204,G53887);
  xor GNAME43204(G43204,G53881,G53884);
  and GNAME43205(G43205,G53881,G53887);
  and GNAME43206(G43206,G53884,G53887);
  and GNAME43207(G43207,G53881,G53884);
  or GNAME43208(G43208,G43207,G43206,G43205);
  xor GNAME43218(G43218,G43219,G53896);
  xor GNAME43219(G43219,G53890,G53893);
  and GNAME43220(G43220,G53890,G53896);
  and GNAME43221(G43221,G53893,G53896);
  and GNAME43222(G43222,G53890,G53893);
  or GNAME43223(G43223,G43222,G43221,G43220);
  xor GNAME43233(G43233,G43234,G53905);
  xor GNAME43234(G43234,G53899,G53902);
  and GNAME43235(G43235,G53899,G53905);
  and GNAME43236(G43236,G53902,G53905);
  and GNAME43237(G43237,G53899,G53902);
  or GNAME43238(G43238,G43237,G43236,G43235);
  xor GNAME43248(G43248,G43249,G53914);
  xor GNAME43249(G43249,G53908,G53911);
  and GNAME43250(G43250,G53908,G53914);
  and GNAME43251(G43251,G53911,G53914);
  and GNAME43252(G43252,G53908,G53911);
  or GNAME43253(G43253,G43252,G43251,G43250);
  xor GNAME43263(G43263,G43264,G53923);
  xor GNAME43264(G43264,G53917,G53920);
  and GNAME43265(G43265,G53917,G53923);
  and GNAME43266(G43266,G53920,G53923);
  and GNAME43267(G43267,G53917,G53920);
  or GNAME43268(G43268,G43267,G43266,G43265);
  xor GNAME43278(G43278,G43279,G53932);
  xor GNAME43279(G43279,G53926,G53929);
  and GNAME43280(G43280,G53926,G53932);
  and GNAME43281(G43281,G53929,G53932);
  and GNAME43282(G43282,G53926,G53929);
  or GNAME43283(G43283,G43282,G43281,G43280);
  xor GNAME43293(G43293,G43294,G53941);
  xor GNAME43294(G43294,G53935,G53938);
  and GNAME43295(G43295,G53935,G53941);
  and GNAME43296(G43296,G53938,G53941);
  and GNAME43297(G43297,G53935,G53938);
  or GNAME43298(G43298,G43297,G43296,G43295);
  xor GNAME43308(G43308,G43309,G53950);
  xor GNAME43309(G43309,G53944,G53947);
  and GNAME43310(G43310,G53944,G53950);
  and GNAME43311(G43311,G53947,G53950);
  and GNAME43312(G43312,G53944,G53947);
  or GNAME43313(G43313,G43312,G43311,G43310);
  xor GNAME43323(G43323,G43324,G53953);
  xor GNAME43324(G43324,G52105,G53956);
  and GNAME43325(G43325,G52105,G53953);
  and GNAME43326(G43326,G53956,G53953);
  and GNAME43327(G43327,G52105,G53956);
  or GNAME43328(G43328,G43327,G43326,G43325);
  xor GNAME43338(G43338,G43339,G53959);
  xor GNAME43339(G43339,G52106,G53962);
  and GNAME43340(G43340,G52106,G53959);
  and GNAME43341(G43341,G53962,G53959);
  and GNAME43342(G43342,G52106,G53962);
  or GNAME43343(G43343,G43342,G43341,G43340);
  xor GNAME43353(G43353,G43354,G53965);
  xor GNAME43354(G43354,G52107,G53968);
  and GNAME43355(G43355,G52107,G53965);
  and GNAME43356(G43356,G53968,G53965);
  and GNAME43357(G43357,G52107,G53968);
  or GNAME43358(G43358,G43357,G43356,G43355);
  xor GNAME43368(G43368,G43369,G53971);
  xor GNAME43369(G43369,G52108,G53974);
  and GNAME43370(G43370,G52108,G53971);
  and GNAME43371(G43371,G53974,G53971);
  and GNAME43372(G43372,G52108,G53974);
  or GNAME43373(G43373,G43372,G43371,G43370);
  xor GNAME43383(G43383,G43384,G53977);
  xor GNAME43384(G43384,G52109,G53980);
  and GNAME43385(G43385,G52109,G53977);
  and GNAME43386(G43386,G53980,G53977);
  and GNAME43387(G43387,G52109,G53980);
  or GNAME43388(G43388,G43387,G43386,G43385);
  xor GNAME43398(G43398,G43399,G53983);
  xor GNAME43399(G43399,G52110,G53986);
  and GNAME43400(G43400,G52110,G53983);
  and GNAME43401(G43401,G53986,G53983);
  and GNAME43402(G43402,G52110,G53986);
  or GNAME43403(G43403,G43402,G43401,G43400);
  xor GNAME43413(G43413,G43414,G53995);
  xor GNAME43414(G43414,G53989,G53992);
  and GNAME43415(G43415,G53989,G53995);
  and GNAME43416(G43416,G53992,G53995);
  and GNAME43417(G43417,G53989,G53992);
  or GNAME43418(G43418,G43417,G43416,G43415);
  xor GNAME43428(G43428,G43429,G54004);
  xor GNAME43429(G43429,G53998,G54001);
  and GNAME43430(G43430,G53998,G54004);
  and GNAME43431(G43431,G54001,G54004);
  and GNAME43432(G43432,G53998,G54001);
  or GNAME43433(G43433,G43432,G43431,G43430);
  xor GNAME43443(G43443,G43444,G54013);
  xor GNAME43444(G43444,G54007,G54010);
  and GNAME43445(G43445,G54007,G54013);
  and GNAME43446(G43446,G54010,G54013);
  and GNAME43447(G43447,G54007,G54010);
  or GNAME43448(G43448,G43447,G43446,G43445);
  xor GNAME43458(G43458,G43459,G54022);
  xor GNAME43459(G43459,G54016,G54019);
  and GNAME43460(G43460,G54016,G54022);
  and GNAME43461(G43461,G54019,G54022);
  and GNAME43462(G43462,G54016,G54019);
  or GNAME43463(G43463,G43462,G43461,G43460);
  xor GNAME43473(G43473,G43474,G54031);
  xor GNAME43474(G43474,G54025,G54028);
  and GNAME43475(G43475,G54025,G54031);
  and GNAME43476(G43476,G54028,G54031);
  and GNAME43477(G43477,G54025,G54028);
  or GNAME43478(G43478,G43477,G43476,G43475);
  xor GNAME43488(G43488,G43489,G54040);
  xor GNAME43489(G43489,G54034,G54037);
  and GNAME43490(G43490,G54034,G54040);
  and GNAME43491(G43491,G54037,G54040);
  and GNAME43492(G43492,G54034,G54037);
  or GNAME43493(G43493,G43492,G43491,G43490);
  xor GNAME43503(G43503,G43504,G43568);
  xor GNAME43504(G43504,G40673,G43748);
  and GNAME43505(G43505,G40673,G43568);
  and GNAME43506(G43506,G43748,G43568);
  and GNAME43507(G43507,G40673,G43748);
  or GNAME43508(G43508,G43507,G43506,G43505);
  xor GNAME43518(G43518,G43519,G43613);
  xor GNAME43519(G43519,G40688,G43793);
  and GNAME43520(G43520,G40688,G43613);
  and GNAME43521(G43521,G43793,G43613);
  and GNAME43522(G43522,G40688,G43793);
  or GNAME43523(G43523,G43522,G43521,G43520);
  xor GNAME43533(G43533,G43534,G43628);
  xor GNAME43534(G43534,G40703,G43808);
  and GNAME43535(G43535,G40703,G43628);
  and GNAME43536(G43536,G43808,G43628);
  and GNAME43537(G43537,G40703,G43808);
  or GNAME43538(G43538,G43537,G43536,G43535);
  xor GNAME43548(G43548,G43549,G54049);
  xor GNAME43549(G43549,G54043,G54046);
  and GNAME43550(G43550,G54043,G54049);
  and GNAME43551(G43551,G54046,G54049);
  and GNAME43552(G43552,G54043,G54046);
  or GNAME43553(G43553,G43552,G43551,G43550);
  xor GNAME43563(G43563,G43564,G54058);
  xor GNAME43564(G43564,G54052,G54055);
  and GNAME43565(G43565,G54052,G54058);
  and GNAME43566(G43566,G54055,G54058);
  and GNAME43567(G43567,G54052,G54055);
  or GNAME43568(G43568,G43567,G43566,G43565);
  xor GNAME43578(G43578,G43579,G54067);
  xor GNAME43579(G43579,G54061,G54064);
  and GNAME43580(G43580,G54061,G54067);
  and GNAME43581(G43581,G54064,G54067);
  and GNAME43582(G43582,G54061,G54064);
  or GNAME43583(G43583,G43582,G43581,G43580);
  xor GNAME43593(G43593,G43594,G54076);
  xor GNAME43594(G43594,G54070,G54073);
  and GNAME43595(G43595,G54070,G54076);
  and GNAME43596(G43596,G54073,G54076);
  and GNAME43597(G43597,G54070,G54073);
  or GNAME43598(G43598,G43597,G43596,G43595);
  xor GNAME43608(G43608,G43609,G54085);
  xor GNAME43609(G43609,G54079,G54082);
  and GNAME43610(G43610,G54079,G54085);
  and GNAME43611(G43611,G54082,G54085);
  and GNAME43612(G43612,G54079,G54082);
  or GNAME43613(G43613,G43612,G43611,G43610);
  xor GNAME43623(G43623,G43624,G54094);
  xor GNAME43624(G43624,G54088,G54091);
  and GNAME43625(G43625,G54088,G54094);
  and GNAME43626(G43626,G54091,G54094);
  and GNAME43627(G43627,G54088,G54091);
  or GNAME43628(G43628,G43627,G43626,G43625);
  xor GNAME43638(G43638,G43639,G43743);
  xor GNAME43639(G43639,G40668,G43563);
  and GNAME43640(G43640,G40668,G43743);
  and GNAME43641(G43641,G43563,G43743);
  and GNAME43642(G43642,G40668,G43563);
  or GNAME43643(G43643,G43642,G43641,G43640);
  xor GNAME43653(G43653,G43654,G43788);
  xor GNAME43654(G43654,G40683,G43608);
  and GNAME43655(G43655,G40683,G43788);
  and GNAME43656(G43656,G43608,G43788);
  and GNAME43657(G43657,G40683,G43608);
  or GNAME43658(G43658,G43657,G43656,G43655);
  xor GNAME43668(G43668,G43669,G43803);
  xor GNAME43669(G43669,G40698,G43623);
  and GNAME43670(G43670,G40698,G43803);
  and GNAME43671(G43671,G43623,G43803);
  and GNAME43672(G43672,G40698,G43623);
  or GNAME43673(G43673,G43672,G43671,G43670);
  xor GNAME43683(G43683,G43684,G54097);
  xor GNAME43684(G43684,G52111,G54100);
  and GNAME43685(G43685,G52111,G54097);
  and GNAME43686(G43686,G54100,G54097);
  and GNAME43687(G43687,G52111,G54100);
  or GNAME43688(G43688,G43687,G43686,G43685);
  xor GNAME43698(G43698,G43699,G54103);
  xor GNAME43699(G43699,G52112,G54106);
  and GNAME43700(G43700,G52112,G54103);
  and GNAME43701(G43701,G54106,G54103);
  and GNAME43702(G43702,G52112,G54106);
  or GNAME43703(G43703,G43702,G43701,G43700);
  xor GNAME43713(G43713,G43714,G54109);
  xor GNAME43714(G43714,G52113,G54112);
  and GNAME43715(G43715,G52113,G54109);
  and GNAME43716(G43716,G54112,G54109);
  and GNAME43717(G43717,G52113,G54112);
  or GNAME43718(G43718,G43717,G43716,G43715);
  xor GNAME43728(G43728,G43729,G54121);
  xor GNAME43729(G43729,G54115,G54118);
  and GNAME43730(G43730,G54115,G54121);
  and GNAME43731(G43731,G54118,G54121);
  and GNAME43732(G43732,G54115,G54118);
  or GNAME43733(G43733,G43732,G43731,G43730);
  xor GNAME43743(G43743,G43744,G54130);
  xor GNAME43744(G43744,G54124,G54127);
  and GNAME43745(G43745,G54124,G54130);
  and GNAME43746(G43746,G54127,G54130);
  and GNAME43747(G43747,G54124,G54127);
  or GNAME43748(G43748,G43747,G43746,G43745);
  xor GNAME43758(G43758,G43759,G54139);
  xor GNAME43759(G43759,G54133,G54136);
  and GNAME43760(G43760,G54133,G54139);
  and GNAME43761(G43761,G54136,G54139);
  and GNAME43762(G43762,G54133,G54136);
  or GNAME43763(G43763,G43762,G43761,G43760);
  xor GNAME43773(G43773,G43774,G54148);
  xor GNAME43774(G43774,G54142,G54145);
  and GNAME43775(G43775,G54142,G54148);
  and GNAME43776(G43776,G54145,G54148);
  and GNAME43777(G43777,G54142,G54145);
  or GNAME43778(G43778,G43777,G43776,G43775);
  xor GNAME43788(G43788,G43789,G54157);
  xor GNAME43789(G43789,G54151,G54154);
  and GNAME43790(G43790,G54151,G54157);
  and GNAME43791(G43791,G54154,G54157);
  and GNAME43792(G43792,G54151,G54154);
  or GNAME43793(G43793,G43792,G43791,G43790);
  xor GNAME43803(G43803,G43804,G54166);
  xor GNAME43804(G43804,G54160,G54163);
  and GNAME43805(G43805,G54160,G54166);
  and GNAME43806(G43806,G54163,G54166);
  and GNAME43807(G43807,G54160,G54163);
  or GNAME43808(G43808,G43807,G43806,G43805);
  xor GNAME43818(G43818,G43819,G54175);
  xor GNAME43819(G43819,G54169,G54172);
  and GNAME43820(G43820,G54169,G54175);
  and GNAME43821(G43821,G54172,G54175);
  and GNAME43822(G43822,G54169,G54172);
  or GNAME43823(G43823,G43822,G43821,G43820);
  xor GNAME43833(G43833,G43834,G54184);
  xor GNAME43834(G43834,G54178,G54181);
  and GNAME43835(G43835,G54178,G54184);
  and GNAME43836(G43836,G54181,G54184);
  and GNAME43837(G43837,G54178,G54181);
  or GNAME43838(G43838,G43837,G43836,G43835);
  xor GNAME43848(G43848,G43849,G54193);
  xor GNAME43849(G43849,G54187,G54190);
  and GNAME43850(G43850,G54187,G54193);
  and GNAME43851(G43851,G54190,G54193);
  and GNAME43852(G43852,G54187,G54190);
  or GNAME43853(G43853,G43852,G43851,G43850);
  xor GNAME43863(G43863,G43864,G43823);
  xor GNAME43864(G43864,G51254,G44048);
  and GNAME43865(G43865,G51254,G43823);
  and GNAME43866(G43866,G44048,G43823);
  and GNAME43867(G43867,G51254,G44048);
  or GNAME43868(G43868,G43867,G43866,G43865);
  xor GNAME43878(G43878,G43879,G43838);
  xor GNAME43879(G43879,G51260,G44078);
  and GNAME43880(G43880,G51260,G43838);
  and GNAME43881(G43881,G44078,G43838);
  and GNAME43882(G43882,G51260,G44078);
  or GNAME43883(G43883,G43882,G43881,G43880);
  xor GNAME43893(G43893,G43894,G43853);
  xor GNAME43894(G43894,G51266,G44093);
  and GNAME43895(G43895,G51266,G43853);
  and GNAME43896(G43896,G44093,G43853);
  and GNAME43897(G43897,G51266,G44093);
  or GNAME43898(G43898,G43897,G43896,G43895);
  xor GNAME43908(G43908,G43909,G51236);
  xor GNAME43909(G43909,G54196,G54199);
  and GNAME43910(G43910,G54196,G51236);
  and GNAME43911(G43911,G54199,G51236);
  and GNAME43912(G43912,G54196,G54199);
  or GNAME43913(G43913,G43912,G43911,G43910);
  xor GNAME43923(G43923,G43924,G51242);
  xor GNAME43924(G43924,G54202,G54205);
  and GNAME43925(G43925,G54202,G51242);
  and GNAME43926(G43926,G54205,G51242);
  and GNAME43927(G43927,G54202,G54205);
  or GNAME43928(G43928,G43927,G43926,G43925);
  xor GNAME43938(G43938,G43939,G51248);
  xor GNAME43939(G43939,G54208,G54211);
  and GNAME43940(G43940,G54208,G51248);
  and GNAME43941(G43941,G54211,G51248);
  and GNAME43942(G43942,G54208,G54211);
  or GNAME43943(G43943,G43942,G43941,G43940);
  xor GNAME43953(G43953,G43954,G40718);
  xor GNAME43954(G43954,G54214,G51253);
  and GNAME43955(G43955,G54214,G40718);
  and GNAME43956(G43956,G51253,G40718);
  and GNAME43957(G43957,G54214,G51253);
  or GNAME43958(G43958,G43957,G43956,G43955);
  xor GNAME43968(G43968,G43969,G40733);
  xor GNAME43969(G43969,G54217,G51259);
  and GNAME43970(G43970,G54217,G40733);
  and GNAME43971(G43971,G51259,G40733);
  and GNAME43972(G43972,G54217,G51259);
  or GNAME43973(G43973,G43972,G43971,G43970);
  xor GNAME43983(G43983,G43984,G40748);
  xor GNAME43984(G43984,G54220,G51265);
  and GNAME43985(G43985,G54220,G40748);
  and GNAME43986(G43986,G51265,G40748);
  and GNAME43987(G43987,G54220,G51265);
  or GNAME43988(G43988,G43987,G43986,G43985);
  xor GNAME43998(G43998,G43999,G40713);
  xor GNAME43999(G43999,G44183,G44408);
  and GNAME44000(G44000,G44183,G40713);
  and GNAME44001(G44001,G44408,G40713);
  and GNAME44002(G44002,G44183,G44408);
  or GNAME44003(G44003,G44002,G44001,G44000);
  xor GNAME44013(G44013,G44014,G40728);
  xor GNAME44014(G44014,G44213,G44423);
  and GNAME44015(G44015,G44213,G40728);
  and GNAME44016(G44016,G44423,G40728);
  and GNAME44017(G44017,G44213,G44423);
  or GNAME44018(G44018,G44017,G44016,G44015);
  xor GNAME44028(G44028,G44029,G40743);
  xor GNAME44029(G44029,G44228,G44438);
  and GNAME44030(G44030,G44228,G40743);
  and GNAME44031(G44031,G44438,G40743);
  and GNAME44032(G44032,G44228,G44438);
  or GNAME44033(G44033,G44032,G44031,G44030);
  xor GNAME44043(G44043,G44044,G54226);
  xor GNAME44044(G44044,G54223,G54229);
  and GNAME44045(G44045,G54223,G54226);
  and GNAME44046(G44046,G54229,G54226);
  and GNAME44047(G44047,G54223,G54229);
  or GNAME44048(G44048,G44047,G44046,G44045);
  xor GNAME44058(G44058,G44059,G54238);
  xor GNAME44059(G44059,G54232,G54235);
  and GNAME44060(G44060,G54232,G54238);
  and GNAME44061(G44061,G54235,G54238);
  and GNAME44062(G44062,G54232,G54235);
  or GNAME44063(G44063,G44062,G44061,G44060);
  xor GNAME44073(G44073,G44074,G54244);
  xor GNAME44074(G44074,G54241,G54247);
  and GNAME44075(G44075,G54241,G54244);
  and GNAME44076(G44076,G54247,G54244);
  and GNAME44077(G44077,G54241,G54247);
  or GNAME44078(G44078,G44077,G44076,G44075);
  xor GNAME44088(G44088,G44089,G54253);
  xor GNAME44089(G44089,G54250,G54256);
  and GNAME44090(G44090,G54250,G54253);
  and GNAME44091(G44091,G54256,G54253);
  and GNAME44092(G44092,G54250,G54256);
  or GNAME44093(G44093,G44092,G44091,G44090);
  xor GNAME44103(G44103,G44104,G54265);
  xor GNAME44104(G44104,G54259,G54262);
  and GNAME44105(G44105,G54259,G54265);
  and GNAME44106(G44106,G54262,G54265);
  and GNAME44107(G44107,G54259,G54262);
  or GNAME44108(G44108,G44107,G44106,G44105);
  xor GNAME44118(G44118,G44119,G54274);
  xor GNAME44119(G44119,G54268,G54271);
  and GNAME44120(G44120,G54268,G54274);
  and GNAME44121(G44121,G54271,G54274);
  and GNAME44122(G44122,G54268,G54271);
  or GNAME44123(G44123,G44122,G44121,G44120);
  xor GNAME44133(G44133,G44134,G44333);
  xor GNAME44134(G44134,G40758,G44193);
  and GNAME44135(G44135,G40758,G44333);
  and GNAME44136(G44136,G44193,G44333);
  and GNAME44137(G44137,G40758,G44193);
  or GNAME44138(G44138,G44137,G44136,G44135);
  xor GNAME44148(G44148,G44149,G44378);
  xor GNAME44149(G44149,G40773,G44238);
  and GNAME44150(G44150,G40773,G44378);
  and GNAME44151(G44151,G44238,G44378);
  and GNAME44152(G44152,G40773,G44238);
  or GNAME44153(G44153,G44152,G44151,G44150);
  xor GNAME44163(G44163,G44164,G44393);
  xor GNAME44164(G44164,G40788,G44253);
  and GNAME44165(G44165,G40788,G44393);
  and GNAME44166(G44166,G44253,G44393);
  and GNAME44167(G44167,G40788,G44253);
  or GNAME44168(G44168,G44167,G44166,G44165);
  xor GNAME44178(G44178,G44179,G54283);
  xor GNAME44179(G44179,G54277,G54280);
  and GNAME44180(G44180,G54277,G54283);
  and GNAME44181(G44181,G54280,G54283);
  and GNAME44182(G44182,G54277,G54280);
  or GNAME44183(G44183,G44182,G44181,G44180);
  xor GNAME44193(G44193,G44194,G54292);
  xor GNAME44194(G44194,G54286,G54289);
  and GNAME44195(G44195,G54286,G54292);
  and GNAME44196(G44196,G54289,G54292);
  and GNAME44197(G44197,G54286,G54289);
  or GNAME44198(G44198,G44197,G44196,G44195);
  xor GNAME44208(G44208,G44209,G54301);
  xor GNAME44209(G44209,G54295,G54298);
  and GNAME44210(G44210,G54295,G54301);
  and GNAME44211(G44211,G54298,G54301);
  and GNAME44212(G44212,G54295,G54298);
  or GNAME44213(G44213,G44212,G44211,G44210);
  xor GNAME44223(G44223,G44224,G54310);
  xor GNAME44224(G44224,G54304,G54307);
  and GNAME44225(G44225,G54304,G54310);
  and GNAME44226(G44226,G54307,G54310);
  and GNAME44227(G44227,G54304,G54307);
  or GNAME44228(G44228,G44227,G44226,G44225);
  xor GNAME44238(G44238,G44239,G54319);
  xor GNAME44239(G44239,G54313,G54316);
  and GNAME44240(G44240,G54313,G54319);
  and GNAME44241(G44241,G54316,G54319);
  and GNAME44242(G44242,G54313,G54316);
  or GNAME44243(G44243,G44242,G44241,G44240);
  xor GNAME44253(G44253,G44254,G54328);
  xor GNAME44254(G44254,G54322,G54325);
  and GNAME44255(G44255,G54322,G54328);
  and GNAME44256(G44256,G54325,G54328);
  and GNAME44257(G44257,G54322,G54325);
  or GNAME44258(G44258,G44257,G44256,G44255);
  xor GNAME44268(G44268,G44269,G44198);
  xor GNAME44269(G44269,G51235,G40763);
  and GNAME44270(G44270,G51235,G44198);
  and GNAME44271(G44271,G40763,G44198);
  and GNAME44272(G44272,G51235,G40763);
  or GNAME44273(G44273,G44272,G44271,G44270);
  xor GNAME44283(G44283,G44284,G44243);
  xor GNAME44284(G44284,G51241,G40778);
  and GNAME44285(G44285,G51241,G44243);
  and GNAME44286(G44286,G40778,G44243);
  and GNAME44287(G44287,G51241,G40778);
  or GNAME44288(G44288,G44287,G44286,G44285);
  xor GNAME44298(G44298,G44299,G44258);
  xor GNAME44299(G44299,G51247,G40793);
  and GNAME44300(G44300,G51247,G44258);
  and GNAME44301(G44301,G40793,G44258);
  and GNAME44302(G44302,G51247,G40793);
  or GNAME44303(G44303,G44302,G44301,G44300);
  xor GNAME44313(G44313,G44314,G44453);
  xor GNAME44314(G44314,G54331,G51272);
  and GNAME44315(G44315,G54331,G44453);
  and GNAME44316(G44316,G51272,G44453);
  and GNAME44317(G44317,G54331,G51272);
  or GNAME44318(G44318,G44317,G44316,G44315);
  xor GNAME44328(G44328,G44329,G51271);
  xor GNAME44329(G44329,G54334,G54337);
  and GNAME44330(G44330,G54334,G51271);
  and GNAME44331(G44331,G54337,G51271);
  and GNAME44332(G44332,G54334,G54337);
  or GNAME44333(G44333,G44332,G44331,G44330);
  xor GNAME44343(G44343,G44344,G44468);
  xor GNAME44344(G44344,G54340,G51278);
  and GNAME44345(G44345,G54340,G44468);
  and GNAME44346(G44346,G51278,G44468);
  and GNAME44347(G44347,G54340,G51278);
  or GNAME44348(G44348,G44347,G44346,G44345);
  xor GNAME44358(G44358,G44359,G44483);
  xor GNAME44359(G44359,G54343,G51284);
  and GNAME44360(G44360,G54343,G44483);
  and GNAME44361(G44361,G51284,G44483);
  and GNAME44362(G44362,G54343,G51284);
  or GNAME44363(G44363,G44362,G44361,G44360);
  xor GNAME44373(G44373,G44374,G51277);
  xor GNAME44374(G44374,G54346,G54349);
  and GNAME44375(G44375,G54346,G51277);
  and GNAME44376(G44376,G54349,G51277);
  and GNAME44377(G44377,G54346,G54349);
  or GNAME44378(G44378,G44377,G44376,G44375);
  xor GNAME44388(G44388,G44389,G51283);
  xor GNAME44389(G44389,G54352,G54355);
  and GNAME44390(G44390,G54352,G51283);
  and GNAME44391(G44391,G54355,G51283);
  and GNAME44392(G44392,G54352,G54355);
  or GNAME44393(G44393,G44392,G44391,G44390);
  xor GNAME44403(G44403,G44404,G54361);
  xor GNAME44404(G44404,G54358,G54364);
  and GNAME44405(G44405,G54358,G54361);
  and GNAME44406(G44406,G54364,G54361);
  and GNAME44407(G44407,G54358,G54364);
  or GNAME44408(G44408,G44407,G44406,G44405);
  xor GNAME44418(G44418,G44419,G54370);
  xor GNAME44419(G44419,G54367,G54373);
  and GNAME44420(G44420,G54367,G54370);
  and GNAME44421(G44421,G54373,G54370);
  and GNAME44422(G44422,G54367,G54373);
  or GNAME44423(G44423,G44422,G44421,G44420);
  xor GNAME44433(G44433,G44434,G54379);
  xor GNAME44434(G44434,G54376,G54382);
  and GNAME44435(G44435,G54376,G54379);
  and GNAME44436(G44436,G54382,G54379);
  and GNAME44437(G44437,G54376,G54382);
  or GNAME44438(G44438,G44437,G44436,G44435);
  xor GNAME44448(G44448,G44449,G54388);
  xor GNAME44449(G44449,G54385,G54391);
  and GNAME44450(G44450,G54385,G54388);
  and GNAME44451(G44451,G54391,G54388);
  and GNAME44452(G44452,G54385,G54391);
  or GNAME44453(G44453,G44452,G44451,G44450);
  xor GNAME44463(G44463,G44464,G54397);
  xor GNAME44464(G44464,G54394,G54400);
  and GNAME44465(G44465,G54394,G54397);
  and GNAME44466(G44466,G54400,G54397);
  and GNAME44467(G44467,G54394,G54400);
  or GNAME44468(G44468,G44467,G44466,G44465);
  xor GNAME44478(G44478,G44479,G54406);
  xor GNAME44479(G44479,G54403,G54409);
  and GNAME44480(G44480,G54403,G54406);
  and GNAME44481(G44481,G54409,G54406);
  and GNAME44482(G44482,G54403,G54409);
  or GNAME44483(G44483,G44482,G44481,G44480);
  xor GNAME44493(G44493,G44494,G44448);
  xor GNAME44494(G44494,G40808,G44633);
  and GNAME44495(G44495,G40808,G44448);
  and GNAME44496(G44496,G44633,G44448);
  and GNAME44497(G44497,G40808,G44633);
  or GNAME44498(G44498,G44497,G44496,G44495);
  xor GNAME44508(G44508,G44509,G40803);
  xor GNAME44509(G44509,G51290,G44588);
  and GNAME44510(G44510,G51290,G40803);
  and GNAME44511(G44511,G44588,G40803);
  and GNAME44512(G44512,G51290,G44588);
  or GNAME44513(G44513,G44512,G44511,G44510);
  xor GNAME44523(G44523,G44524,G44463);
  xor GNAME44524(G44524,G40823,G44648);
  and GNAME44525(G44525,G40823,G44463);
  and GNAME44526(G44526,G44648,G44463);
  and GNAME44527(G44527,G40823,G44648);
  or GNAME44528(G44528,G44527,G44526,G44525);
  xor GNAME44538(G44538,G44539,G44478);
  xor GNAME44539(G44539,G40838,G44663);
  and GNAME44540(G44540,G40838,G44478);
  and GNAME44541(G44541,G44663,G44478);
  and GNAME44542(G44542,G40838,G44663);
  or GNAME44543(G44543,G44542,G44541,G44540);
  xor GNAME44553(G44553,G44554,G40818);
  xor GNAME44554(G44554,G51296,G44603);
  and GNAME44555(G44555,G51296,G40818);
  and GNAME44556(G44556,G44603,G40818);
  and GNAME44557(G44557,G51296,G44603);
  or GNAME44558(G44558,G44557,G44556,G44555);
  xor GNAME44568(G44568,G44569,G40833);
  xor GNAME44569(G44569,G51302,G44618);
  and GNAME44570(G44570,G51302,G40833);
  and GNAME44571(G44571,G44618,G40833);
  and GNAME44572(G44572,G51302,G44618);
  or GNAME44573(G44573,G44572,G44571,G44570);
  xor GNAME44583(G44583,G44584,G54415);
  xor GNAME44584(G44584,G54412,G54418);
  and GNAME44585(G44585,G54412,G54415);
  and GNAME44586(G44586,G54418,G54415);
  and GNAME44587(G44587,G54412,G54418);
  or GNAME44588(G44588,G44587,G44586,G44585);
  xor GNAME44598(G44598,G44599,G54424);
  xor GNAME44599(G44599,G54421,G54427);
  and GNAME44600(G44600,G54421,G54424);
  and GNAME44601(G44601,G54427,G54424);
  and GNAME44602(G44602,G54421,G54427);
  or GNAME44603(G44603,G44602,G44601,G44600);
  xor GNAME44613(G44613,G44614,G54433);
  xor GNAME44614(G44614,G54430,G54436);
  and GNAME44615(G44615,G54430,G54433);
  and GNAME44616(G44616,G54436,G54433);
  and GNAME44617(G44617,G54430,G54436);
  or GNAME44618(G44618,G44617,G44616,G44615);
  xor GNAME44628(G44628,G44629,G54445);
  xor GNAME44629(G44629,G54439,G54442);
  and GNAME44630(G44630,G54439,G54445);
  and GNAME44631(G44631,G54442,G54445);
  and GNAME44632(G44632,G54439,G54442);
  or GNAME44633(G44633,G44632,G44631,G44630);
  xor GNAME44643(G44643,G44644,G54454);
  xor GNAME44644(G44644,G54448,G54451);
  and GNAME44645(G44645,G54448,G54454);
  and GNAME44646(G44646,G54451,G54454);
  and GNAME44647(G44647,G54448,G54451);
  or GNAME44648(G44648,G44647,G44646,G44645);
  xor GNAME44658(G44658,G44659,G54463);
  xor GNAME44659(G44659,G54457,G54460);
  and GNAME44660(G44660,G54457,G54463);
  and GNAME44661(G44661,G54460,G54463);
  and GNAME44662(G44662,G54457,G54460);
  or GNAME44663(G44663,G44662,G44661,G44660);
  xor GNAME44673(G44673,G44674,G54469);
  xor GNAME44674(G44674,G54466,G54472);
  and GNAME44675(G44675,G54466,G54469);
  and GNAME44676(G44676,G54472,G54469);
  and GNAME44677(G44677,G54466,G54472);
  or GNAME44678(G44678,G44677,G44676,G44675);
  xor GNAME44688(G44688,G44689,G54478);
  xor GNAME44689(G44689,G54475,G54481);
  and GNAME44690(G44690,G54475,G54478);
  and GNAME44691(G44691,G54481,G54478);
  and GNAME44692(G44692,G54475,G54481);
  or GNAME44693(G44693,G44692,G44691,G44690);
  xor GNAME44703(G44703,G44704,G54487);
  xor GNAME44704(G44704,G54484,G54490);
  and GNAME44705(G44705,G54484,G54487);
  and GNAME44706(G44706,G54490,G54487);
  and GNAME44707(G44707,G54484,G54490);
  or GNAME44708(G44708,G44707,G44706,G44705);
  xor GNAME44718(G44718,G44719,G51308);
  xor GNAME44719(G44719,G54493,G54496);
  and GNAME44720(G44720,G54493,G51308);
  and GNAME44721(G44721,G54496,G51308);
  and GNAME44722(G44722,G54493,G54496);
  or GNAME44723(G44723,G44722,G44721,G44720);
  xor GNAME44733(G44733,G44734,G51314);
  xor GNAME44734(G44734,G54499,G54502);
  and GNAME44735(G44735,G54499,G51314);
  and GNAME44736(G44736,G54502,G51314);
  and GNAME44737(G44737,G54499,G54502);
  or GNAME44738(G44738,G44737,G44736,G44735);
  xor GNAME44748(G44748,G44749,G51320);
  xor GNAME44749(G44749,G54505,G54508);
  and GNAME44750(G44750,G54505,G51320);
  and GNAME44751(G44751,G54508,G51320);
  and GNAME44752(G44752,G54505,G54508);
  or GNAME44753(G44753,G44752,G44751,G44750);
  xor GNAME44763(G44763,G44764,G40853);
  xor GNAME44764(G44764,G54511,G51289);
  and GNAME44765(G44765,G54511,G40853);
  and GNAME44766(G44766,G51289,G40853);
  and GNAME44767(G44767,G54511,G51289);
  or GNAME44768(G44768,G44767,G44766,G44765);
  xor GNAME44778(G44778,G44779,G40868);
  xor GNAME44779(G44779,G54514,G51295);
  and GNAME44780(G44780,G54514,G40868);
  and GNAME44781(G44781,G51295,G40868);
  and GNAME44782(G44782,G54514,G51295);
  or GNAME44783(G44783,G44782,G44781,G44780);
  xor GNAME44793(G44793,G44794,G40883);
  xor GNAME44794(G44794,G54517,G51301);
  and GNAME44795(G44795,G54517,G40883);
  and GNAME44796(G44796,G51301,G40883);
  and GNAME44797(G44797,G54517,G51301);
  or GNAME44798(G44798,G44797,G44796,G44795);
  xor GNAME44808(G44808,G44809,G44673);
  xor GNAME44809(G44809,G51307,G40898);
  and GNAME44810(G44810,G51307,G44673);
  and GNAME44811(G44811,G40898,G44673);
  and GNAME44812(G44812,G51307,G40898);
  or GNAME44813(G44813,G44812,G44811,G44810);
  xor GNAME44823(G44823,G44824,G44718);
  xor GNAME44824(G44824,G44678,G40848);
  and GNAME44825(G44825,G44678,G44718);
  and GNAME44826(G44826,G40848,G44718);
  and GNAME44827(G44827,G44678,G40848);
  or GNAME44828(G44828,G44827,G44826,G44825);
  xor GNAME44838(G44838,G44839,G44733);
  xor GNAME44839(G44839,G44693,G40863);
  and GNAME44840(G44840,G44693,G44733);
  and GNAME44841(G44841,G40863,G44733);
  and GNAME44842(G44842,G44693,G40863);
  or GNAME44843(G44843,G44842,G44841,G44840);
  xor GNAME44853(G44853,G44854,G44748);
  xor GNAME44854(G44854,G44708,G40878);
  and GNAME44855(G44855,G44708,G44748);
  and GNAME44856(G44856,G40878,G44748);
  and GNAME44857(G44857,G44708,G40878);
  or GNAME44858(G44858,G44857,G44856,G44855);
  xor GNAME44868(G44868,G44869,G44688);
  xor GNAME44869(G44869,G51313,G40913);
  and GNAME44870(G44870,G51313,G44688);
  and GNAME44871(G44871,G40913,G44688);
  and GNAME44872(G44872,G51313,G40913);
  or GNAME44873(G44873,G44872,G44871,G44870);
  xor GNAME44883(G44883,G44884,G44703);
  xor GNAME44884(G44884,G51319,G40928);
  and GNAME44885(G44885,G51319,G44703);
  and GNAME44886(G44886,G40928,G44703);
  and GNAME44887(G44887,G51319,G40928);
  or GNAME44888(G44888,G44887,G44886,G44885);
  xor GNAME44898(G44898,G44899,G40893);
  xor GNAME44899(G44899,G54520,G51344);
  and GNAME44900(G44900,G54520,G40893);
  and GNAME44901(G44901,G51344,G40893);
  and GNAME44902(G44902,G54520,G51344);
  or GNAME44903(G44903,G44902,G44901,G44900);
  xor GNAME44913(G44913,G44914,G52006);
  xor GNAME44914(G44914,G44903,G44808);
  and GNAME44915(G44915,G44903,G52006);
  and GNAME44916(G44916,G44808,G52006);
  and GNAME44917(G44917,G44903,G44808);
  or GNAME44918(G44918,G44917,G44916,G44915);
  xor GNAME44928(G44928,G44929,G40908);
  xor GNAME44929(G44929,G54523,G51350);
  and GNAME44930(G44930,G54523,G40908);
  and GNAME44931(G44931,G51350,G40908);
  and GNAME44932(G44932,G54523,G51350);
  or GNAME44933(G44933,G44932,G44931,G44930);
  xor GNAME44943(G44943,G44944,G52026);
  xor GNAME44944(G44944,G44933,G44868);
  and GNAME44945(G44945,G44933,G52026);
  and GNAME44946(G44946,G44868,G52026);
  and GNAME44947(G44947,G44933,G44868);
  or GNAME44948(G44948,G44947,G44946,G44945);
  xor GNAME44958(G44958,G44959,G40923);
  xor GNAME44959(G44959,G54526,G51356);
  and GNAME44960(G44960,G54526,G40923);
  and GNAME44961(G44961,G51356,G40923);
  and GNAME44962(G44962,G54526,G51356);
  or GNAME44963(G44963,G44962,G44961,G44960);
  xor GNAME44973(G44973,G44974,G52046);
  xor GNAME44974(G44974,G44963,G44883);
  and GNAME44975(G44975,G44963,G52046);
  and GNAME44976(G44976,G44883,G52046);
  and GNAME44977(G44977,G44963,G44883);
  or GNAME44978(G44978,G44977,G44976,G44975);
  xor GNAME44988(G44988,G44989,G41438);
  xor GNAME44989(G44989,G41343,G41298);
  and GNAME44990(G44990,G41343,G41438);
  and GNAME44991(G44991,G41298,G41438);
  and GNAME44992(G44992,G41343,G41298);
  or GNAME44993(G44993,G44992,G44991,G44990);
  xor GNAME45003(G45003,G45004,G41453);
  xor GNAME45004(G45004,G41358,G41313);
  and GNAME45005(G45005,G41358,G41453);
  and GNAME45006(G45006,G41313,G41453);
  and GNAME45007(G45007,G41358,G41313);
  or GNAME45008(G45008,G45007,G45006,G45005);
  xor GNAME45018(G45018,G45019,G41468);
  xor GNAME45019(G45019,G41373,G41328);
  and GNAME45020(G45020,G41373,G41468);
  and GNAME45021(G45021,G41328,G41468);
  and GNAME45022(G45022,G41373,G41328);
  or GNAME45023(G45023,G45022,G45021,G45020);
  xor GNAME45033(G45033,G45034,G45083);
  xor GNAME45034(G45034,G41528,G41433);
  and GNAME45035(G45035,G41528,G45083);
  and GNAME45036(G45036,G41433,G45083);
  and GNAME45037(G45037,G41528,G41433);
  or GNAME45038(G45038,G45037,G45036,G45035);
  xor GNAME45048(G45048,G45049,G45098);
  xor GNAME45049(G45049,G41543,G41448);
  and GNAME45050(G45050,G41543,G45098);
  and GNAME45051(G45051,G41448,G45098);
  and GNAME45052(G45052,G41543,G41448);
  or GNAME45053(G45053,G45052,G45051,G45050);
  xor GNAME45063(G45063,G45064,G45113);
  xor GNAME45064(G45064,G41558,G41463);
  and GNAME45065(G45065,G41558,G45113);
  and GNAME45066(G45066,G41463,G45113);
  and GNAME45067(G45067,G41558,G41463);
  or GNAME45068(G45068,G45067,G45066,G45065);
  xor GNAME45078(G45078,G45079,G41708);
  xor GNAME45079(G45079,G41798,G41478);
  and GNAME45080(G45080,G41798,G41708);
  and GNAME45081(G45081,G41478,G41708);
  and GNAME45082(G45082,G41798,G41478);
  or GNAME45083(G45083,G45082,G45081,G45080);
  xor GNAME45093(G45093,G45094,G41723);
  xor GNAME45094(G45094,G41813,G41493);
  and GNAME45095(G45095,G41813,G41723);
  and GNAME45096(G45096,G41493,G41723);
  and GNAME45097(G45097,G41813,G41493);
  or GNAME45098(G45098,G45097,G45096,G45095);
  xor GNAME45108(G45108,G45109,G41738);
  xor GNAME45109(G45109,G41828,G41508);
  and GNAME45110(G45110,G41828,G41738);
  and GNAME45111(G45111,G41508,G41738);
  and GNAME45112(G45112,G41828,G41508);
  or GNAME45113(G45113,G45112,G45111,G45110);
  xor GNAME45123(G45123,G45124,G45078);
  xor GNAME45124(G45124,G41523,G41573);
  and GNAME45125(G45125,G41523,G45078);
  and GNAME45126(G45126,G41573,G45078);
  and GNAME45127(G45127,G41523,G41573);
  or GNAME45128(G45128,G45127,G45126,G45125);
  xor GNAME45138(G45138,G45139,G41568);
  xor GNAME45139(G45139,G41703,G45218);
  and GNAME45140(G45140,G41703,G41568);
  and GNAME45141(G45141,G45218,G41568);
  and GNAME45142(G45142,G41703,G45218);
  or GNAME45143(G45143,G45142,G45141,G45140);
  xor GNAME45153(G45153,G45154,G45093);
  xor GNAME45154(G45154,G41538,G41588);
  and GNAME45155(G45155,G41538,G45093);
  and GNAME45156(G45156,G41588,G45093);
  and GNAME45157(G45157,G41538,G41588);
  or GNAME45158(G45158,G45157,G45156,G45155);
  xor GNAME45168(G45168,G45169,G45108);
  xor GNAME45169(G45169,G41553,G41603);
  and GNAME45170(G45170,G41553,G45108);
  and GNAME45171(G45171,G41603,G45108);
  and GNAME45172(G45172,G41553,G41603);
  or GNAME45173(G45173,G45172,G45171,G45170);
  xor GNAME45183(G45183,G45184,G41583);
  xor GNAME45184(G45184,G41718,G45248);
  and GNAME45185(G45185,G41718,G41583);
  and GNAME45186(G45186,G45248,G41583);
  and GNAME45187(G45187,G41718,G45248);
  or GNAME45188(G45188,G45187,G45186,G45185);
  xor GNAME45198(G45198,G45199,G41598);
  xor GNAME45199(G45199,G41733,G45278);
  and GNAME45200(G45200,G41733,G41598);
  and GNAME45201(G45201,G45278,G41598);
  and GNAME45202(G45202,G41733,G45278);
  or GNAME45203(G45203,G45202,G45201,G45200);
  xor GNAME45213(G45213,G45214,G41978);
  xor GNAME45214(G45214,G41748,G41888);
  and GNAME45215(G45215,G41748,G41978);
  and GNAME45216(G45216,G41888,G41978);
  and GNAME45217(G45217,G41748,G41888);
  or GNAME45218(G45218,G45217,G45216,G45215);
  xor GNAME45228(G45228,G45229,G45398);
  xor GNAME45229(G45229,G42113,G41883);
  and GNAME45230(G45230,G42113,G45398);
  and GNAME45231(G45231,G41883,G45398);
  and GNAME45232(G45232,G42113,G41883);
  or GNAME45233(G45233,G45232,G45231,G45230);
  xor GNAME45243(G45243,G45244,G41993);
  xor GNAME45244(G45244,G41763,G41903);
  and GNAME45245(G45245,G41763,G41993);
  and GNAME45246(G45246,G41903,G41993);
  and GNAME45247(G45247,G41763,G41903);
  or GNAME45248(G45248,G45247,G45246,G45245);
  xor GNAME45258(G45258,G45259,G45413);
  xor GNAME45259(G45259,G42143,G41898);
  and GNAME45260(G45260,G42143,G45413);
  and GNAME45261(G45261,G41898,G45413);
  and GNAME45262(G45262,G42143,G41898);
  or GNAME45263(G45263,G45262,G45261,G45260);
  xor GNAME45273(G45273,G45274,G42008);
  xor GNAME45274(G45274,G41778,G41918);
  and GNAME45275(G45275,G41778,G42008);
  and GNAME45276(G45276,G41918,G42008);
  and GNAME45277(G45277,G41778,G41918);
  or GNAME45278(G45278,G45277,G45276,G45275);
  xor GNAME45288(G45288,G45289,G45428);
  xor GNAME45289(G45289,G42158,G41913);
  and GNAME45290(G45290,G42158,G45428);
  and GNAME45291(G45291,G41913,G45428);
  and GNAME45292(G45292,G42158,G41913);
  or GNAME45293(G45293,G45292,G45291,G45290);
  xor GNAME45303(G45303,G45304,G45213);
  xor GNAME45304(G45304,G41658,G45233);
  and GNAME45305(G45305,G41658,G45213);
  and GNAME45306(G45306,G45233,G45213);
  and GNAME45307(G45307,G41658,G45233);
  or GNAME45308(G45308,G45307,G45306,G45305);
  xor GNAME45318(G45318,G45319,G45228);
  xor GNAME45319(G45319,G41973,G45443);
  and GNAME45320(G45320,G41973,G45228);
  and GNAME45321(G45321,G45443,G45228);
  and GNAME45322(G45322,G41973,G45443);
  or GNAME45323(G45323,G45322,G45321,G45320);
  xor GNAME45333(G45333,G45334,G45243);
  xor GNAME45334(G45334,G41673,G45263);
  and GNAME45335(G45335,G41673,G45243);
  and GNAME45336(G45336,G45263,G45243);
  and GNAME45337(G45337,G41673,G45263);
  or GNAME45338(G45338,G45337,G45336,G45335);
  xor GNAME45348(G45348,G45349,G45273);
  xor GNAME45349(G45349,G41688,G45293);
  and GNAME45350(G45350,G41688,G45273);
  and GNAME45351(G45351,G45293,G45273);
  and GNAME45352(G45352,G41688,G45293);
  or GNAME45353(G45353,G45352,G45351,G45350);
  xor GNAME45363(G45363,G45364,G45258);
  xor GNAME45364(G45364,G41988,G45473);
  and GNAME45365(G45365,G41988,G45258);
  and GNAME45366(G45366,G45473,G45258);
  and GNAME45367(G45367,G41988,G45473);
  or GNAME45368(G45368,G45367,G45366,G45365);
  xor GNAME45378(G45378,G45379,G45288);
  xor GNAME45379(G45379,G42003,G45503);
  and GNAME45380(G45380,G42003,G45288);
  and GNAME45381(G45381,G45503,G45288);
  and GNAME45382(G45382,G42003,G45503);
  or GNAME45383(G45383,G45382,G45381,G45380);
  xor GNAME45393(G45393,G45394,G42018);
  xor GNAME45394(G45394,G42203,G41928);
  and GNAME45395(G45395,G42203,G42018);
  and GNAME45396(G45396,G41928,G42018);
  and GNAME45397(G45397,G42203,G41928);
  or GNAME45398(G45398,G45397,G45396,G45395);
  xor GNAME45408(G45408,G45409,G42033);
  xor GNAME45409(G45409,G42233,G41943);
  and GNAME45410(G45410,G42233,G42033);
  and GNAME45411(G45411,G41943,G42033);
  and GNAME45412(G45412,G42233,G41943);
  or GNAME45413(G45413,G45412,G45411,G45410);
  xor GNAME45423(G45423,G45424,G42048);
  xor GNAME45424(G45424,G42248,G41958);
  and GNAME45425(G45425,G42248,G42048);
  and GNAME45426(G45426,G41958,G42048);
  and GNAME45427(G45427,G42248,G41958);
  or GNAME45428(G45428,G45427,G45426,G45425);
  xor GNAME45438(G45438,G45439,G42293);
  xor GNAME45439(G45439,G42128,G42108);
  and GNAME45440(G45440,G42128,G42293);
  and GNAME45441(G45441,G42108,G42293);
  and GNAME45442(G45442,G42128,G42108);
  or GNAME45443(G45443,G45442,G45441,G45440);
  xor GNAME45453(G45453,G45454,G42308);
  xor GNAME45454(G45454,G45578,G42123);
  and GNAME45455(G45455,G45578,G42308);
  and GNAME45456(G45456,G42123,G42308);
  and GNAME45457(G45457,G45578,G42123);
  or GNAME45458(G45458,G45457,G45456,G45455);
  xor GNAME45468(G45468,G45469,G42323);
  xor GNAME45469(G45469,G42173,G42138);
  and GNAME45470(G45470,G42173,G42323);
  and GNAME45471(G45471,G42138,G42323);
  and GNAME45472(G45472,G42173,G42138);
  or GNAME45473(G45473,G45472,G45471,G45470);
  xor GNAME45483(G45483,G45484,G42338);
  xor GNAME45484(G45484,G45593,G42168);
  and GNAME45485(G45485,G45593,G42338);
  and GNAME45486(G45486,G42168,G42338);
  and GNAME45487(G45487,G45593,G42168);
  or GNAME45488(G45488,G45487,G45486,G45485);
  xor GNAME45498(G45498,G45499,G42353);
  xor GNAME45499(G45499,G42188,G42153);
  and GNAME45500(G45500,G42188,G42353);
  and GNAME45501(G45501,G42153,G42353);
  and GNAME45502(G45502,G42188,G42153);
  or GNAME45503(G45503,G45502,G45501,G45500);
  xor GNAME45513(G45513,G45514,G42368);
  xor GNAME45514(G45514,G45608,G42183);
  and GNAME45515(G45515,G45608,G42368);
  and GNAME45516(G45516,G42183,G42368);
  and GNAME45517(G45517,G45608,G42183);
  or GNAME45518(G45518,G45517,G45516,G45515);
  xor GNAME45528(G45528,G45529,G45453);
  xor GNAME45529(G45529,G42288,G47378);
  and GNAME45530(G45530,G42288,G45453);
  and GNAME45531(G45531,G47378,G45453);
  and GNAME45532(G45532,G42288,G47378);
  or GNAME45533(G45533,G45532,G45531,G45530);
  xor GNAME45543(G45543,G45544,G45483);
  xor GNAME45544(G45544,G42318,G47408);
  and GNAME45545(G45545,G42318,G45483);
  and GNAME45546(G45546,G47408,G45483);
  and GNAME45547(G45547,G42318,G47408);
  or GNAME45548(G45548,G45547,G45546,G45545);
  xor GNAME45558(G45558,G45559,G45513);
  xor GNAME45559(G45559,G42348,G47438);
  and GNAME45560(G45560,G42348,G45513);
  and GNAME45561(G45561,G47438,G45513);
  and GNAME45562(G45562,G42348,G47438);
  or GNAME45563(G45563,G45562,G45561,G45560);
  xor GNAME45573(G45573,G45574,G42428);
  xor GNAME45574(G45574,G42563,G42608);
  and GNAME45575(G45575,G42563,G42428);
  and GNAME45576(G45576,G42608,G42428);
  and GNAME45577(G45577,G42563,G42608);
  or GNAME45578(G45578,G45577,G45576,G45575);
  xor GNAME45588(G45588,G45589,G42443);
  xor GNAME45589(G45589,G42578,G42638);
  and GNAME45590(G45590,G42578,G42443);
  and GNAME45591(G45591,G42638,G42443);
  and GNAME45592(G45592,G42578,G42638);
  or GNAME45593(G45593,G45592,G45591,G45590);
  xor GNAME45603(G45603,G45604,G42458);
  xor GNAME45604(G45604,G42593,G42653);
  and GNAME45605(G45605,G42593,G42458);
  and GNAME45606(G45606,G42653,G42458);
  and GNAME45607(G45607,G42593,G42653);
  or GNAME45608(G45608,G45607,G45606,G45605);
  xor GNAME45618(G45618,G45619,G47373);
  xor GNAME45619(G45619,G42303,G47393);
  and GNAME45620(G45620,G42303,G47373);
  and GNAME45621(G45621,G47393,G47373);
  and GNAME45622(G45622,G42303,G47393);
  or GNAME45623(G45623,G45622,G45621,G45620);
  xor GNAME45633(G45633,G45634,G47403);
  xor GNAME45634(G45634,G42333,G47423);
  and GNAME45635(G45635,G42333,G47403);
  and GNAME45636(G45636,G47423,G47403);
  and GNAME45637(G45637,G42333,G47423);
  or GNAME45638(G45638,G45637,G45636,G45635);
  xor GNAME45648(G45648,G45649,G47433);
  xor GNAME45649(G45649,G42363,G47453);
  and GNAME45650(G45650,G42363,G47433);
  and GNAME45651(G45651,G47453,G47433);
  and GNAME45652(G45652,G42363,G47453);
  or GNAME45653(G45653,G45652,G45651,G45650);
  xor GNAME45663(G45663,G45664,G42473);
  xor GNAME45664(G45664,G42518,G42623);
  and GNAME45665(G45665,G42518,G42473);
  and GNAME45666(G45666,G42623,G42473);
  and GNAME45667(G45667,G42518,G42623);
  or GNAME45668(G45668,G45667,G45666,G45665);
  xor GNAME45678(G45678,G45679,G42488);
  xor GNAME45679(G45679,G42533,G42668);
  and GNAME45680(G45680,G42533,G42488);
  and GNAME45681(G45681,G42668,G42488);
  and GNAME45682(G45682,G42533,G42668);
  or GNAME45683(G45683,G45682,G45681,G45680);
  xor GNAME45693(G45693,G45694,G42503);
  xor GNAME45694(G45694,G42548,G42683);
  and GNAME45695(G45695,G42548,G42503);
  and GNAME45696(G45696,G42683,G42503);
  and GNAME45697(G45697,G42548,G42683);
  or GNAME45698(G45698,G45697,G45696,G45695);
  xor GNAME45708(G45708,G45709,G42603);
  xor GNAME45709(G45709,G42558,G42423);
  and GNAME45710(G45710,G42558,G42603);
  and GNAME45711(G45711,G42423,G42603);
  and GNAME45712(G45712,G42558,G42423);
  or GNAME45713(G45713,G45712,G45711,G45710);
  xor GNAME45723(G45723,G45724,G42618);
  xor GNAME45724(G45724,G42513,G42468);
  and GNAME45725(G45725,G42513,G42618);
  and GNAME45726(G45726,G42468,G42618);
  and GNAME45727(G45727,G42513,G42468);
  or GNAME45728(G45728,G45727,G45726,G45725);
  xor GNAME45738(G45738,G45739,G42633);
  xor GNAME45739(G45739,G42573,G42438);
  and GNAME45740(G45740,G42573,G42633);
  and GNAME45741(G45741,G42438,G42633);
  and GNAME45742(G45742,G42573,G42438);
  or GNAME45743(G45743,G45742,G45741,G45740);
  xor GNAME45753(G45753,G45754,G42663);
  xor GNAME45754(G45754,G42528,G42483);
  and GNAME45755(G45755,G42528,G42663);
  and GNAME45756(G45756,G42483,G42663);
  and GNAME45757(G45757,G42528,G42483);
  or GNAME45758(G45758,G45757,G45756,G45755);
  xor GNAME45768(G45768,G45769,G42648);
  xor GNAME45769(G45769,G42588,G42453);
  and GNAME45770(G45770,G42588,G42648);
  and GNAME45771(G45771,G42453,G42648);
  and GNAME45772(G45772,G42588,G42453);
  or GNAME45773(G45773,G45772,G45771,G45770);
  xor GNAME45783(G45783,G45784,G42678);
  xor GNAME45784(G45784,G42543,G42498);
  and GNAME45785(G45785,G42543,G42678);
  and GNAME45786(G45786,G42498,G42678);
  and GNAME45787(G45787,G42543,G42498);
  or GNAME45788(G45788,G45787,G45786,G45785);
  xor GNAME45798(G45798,G45799,G42698);
  xor GNAME45799(G45799,G42788,G42878);
  and GNAME45800(G45800,G42788,G42698);
  and GNAME45801(G45801,G42878,G42698);
  and GNAME45802(G45802,G42788,G42878);
  or GNAME45803(G45803,G45802,G45801,G45800);
  xor GNAME45813(G45813,G45814,G42713);
  xor GNAME45814(G45814,G42803,G42893);
  and GNAME45815(G45815,G42803,G42713);
  and GNAME45816(G45816,G42893,G42713);
  and GNAME45817(G45817,G42803,G42893);
  or GNAME45818(G45818,G45817,G45816,G45815);
  xor GNAME45828(G45828,G45829,G42728);
  xor GNAME45829(G45829,G42818,G42908);
  and GNAME45830(G45830,G42818,G42728);
  and GNAME45831(G45831,G42908,G42728);
  and GNAME45832(G45832,G42818,G42908);
  or GNAME45833(G45833,G45832,G45831,G45830);
  xor GNAME45843(G45843,G45844,G42743);
  xor GNAME45844(G45844,G42833,G42923);
  and GNAME45845(G45845,G42833,G42743);
  and GNAME45846(G45846,G42923,G42743);
  and GNAME45847(G45847,G42833,G42923);
  or GNAME45848(G45848,G45847,G45846,G45845);
  xor GNAME45858(G45858,G45859,G42758);
  xor GNAME45859(G45859,G42848,G42938);
  and GNAME45860(G45860,G42848,G42758);
  and GNAME45861(G45861,G42938,G42758);
  and GNAME45862(G45862,G42848,G42938);
  or GNAME45863(G45863,G45862,G45861,G45860);
  xor GNAME45873(G45873,G45874,G42773);
  xor GNAME45874(G45874,G42863,G42953);
  and GNAME45875(G45875,G42863,G42773);
  and GNAME45876(G45876,G42953,G42773);
  and GNAME45877(G45877,G42863,G42953);
  or GNAME45878(G45878,G45877,G45876,G45875);
  xor GNAME45888(G45888,G45889,G42873);
  xor GNAME45889(G45889,G42783,G42693);
  and GNAME45890(G45890,G42783,G42873);
  and GNAME45891(G45891,G42693,G42873);
  and GNAME45892(G45892,G42783,G42693);
  or GNAME45893(G45893,G45892,G45891,G45890);
  xor GNAME45903(G45903,G45904,G42888);
  xor GNAME45904(G45904,G42798,G42708);
  and GNAME45905(G45905,G42798,G42888);
  and GNAME45906(G45906,G42708,G42888);
  and GNAME45907(G45907,G42798,G42708);
  or GNAME45908(G45908,G45907,G45906,G45905);
  xor GNAME45918(G45918,G45919,G42903);
  xor GNAME45919(G45919,G42813,G42723);
  and GNAME45920(G45920,G42813,G42903);
  and GNAME45921(G45921,G42723,G42903);
  and GNAME45922(G45922,G42813,G42723);
  or GNAME45923(G45923,G45922,G45921,G45920);
  xor GNAME45933(G45933,G45934,G42933);
  xor GNAME45934(G45934,G42843,G42753);
  and GNAME45935(G45935,G42843,G42933);
  and GNAME45936(G45936,G42753,G42933);
  and GNAME45937(G45937,G42843,G42753);
  or GNAME45938(G45938,G45937,G45936,G45935);
  xor GNAME45948(G45948,G45949,G42918);
  xor GNAME45949(G45949,G42828,G42738);
  and GNAME45950(G45950,G42828,G42918);
  and GNAME45951(G45951,G42738,G42918);
  and GNAME45952(G45952,G42828,G42738);
  or GNAME45953(G45953,G45952,G45951,G45950);
  xor GNAME45963(G45963,G45964,G42948);
  xor GNAME45964(G45964,G42858,G42768);
  and GNAME45965(G45965,G42858,G42948);
  and GNAME45966(G45966,G42768,G42948);
  and GNAME45967(G45967,G42858,G42768);
  or GNAME45968(G45968,G45967,G45966,G45965);
  xor GNAME45978(G45978,G45979,G42968);
  xor GNAME45979(G45979,G43058,G43148);
  and GNAME45980(G45980,G43058,G42968);
  and GNAME45981(G45981,G43148,G42968);
  and GNAME45982(G45982,G43058,G43148);
  or GNAME45983(G45983,G45982,G45981,G45980);
  xor GNAME45993(G45993,G45994,G42983);
  xor GNAME45994(G45994,G43073,G43163);
  and GNAME45995(G45995,G43073,G42983);
  and GNAME45996(G45996,G43163,G42983);
  and GNAME45997(G45997,G43073,G43163);
  or GNAME45998(G45998,G45997,G45996,G45995);
  xor GNAME46008(G46008,G46009,G42998);
  xor GNAME46009(G46009,G43088,G43178);
  and GNAME46010(G46010,G43088,G42998);
  and GNAME46011(G46011,G43178,G42998);
  and GNAME46012(G46012,G43088,G43178);
  or GNAME46013(G46013,G46012,G46011,G46010);
  xor GNAME46023(G46023,G46024,G43013);
  xor GNAME46024(G46024,G43103,G43193);
  and GNAME46025(G46025,G43103,G43013);
  and GNAME46026(G46026,G43193,G43013);
  and GNAME46027(G46027,G43103,G43193);
  or GNAME46028(G46028,G46027,G46026,G46025);
  xor GNAME46038(G46038,G46039,G43028);
  xor GNAME46039(G46039,G43118,G43208);
  and GNAME46040(G46040,G43118,G43028);
  and GNAME46041(G46041,G43208,G43028);
  and GNAME46042(G46042,G43118,G43208);
  or GNAME46043(G46043,G46042,G46041,G46040);
  xor GNAME46053(G46053,G46054,G43043);
  xor GNAME46054(G46054,G43133,G43223);
  and GNAME46055(G46055,G43133,G43043);
  and GNAME46056(G46056,G43223,G43043);
  and GNAME46057(G46057,G43133,G43223);
  or GNAME46058(G46058,G46057,G46056,G46055);
  xor GNAME46068(G46068,G46069,G43143);
  xor GNAME46069(G46069,G43053,G42963);
  and GNAME46070(G46070,G43053,G43143);
  and GNAME46071(G46071,G42963,G43143);
  and GNAME46072(G46072,G43053,G42963);
  or GNAME46073(G46073,G46072,G46071,G46070);
  xor GNAME46083(G46083,G46084,G43158);
  xor GNAME46084(G46084,G43068,G42978);
  and GNAME46085(G46085,G43068,G43158);
  and GNAME46086(G46086,G42978,G43158);
  and GNAME46087(G46087,G43068,G42978);
  or GNAME46088(G46088,G46087,G46086,G46085);
  xor GNAME46098(G46098,G46099,G43173);
  xor GNAME46099(G46099,G43083,G42993);
  and GNAME46100(G46100,G43083,G43173);
  and GNAME46101(G46101,G42993,G43173);
  and GNAME46102(G46102,G43083,G42993);
  or GNAME46103(G46103,G46102,G46101,G46100);
  xor GNAME46113(G46113,G46114,G43203);
  xor GNAME46114(G46114,G43113,G43023);
  and GNAME46115(G46115,G43113,G43203);
  and GNAME46116(G46116,G43023,G43203);
  and GNAME46117(G46117,G43113,G43023);
  or GNAME46118(G46118,G46117,G46116,G46115);
  xor GNAME46128(G46128,G46129,G43188);
  xor GNAME46129(G46129,G43098,G43008);
  and GNAME46130(G46130,G43098,G43188);
  and GNAME46131(G46131,G43008,G43188);
  and GNAME46132(G46132,G43098,G43008);
  or GNAME46133(G46133,G46132,G46131,G46130);
  xor GNAME46143(G46143,G46144,G43218);
  xor GNAME46144(G46144,G43128,G43038);
  and GNAME46145(G46145,G43128,G43218);
  and GNAME46146(G46146,G43038,G43218);
  and GNAME46147(G46147,G43128,G43038);
  or GNAME46148(G46148,G46147,G46146,G46145);
  xor GNAME46158(G46158,G46159,G43238);
  xor GNAME46159(G46159,G43328,G43418);
  and GNAME46160(G46160,G43328,G43238);
  and GNAME46161(G46161,G43418,G43238);
  and GNAME46162(G46162,G43328,G43418);
  or GNAME46163(G46163,G46162,G46161,G46160);
  xor GNAME46173(G46173,G46174,G43253);
  xor GNAME46174(G46174,G43343,G43433);
  and GNAME46175(G46175,G43343,G43253);
  and GNAME46176(G46176,G43433,G43253);
  and GNAME46177(G46177,G43343,G43433);
  or GNAME46178(G46178,G46177,G46176,G46175);
  xor GNAME46188(G46188,G46189,G43268);
  xor GNAME46189(G46189,G43358,G43448);
  and GNAME46190(G46190,G43358,G43268);
  and GNAME46191(G46191,G43448,G43268);
  and GNAME46192(G46192,G43358,G43448);
  or GNAME46193(G46193,G46192,G46191,G46190);
  xor GNAME46203(G46203,G46204,G43283);
  xor GNAME46204(G46204,G43373,G43463);
  and GNAME46205(G46205,G43373,G43283);
  and GNAME46206(G46206,G43463,G43283);
  and GNAME46207(G46207,G43373,G43463);
  or GNAME46208(G46208,G46207,G46206,G46205);
  xor GNAME46218(G46218,G46219,G43298);
  xor GNAME46219(G46219,G43388,G43478);
  and GNAME46220(G46220,G43388,G43298);
  and GNAME46221(G46221,G43478,G43298);
  and GNAME46222(G46222,G43388,G43478);
  or GNAME46223(G46223,G46222,G46221,G46220);
  xor GNAME46233(G46233,G46234,G43313);
  xor GNAME46234(G46234,G43403,G43493);
  and GNAME46235(G46235,G43403,G43313);
  and GNAME46236(G46236,G43493,G43313);
  and GNAME46237(G46237,G43403,G43493);
  or GNAME46238(G46238,G46237,G46236,G46235);
  xor GNAME46248(G46248,G46249,G43413);
  xor GNAME46249(G46249,G43323,G43233);
  and GNAME46250(G46250,G43323,G43413);
  and GNAME46251(G46251,G43233,G43413);
  and GNAME46252(G46252,G43323,G43233);
  or GNAME46253(G46253,G46252,G46251,G46250);
  xor GNAME46263(G46263,G46264,G43428);
  xor GNAME46264(G46264,G43338,G43248);
  and GNAME46265(G46265,G43338,G43428);
  and GNAME46266(G46266,G43248,G43428);
  and GNAME46267(G46267,G43338,G43248);
  or GNAME46268(G46268,G46267,G46266,G46265);
  xor GNAME46278(G46278,G46279,G43443);
  xor GNAME46279(G46279,G43353,G43263);
  and GNAME46280(G46280,G43353,G43443);
  and GNAME46281(G46281,G43263,G43443);
  and GNAME46282(G46282,G43353,G43263);
  or GNAME46283(G46283,G46282,G46281,G46280);
  xor GNAME46293(G46293,G46294,G43473);
  xor GNAME46294(G46294,G43383,G43293);
  and GNAME46295(G46295,G43383,G43473);
  and GNAME46296(G46296,G43293,G43473);
  and GNAME46297(G46297,G43383,G43293);
  or GNAME46298(G46298,G46297,G46296,G46295);
  xor GNAME46308(G46308,G46309,G43458);
  xor GNAME46309(G46309,G43368,G43278);
  and GNAME46310(G46310,G43368,G43458);
  and GNAME46311(G46311,G43278,G43458);
  and GNAME46312(G46312,G43368,G43278);
  or GNAME46313(G46313,G46312,G46311,G46310);
  xor GNAME46323(G46323,G46324,G43488);
  xor GNAME46324(G46324,G43398,G43308);
  and GNAME46325(G46325,G43398,G43488);
  and GNAME46326(G46326,G43308,G43488);
  and GNAME46327(G46327,G43398,G43308);
  or GNAME46328(G46328,G46327,G46326,G46325);
  xor GNAME46338(G46338,G46339,G46478);
  xor GNAME46339(G46339,G43508,G46428);
  and GNAME46340(G46340,G43508,G46478);
  and GNAME46341(G46341,G46428,G46478);
  and GNAME46342(G46342,G43508,G46428);
  or GNAME46343(G46343,G46342,G46341,G46340);
  xor GNAME46353(G46353,G46354,G43643);
  xor GNAME46354(G46354,G43868,G43503);
  and GNAME46355(G46355,G43868,G43643);
  and GNAME46356(G46356,G43503,G43643);
  and GNAME46357(G46357,G43868,G43503);
  or GNAME46358(G46358,G46357,G46356,G46355);
  xor GNAME46368(G46368,G46369,G46493);
  xor GNAME46369(G46369,G43523,G46443);
  and GNAME46370(G46370,G43523,G46493);
  and GNAME46371(G46371,G46443,G46493);
  and GNAME46372(G46372,G43523,G46443);
  or GNAME46373(G46373,G46372,G46371,G46370);
  xor GNAME46383(G46383,G46384,G43658);
  xor GNAME46384(G46384,G43883,G43518);
  and GNAME46385(G46385,G43883,G43658);
  and GNAME46386(G46386,G43518,G43658);
  and GNAME46387(G46387,G43883,G43518);
  or GNAME46388(G46388,G46387,G46386,G46385);
  xor GNAME46398(G46398,G46399,G46508);
  xor GNAME46399(G46399,G43538,G46458);
  and GNAME46400(G46400,G43538,G46508);
  and GNAME46401(G46401,G46458,G46508);
  and GNAME46402(G46402,G43538,G46458);
  or GNAME46403(G46403,G46402,G46401,G46400);
  xor GNAME46413(G46413,G46414,G43673);
  xor GNAME46414(G46414,G43898,G43533);
  and GNAME46415(G46415,G43898,G43673);
  and GNAME46416(G46416,G43533,G43673);
  and GNAME46417(G46417,G43898,G43533);
  or GNAME46418(G46418,G46417,G46416,G46415);
  xor GNAME46428(G46428,G46429,G43553);
  xor GNAME46429(G46429,G43688,G43733);
  and GNAME46430(G46430,G43688,G43553);
  and GNAME46431(G46431,G43733,G43553);
  and GNAME46432(G46432,G43688,G43733);
  or GNAME46433(G46433,G46432,G46431,G46430);
  xor GNAME46443(G46443,G46444,G43583);
  xor GNAME46444(G46444,G43703,G43763);
  and GNAME46445(G46445,G43703,G43583);
  and GNAME46446(G46446,G43763,G43583);
  and GNAME46447(G46447,G43703,G43763);
  or GNAME46448(G46448,G46447,G46446,G46445);
  xor GNAME46458(G46458,G46459,G43598);
  xor GNAME46459(G46459,G43718,G43778);
  and GNAME46460(G46460,G43718,G43598);
  and GNAME46461(G46461,G43778,G43598);
  and GNAME46462(G46462,G43718,G43778);
  or GNAME46463(G46463,G46462,G46461,G46460);
  xor GNAME46473(G46473,G46474,G43728);
  xor GNAME46474(G46474,G43683,G43548);
  and GNAME46475(G46475,G43683,G43728);
  and GNAME46476(G46476,G43548,G43728);
  and GNAME46477(G46477,G43683,G43548);
  or GNAME46478(G46478,G46477,G46476,G46475);
  xor GNAME46488(G46488,G46489,G43758);
  xor GNAME46489(G46489,G43698,G43578);
  and GNAME46490(G46490,G43698,G43758);
  and GNAME46491(G46491,G43578,G43758);
  and GNAME46492(G46492,G43698,G43578);
  or GNAME46493(G46493,G46492,G46491,G46490);
  xor GNAME46503(G46503,G46504,G43773);
  xor GNAME46504(G46504,G43713,G43593);
  and GNAME46505(G46505,G43713,G43773);
  and GNAME46506(G46506,G43593,G43773);
  and GNAME46507(G46507,G43713,G43593);
  or GNAME46508(G46508,G46507,G46506,G46505);
  xor GNAME46518(G46518,G46519,G43863);
  xor GNAME46519(G46519,G43958,G46658);
  and GNAME46520(G46520,G43958,G43863);
  and GNAME46521(G46521,G46658,G43863);
  and GNAME46522(G46522,G43958,G46658);
  or GNAME46523(G46523,G46522,G46521,G46520);
  xor GNAME46533(G46533,G46534,G44003);
  xor GNAME46534(G46534,G44043,G43953);
  and GNAME46535(G46535,G44043,G44003);
  and GNAME46536(G46536,G43953,G44003);
  and GNAME46537(G46537,G44043,G43953);
  or GNAME46538(G46538,G46537,G46536,G46535);
  xor GNAME46548(G46548,G46549,G43878);
  xor GNAME46549(G46549,G43973,G46673);
  and GNAME46550(G46550,G43973,G43878);
  and GNAME46551(G46551,G46673,G43878);
  and GNAME46552(G46552,G43973,G46673);
  or GNAME46553(G46553,G46552,G46551,G46550);
  xor GNAME46563(G46563,G46564,G44018);
  xor GNAME46564(G46564,G44073,G43968);
  and GNAME46565(G46565,G44073,G44018);
  and GNAME46566(G46566,G43968,G44018);
  and GNAME46567(G46567,G44073,G43968);
  or GNAME46568(G46568,G46567,G46566,G46565);
  xor GNAME46578(G46578,G46579,G43893);
  xor GNAME46579(G46579,G43988,G46688);
  and GNAME46580(G46580,G43988,G43893);
  and GNAME46581(G46581,G46688,G43893);
  and GNAME46582(G46582,G43988,G46688);
  or GNAME46583(G46583,G46582,G46581,G46580);
  xor GNAME46593(G46593,G46594,G44033);
  xor GNAME46594(G46594,G44088,G43983);
  and GNAME46595(G46595,G44088,G44033);
  and GNAME46596(G46596,G43983,G44033);
  and GNAME46597(G46597,G44088,G43983);
  or GNAME46598(G46598,G46597,G46596,G46595);
  xor GNAME46608(G46608,G46609,G46518);
  xor GNAME46609(G46609,G43638,G46538);
  and GNAME46610(G46610,G43638,G46518);
  and GNAME46611(G46611,G46538,G46518);
  and GNAME46612(G46612,G43638,G46538);
  or GNAME46613(G46613,G46612,G46611,G46610);
  xor GNAME46623(G46623,G46624,G46548);
  xor GNAME46624(G46624,G43653,G46568);
  and GNAME46625(G46625,G43653,G46548);
  and GNAME46626(G46626,G46568,G46548);
  and GNAME46627(G46627,G43653,G46568);
  or GNAME46628(G46628,G46627,G46626,G46625);
  xor GNAME46638(G46638,G46639,G46578);
  xor GNAME46639(G46639,G43668,G46598);
  and GNAME46640(G46640,G43668,G46578);
  and GNAME46641(G46641,G46598,G46578);
  and GNAME46642(G46642,G43668,G46598);
  or GNAME46643(G46643,G46642,G46641,G46640);
  xor GNAME46653(G46653,G46654,G43818);
  xor GNAME46654(G46654,G44063,G43913);
  and GNAME46655(G46655,G44063,G43818);
  and GNAME46656(G46656,G43913,G43818);
  and GNAME46657(G46657,G44063,G43913);
  or GNAME46658(G46658,G46657,G46656,G46655);
  xor GNAME46668(G46668,G46669,G43833);
  xor GNAME46669(G46669,G44108,G43928);
  and GNAME46670(G46670,G44108,G43833);
  and GNAME46671(G46671,G43928,G43833);
  and GNAME46672(G46672,G44108,G43928);
  or GNAME46673(G46673,G46672,G46671,G46670);
  xor GNAME46683(G46683,G46684,G43848);
  xor GNAME46684(G46684,G44123,G43943);
  and GNAME46685(G46685,G44123,G43848);
  and GNAME46686(G46686,G43943,G43848);
  and GNAME46687(G46687,G44123,G43943);
  or GNAME46688(G46688,G46687,G46686,G46685);
  xor GNAME46698(G46698,G46699,G44273);
  xor GNAME46699(G46699,G44058,G43908);
  and GNAME46700(G46700,G44058,G44273);
  and GNAME46701(G46701,G43908,G44273);
  and GNAME46702(G46702,G44058,G43908);
  or GNAME46703(G46703,G46702,G46701,G46700);
  xor GNAME46713(G46713,G46714,G44318);
  xor GNAME46714(G46714,G44403,G44178);
  and GNAME46715(G46715,G44403,G44318);
  and GNAME46716(G46716,G44178,G44318);
  and GNAME46717(G46717,G44403,G44178);
  or GNAME46718(G46718,G46717,G46716,G46715);
  xor GNAME46728(G46728,G46729,G44288);
  xor GNAME46729(G46729,G44103,G43923);
  and GNAME46730(G46730,G44103,G44288);
  and GNAME46731(G46731,G43923,G44288);
  and GNAME46732(G46732,G44103,G43923);
  or GNAME46733(G46733,G46732,G46731,G46730);
  xor GNAME46743(G46743,G46744,G44348);
  xor GNAME46744(G46744,G44418,G44208);
  and GNAME46745(G46745,G44418,G44348);
  and GNAME46746(G46746,G44208,G44348);
  and GNAME46747(G46747,G44418,G44208);
  or GNAME46748(G46748,G46747,G46746,G46745);
  xor GNAME46758(G46758,G46759,G44303);
  xor GNAME46759(G46759,G44118,G43938);
  and GNAME46760(G46760,G44118,G44303);
  and GNAME46761(G46761,G43938,G44303);
  and GNAME46762(G46762,G44118,G43938);
  or GNAME46763(G46763,G46762,G46761,G46760);
  xor GNAME46773(G46773,G46774,G44363);
  xor GNAME46774(G46774,G44433,G44223);
  and GNAME46775(G46775,G44433,G44363);
  and GNAME46776(G46776,G44223,G44363);
  and GNAME46777(G46777,G44433,G44223);
  or GNAME46778(G46778,G46777,G46776,G46775);
  xor GNAME46788(G46788,G46789,G46698);
  xor GNAME46789(G46789,G43998,G46718);
  and GNAME46790(G46790,G43998,G46698);
  and GNAME46791(G46791,G46718,G46698);
  and GNAME46792(G46792,G43998,G46718);
  or GNAME46793(G46793,G46792,G46791,G46790);
  xor GNAME46803(G46803,G46804,G46713);
  xor GNAME46804(G46804,G44268,G44138);
  and GNAME46805(G46805,G44268,G46713);
  and GNAME46806(G46806,G44138,G46713);
  and GNAME46807(G46807,G44268,G44138);
  or GNAME46808(G46808,G46807,G46806,G46805);
  xor GNAME46818(G46818,G46819,G44133);
  xor GNAME46819(G46819,G44313,G44498);
  and GNAME46820(G46820,G44313,G44133);
  and GNAME46821(G46821,G44498,G44133);
  and GNAME46822(G46822,G44313,G44498);
  or GNAME46823(G46823,G46822,G46821,G46820);
  xor GNAME46833(G46833,G46834,G46728);
  xor GNAME46834(G46834,G44013,G46748);
  and GNAME46835(G46835,G44013,G46728);
  and GNAME46836(G46836,G46748,G46728);
  and GNAME46837(G46837,G44013,G46748);
  or GNAME46838(G46838,G46837,G46836,G46835);
  xor GNAME46848(G46848,G46849,G46758);
  xor GNAME46849(G46849,G44028,G46778);
  and GNAME46850(G46850,G44028,G46758);
  and GNAME46851(G46851,G46778,G46758);
  and GNAME46852(G46852,G44028,G46778);
  or GNAME46853(G46853,G46852,G46851,G46850);
  xor GNAME46863(G46863,G46864,G46743);
  xor GNAME46864(G46864,G44283,G44153);
  and GNAME46865(G46865,G44283,G46743);
  and GNAME46866(G46866,G44153,G46743);
  and GNAME46867(G46867,G44283,G44153);
  or GNAME46868(G46868,G46867,G46866,G46865);
  xor GNAME46878(G46878,G46879,G44148);
  xor GNAME46879(G46879,G44343,G44528);
  and GNAME46880(G46880,G44343,G44148);
  and GNAME46881(G46881,G44528,G44148);
  and GNAME46882(G46882,G44343,G44528);
  or GNAME46883(G46883,G46882,G46881,G46880);
  xor GNAME46893(G46893,G46894,G46773);
  xor GNAME46894(G46894,G44298,G44168);
  and GNAME46895(G46895,G44298,G46773);
  and GNAME46896(G46896,G44168,G46773);
  and GNAME46897(G46897,G44298,G44168);
  or GNAME46898(G46898,G46897,G46896,G46895);
  xor GNAME46908(G46908,G46909,G44163);
  xor GNAME46909(G46909,G44358,G44543);
  and GNAME46910(G46910,G44358,G44163);
  and GNAME46911(G46911,G44543,G44163);
  and GNAME46912(G46912,G44358,G44543);
  or GNAME46913(G46913,G46912,G46911,G46910);
  xor GNAME46923(G46923,G46924,G44493);
  xor GNAME46924(G46924,G44328,G44513);
  and GNAME46925(G46925,G44328,G44493);
  and GNAME46926(G46926,G44513,G44493);
  and GNAME46927(G46927,G44328,G44513);
  or GNAME46928(G46928,G46927,G46926,G46925);
  xor GNAME46938(G46938,G46939,G44508);
  xor GNAME46939(G46939,G44628,G44768);
  and GNAME46940(G46940,G44628,G44508);
  and GNAME46941(G46941,G44768,G44508);
  and GNAME46942(G46942,G44628,G44768);
  or GNAME46943(G46943,G46942,G46941,G46940);
  xor GNAME46953(G46953,G46954,G44523);
  xor GNAME46954(G46954,G44373,G44558);
  and GNAME46955(G46955,G44373,G44523);
  and GNAME46956(G46956,G44558,G44523);
  and GNAME46957(G46957,G44373,G44558);
  or GNAME46958(G46958,G46957,G46956,G46955);
  xor GNAME46968(G46968,G46969,G44553);
  xor GNAME46969(G46969,G44643,G44783);
  and GNAME46970(G46970,G44643,G44553);
  and GNAME46971(G46971,G44783,G44553);
  and GNAME46972(G46972,G44643,G44783);
  or GNAME46973(G46973,G46972,G46971,G46970);
  xor GNAME46983(G46983,G46984,G44538);
  xor GNAME46984(G46984,G44388,G44573);
  and GNAME46985(G46985,G44388,G44538);
  and GNAME46986(G46986,G44573,G44538);
  and GNAME46987(G46987,G44388,G44573);
  or GNAME46988(G46988,G46987,G46986,G46985);
  xor GNAME46998(G46998,G46999,G44568);
  xor GNAME46999(G46999,G44658,G44798);
  and GNAME47000(G47000,G44658,G44568);
  and GNAME47001(G47001,G44798,G44568);
  and GNAME47002(G47002,G44658,G44798);
  or GNAME47003(G47003,G47002,G47001,G47000);
  xor GNAME47013(G47013,G47014,G44763);
  xor GNAME47014(G47014,G44723,G44583);
  and GNAME47015(G47015,G44723,G44763);
  and GNAME47016(G47016,G44583,G44763);
  and GNAME47017(G47017,G44723,G44583);
  or GNAME47018(G47018,G47017,G47016,G47015);
  xor GNAME47028(G47028,G47029,G44778);
  xor GNAME47029(G47029,G44738,G44598);
  and GNAME47030(G47030,G44738,G44778);
  and GNAME47031(G47031,G44598,G44778);
  and GNAME47032(G47032,G44738,G44598);
  or GNAME47033(G47033,G47032,G47031,G47030);
  xor GNAME47043(G47043,G47044,G44793);
  xor GNAME47044(G47044,G44753,G44613);
  and GNAME47045(G47045,G44753,G44793);
  and GNAME47046(G47046,G44613,G44793);
  and GNAME47047(G47047,G44753,G44613);
  or GNAME47048(G47048,G47047,G47046,G47045);
  xor GNAME47058(G47058,G47059,G47078);
  xor GNAME47059(G47059,G41073,G41123);
  and GNAME47060(G47060,G41073,G47078);
  and GNAME47061(G47061,G41123,G47078);
  and GNAME47062(G47062,G41073,G41123);
  or GNAME47063(G47063,G47062,G47061,G47060);
  xor GNAME47073(G47073,G47074,G47093);
  xor GNAME47074(G47074,G41258,G41118);
  and GNAME47075(G47075,G41258,G47093);
  and GNAME47076(G47076,G41118,G47093);
  and GNAME47077(G47077,G41258,G41118);
  or GNAME47078(G47078,G47077,G47076,G47075);
  xor GNAME47088(G47088,G47089,G48188);
  xor GNAME47089(G47089,G44993,G41253);
  and GNAME47090(G47090,G44993,G48188);
  and GNAME47091(G47091,G41253,G48188);
  and GNAME47092(G47092,G44993,G41253);
  or GNAME47093(G47093,G47092,G47091,G47090);
  xor GNAME47103(G47103,G47104,G47138);
  xor GNAME47104(G47104,G41088,G41138);
  and GNAME47105(G47105,G41088,G47138);
  and GNAME47106(G47106,G41138,G47138);
  and GNAME47107(G47107,G41088,G41138);
  or GNAME47108(G47108,G47107,G47106,G47105);
  xor GNAME47118(G47118,G47119,G47168);
  xor GNAME47119(G47119,G41103,G41153);
  and GNAME47120(G47120,G41103,G47168);
  and GNAME47121(G47121,G41153,G47168);
  and GNAME47122(G47122,G41103,G41153);
  or GNAME47123(G47123,G47122,G47121,G47120);
  xor GNAME47133(G47133,G47134,G47153);
  xor GNAME47134(G47134,G41273,G41133);
  and GNAME47135(G47135,G41273,G47153);
  and GNAME47136(G47136,G41133,G47153);
  and GNAME47137(G47137,G41273,G41133);
  or GNAME47138(G47138,G47137,G47136,G47135);
  xor GNAME47148(G47148,G47149,G48323);
  xor GNAME47149(G47149,G45008,G41268);
  and GNAME47150(G47150,G45008,G48323);
  and GNAME47151(G47151,G41268,G48323);
  and GNAME47152(G47152,G45008,G41268);
  or GNAME47153(G47153,G47152,G47151,G47150);
  xor GNAME47163(G47163,G47164,G47183);
  xor GNAME47164(G47164,G41288,G41148);
  and GNAME47165(G47165,G41288,G47183);
  and GNAME47166(G47166,G41148,G47183);
  and GNAME47167(G47167,G41288,G41148);
  or GNAME47168(G47168,G47167,G47166,G47165);
  xor GNAME47178(G47178,G47179,G48353);
  xor GNAME47179(G47179,G45023,G41283);
  and GNAME47180(G47180,G45023,G48353);
  and GNAME47181(G47181,G41283,G48353);
  and GNAME47182(G47182,G45023,G41283);
  or GNAME47183(G47183,G47182,G47181,G47180);
  xor GNAME47193(G47193,G47194,G47213);
  xor GNAME47194(G47194,G44828,G47013);
  and GNAME47195(G47195,G44828,G47213);
  and GNAME47196(G47196,G47013,G47213);
  and GNAME47197(G47197,G44828,G47013);
  or GNAME47198(G47198,G47197,G47196,G47195);
  xor GNAME47208(G47208,G47209,G44918);
  xor GNAME47209(G47209,G44813,G44823);
  and GNAME47210(G47210,G44813,G44918);
  and GNAME47211(G47211,G44823,G44918);
  and GNAME47212(G47212,G44813,G44823);
  or GNAME47213(G47213,G47212,G47211,G47210);
  xor GNAME47223(G47223,G47224,G47258);
  xor GNAME47224(G47224,G44843,G47028);
  and GNAME47225(G47225,G44843,G47258);
  and GNAME47226(G47226,G47028,G47258);
  and GNAME47227(G47227,G44843,G47028);
  or GNAME47228(G47228,G47227,G47226,G47225);
  xor GNAME47238(G47238,G47239,G47273);
  xor GNAME47239(G47239,G44858,G47043);
  and GNAME47240(G47240,G44858,G47273);
  and GNAME47241(G47241,G47043,G47273);
  and GNAME47242(G47242,G44858,G47043);
  or GNAME47243(G47243,G47242,G47241,G47240);
  xor GNAME47253(G47253,G47254,G44948);
  xor GNAME47254(G47254,G44873,G44838);
  and GNAME47255(G47255,G44873,G44948);
  and GNAME47256(G47256,G44838,G44948);
  and GNAME47257(G47257,G44873,G44838);
  or GNAME47258(G47258,G47257,G47256,G47255);
  xor GNAME47268(G47268,G47269,G44978);
  xor GNAME47269(G47269,G44888,G44853);
  and GNAME47270(G47270,G44888,G44978);
  and GNAME47271(G47271,G44853,G44978);
  and GNAME47272(G47272,G44888,G44853);
  or GNAME47273(G47273,G47272,G47271,G47270);
  xor GNAME47283(G47283,G47284,G47063);
  xor GNAME47284(G47284,G41078,G41028);
  and GNAME47285(G47285,G41078,G47063);
  and GNAME47286(G47286,G41028,G47063);
  and GNAME47287(G47287,G41078,G41028);
  or GNAME47288(G47288,G47287,G47286,G47285);
  xor GNAME47298(G47298,G47299,G47108);
  xor GNAME47299(G47299,G41093,G41043);
  and GNAME47300(G47300,G41093,G47108);
  and GNAME47301(G47301,G41043,G47108);
  and GNAME47302(G47302,G41093,G41043);
  or GNAME47303(G47303,G47302,G47301,G47300);
  xor GNAME47313(G47313,G47314,G47123);
  xor GNAME47314(G47314,G41108,G41058);
  and GNAME47315(G47315,G41108,G47123);
  and GNAME47316(G47316,G41058,G47123);
  and GNAME47317(G47317,G41108,G41058);
  or GNAME47318(G47318,G47317,G47316,G47315);
  xor GNAME47328(G47328,G47329,G45438);
  xor GNAME47329(G47329,G45393,G45458);
  and GNAME47330(G47330,G45393,G45438);
  and GNAME47331(G47331,G45458,G45438);
  and GNAME47332(G47332,G45393,G45458);
  or GNAME47333(G47333,G47332,G47331,G47330);
  xor GNAME47343(G47343,G47344,G45468);
  xor GNAME47344(G47344,G45408,G45488);
  and GNAME47345(G47345,G45408,G45468);
  and GNAME47346(G47346,G45488,G45468);
  and GNAME47347(G47347,G45408,G45488);
  or GNAME47348(G47348,G47347,G47346,G47345);
  xor GNAME47358(G47358,G47359,G45498);
  xor GNAME47359(G47359,G45423,G45518);
  and GNAME47360(G47360,G45423,G45498);
  and GNAME47361(G47361,G45518,G45498);
  and GNAME47362(G47362,G45423,G45518);
  or GNAME47363(G47363,G47362,G47361,G47360);
  xor GNAME47373(G47373,G47374,G45573);
  xor GNAME47374(G47374,G45668,G45713);
  and GNAME47375(G47375,G45668,G45573);
  and GNAME47376(G47376,G45713,G45573);
  and GNAME47377(G47377,G45668,G45713);
  or GNAME47378(G47378,G47377,G47376,G47375);
  xor GNAME47388(G47388,G47389,G45728);
  xor GNAME47389(G47389,G45803,G45663);
  and GNAME47390(G47390,G45803,G45728);
  and GNAME47391(G47391,G45663,G45728);
  and GNAME47392(G47392,G45803,G45663);
  or GNAME47393(G47393,G47392,G47391,G47390);
  xor GNAME47403(G47403,G47404,G45588);
  xor GNAME47404(G47404,G45683,G45743);
  and GNAME47405(G47405,G45683,G45588);
  and GNAME47406(G47406,G45743,G45588);
  and GNAME47407(G47407,G45683,G45743);
  or GNAME47408(G47408,G47407,G47406,G47405);
  xor GNAME47418(G47418,G47419,G45758);
  xor GNAME47419(G47419,G45833,G45678);
  and GNAME47420(G47420,G45833,G45758);
  and GNAME47421(G47421,G45678,G45758);
  and GNAME47422(G47422,G45833,G45678);
  or GNAME47423(G47423,G47422,G47421,G47420);
  xor GNAME47433(G47433,G47434,G45603);
  xor GNAME47434(G47434,G45698,G45773);
  and GNAME47435(G47435,G45698,G45603);
  and GNAME47436(G47436,G45773,G45603);
  and GNAME47437(G47437,G45698,G45773);
  or GNAME47438(G47438,G47437,G47436,G47435);
  xor GNAME47448(G47448,G47449,G45788);
  xor GNAME47449(G47449,G45848,G45693);
  and GNAME47450(G47450,G45848,G45788);
  and GNAME47451(G47451,G45693,G45788);
  and GNAME47452(G47452,G45848,G45693);
  or GNAME47453(G47453,G47452,G47451,G47450);
  xor GNAME47463(G47463,G47464,G47388);
  xor GNAME47464(G47464,G45708,G47513);
  and GNAME47465(G47465,G45708,G47388);
  and GNAME47466(G47466,G47513,G47388);
  and GNAME47467(G47467,G45708,G47513);
  or GNAME47468(G47468,G47467,G47466,G47465);
  xor GNAME47478(G47478,G47479,G47418);
  xor GNAME47479(G47479,G45738,G47543);
  and GNAME47480(G47480,G45738,G47418);
  and GNAME47481(G47481,G47543,G47418);
  and GNAME47482(G47482,G45738,G47543);
  or GNAME47483(G47483,G47482,G47481,G47480);
  xor GNAME47493(G47493,G47494,G47448);
  xor GNAME47494(G47494,G45768,G47573);
  and GNAME47495(G47495,G45768,G47448);
  and GNAME47496(G47496,G47573,G47448);
  and GNAME47497(G47497,G45768,G47573);
  or GNAME47498(G47498,G47497,G47496,G47495);
  xor GNAME47508(G47508,G47509,G45893);
  xor GNAME47509(G47509,G45818,G45798);
  and GNAME47510(G47510,G45818,G45893);
  and GNAME47511(G47511,G45798,G45893);
  and GNAME47512(G47512,G45818,G45798);
  or GNAME47513(G47513,G47512,G47511,G47510);
  xor GNAME47523(G47523,G47524,G45908);
  xor GNAME47524(G47524,G45983,G45813);
  and GNAME47525(G47525,G45983,G45908);
  and GNAME47526(G47526,G45813,G45908);
  and GNAME47527(G47527,G45983,G45813);
  or GNAME47528(G47528,G47527,G47526,G47525);
  xor GNAME47538(G47538,G47539,G45923);
  xor GNAME47539(G47539,G45863,G45828);
  and GNAME47540(G47540,G45863,G45923);
  and GNAME47541(G47541,G45828,G45923);
  and GNAME47542(G47542,G45863,G45828);
  or GNAME47543(G47543,G47542,G47541,G47540);
  xor GNAME47553(G47553,G47554,G45938);
  xor GNAME47554(G47554,G46013,G45858);
  and GNAME47555(G47555,G46013,G45938);
  and GNAME47556(G47556,G45858,G45938);
  and GNAME47557(G47557,G46013,G45858);
  or GNAME47558(G47558,G47557,G47556,G47555);
  xor GNAME47568(G47568,G47569,G45953);
  xor GNAME47569(G47569,G45878,G45843);
  and GNAME47570(G47570,G45878,G45953);
  and GNAME47571(G47571,G45843,G45953);
  and GNAME47572(G47572,G45878,G45843);
  or GNAME47573(G47573,G47572,G47571,G47570);
  xor GNAME47583(G47583,G47584,G45968);
  xor GNAME47584(G47584,G46028,G45873);
  and GNAME47585(G47585,G46028,G45968);
  and GNAME47586(G47586,G45873,G45968);
  and GNAME47587(G47587,G46028,G45873);
  or GNAME47588(G47588,G47587,G47586,G47585);
  xor GNAME47598(G47598,G47599,G47508);
  xor GNAME47599(G47599,G45723,G47528);
  and GNAME47600(G47600,G45723,G47508);
  and GNAME47601(G47601,G47528,G47508);
  and GNAME47602(G47602,G45723,G47528);
  or GNAME47603(G47603,G47602,G47601,G47600);
  xor GNAME47613(G47613,G47614,G47523);
  xor GNAME47614(G47614,G45888,G47693);
  and GNAME47615(G47615,G45888,G47523);
  and GNAME47616(G47616,G47693,G47523);
  and GNAME47617(G47617,G45888,G47693);
  or GNAME47618(G47618,G47617,G47616,G47615);
  xor GNAME47628(G47628,G47629,G47538);
  xor GNAME47629(G47629,G45753,G47558);
  and GNAME47630(G47630,G45753,G47538);
  and GNAME47631(G47631,G47558,G47538);
  and GNAME47632(G47632,G45753,G47558);
  or GNAME47633(G47633,G47632,G47631,G47630);
  xor GNAME47643(G47643,G47644,G47568);
  xor GNAME47644(G47644,G45783,G47588);
  and GNAME47645(G47645,G45783,G47568);
  and GNAME47646(G47646,G47588,G47568);
  and GNAME47647(G47647,G45783,G47588);
  or GNAME47648(G47648,G47647,G47646,G47645);
  xor GNAME47658(G47658,G47659,G47553);
  xor GNAME47659(G47659,G45918,G47723);
  and GNAME47660(G47660,G45918,G47553);
  and GNAME47661(G47661,G47723,G47553);
  and GNAME47662(G47662,G45918,G47723);
  or GNAME47663(G47663,G47662,G47661,G47660);
  xor GNAME47673(G47673,G47674,G47583);
  xor GNAME47674(G47674,G45948,G47753);
  and GNAME47675(G47675,G45948,G47583);
  and GNAME47676(G47676,G47753,G47583);
  and GNAME47677(G47677,G45948,G47753);
  or GNAME47678(G47678,G47677,G47676,G47675);
  xor GNAME47688(G47688,G47689,G46073);
  xor GNAME47689(G47689,G45998,G45978);
  and GNAME47690(G47690,G45998,G46073);
  and GNAME47691(G47691,G45978,G46073);
  and GNAME47692(G47692,G45998,G45978);
  or GNAME47693(G47693,G47692,G47691,G47690);
  xor GNAME47703(G47703,G47704,G46088);
  xor GNAME47704(G47704,G46163,G45993);
  and GNAME47705(G47705,G46163,G46088);
  and GNAME47706(G47706,G45993,G46088);
  and GNAME47707(G47707,G46163,G45993);
  or GNAME47708(G47708,G47707,G47706,G47705);
  xor GNAME47718(G47718,G47719,G46103);
  xor GNAME47719(G47719,G46043,G46008);
  and GNAME47720(G47720,G46043,G46103);
  and GNAME47721(G47721,G46008,G46103);
  and GNAME47722(G47722,G46043,G46008);
  or GNAME47723(G47723,G47722,G47721,G47720);
  xor GNAME47733(G47733,G47734,G46118);
  xor GNAME47734(G47734,G46193,G46038);
  and GNAME47735(G47735,G46193,G46118);
  and GNAME47736(G47736,G46038,G46118);
  and GNAME47737(G47737,G46193,G46038);
  or GNAME47738(G47738,G47737,G47736,G47735);
  xor GNAME47748(G47748,G47749,G46133);
  xor GNAME47749(G47749,G46058,G46023);
  and GNAME47750(G47750,G46058,G46133);
  and GNAME47751(G47751,G46023,G46133);
  and GNAME47752(G47752,G46058,G46023);
  or GNAME47753(G47753,G47752,G47751,G47750);
  xor GNAME47763(G47763,G47764,G46148);
  xor GNAME47764(G47764,G46208,G46053);
  and GNAME47765(G47765,G46208,G46148);
  and GNAME47766(G47766,G46053,G46148);
  and GNAME47767(G47767,G46208,G46053);
  or GNAME47768(G47768,G47767,G47766,G47765);
  xor GNAME47778(G47778,G47779,G47688);
  xor GNAME47779(G47779,G45903,G47708);
  and GNAME47780(G47780,G45903,G47688);
  and GNAME47781(G47781,G47708,G47688);
  and GNAME47782(G47782,G45903,G47708);
  or GNAME47783(G47783,G47782,G47781,G47780);
  xor GNAME47793(G47793,G47794,G47703);
  xor GNAME47794(G47794,G46068,G47873);
  and GNAME47795(G47795,G46068,G47703);
  and GNAME47796(G47796,G47873,G47703);
  and GNAME47797(G47797,G46068,G47873);
  or GNAME47798(G47798,G47797,G47796,G47795);
  xor GNAME47808(G47808,G47809,G47718);
  xor GNAME47809(G47809,G45933,G47738);
  and GNAME47810(G47810,G45933,G47718);
  and GNAME47811(G47811,G47738,G47718);
  and GNAME47812(G47812,G45933,G47738);
  or GNAME47813(G47813,G47812,G47811,G47810);
  xor GNAME47823(G47823,G47824,G47748);
  xor GNAME47824(G47824,G45963,G47768);
  and GNAME47825(G47825,G45963,G47748);
  and GNAME47826(G47826,G47768,G47748);
  and GNAME47827(G47827,G45963,G47768);
  or GNAME47828(G47828,G47827,G47826,G47825);
  xor GNAME47838(G47838,G47839,G47733);
  xor GNAME47839(G47839,G46098,G47903);
  and GNAME47840(G47840,G46098,G47733);
  and GNAME47841(G47841,G47903,G47733);
  and GNAME47842(G47842,G46098,G47903);
  or GNAME47843(G47843,G47842,G47841,G47840);
  xor GNAME47853(G47853,G47854,G47763);
  xor GNAME47854(G47854,G46128,G47933);
  and GNAME47855(G47855,G46128,G47763);
  and GNAME47856(G47856,G47933,G47763);
  and GNAME47857(G47857,G46128,G47933);
  or GNAME47858(G47858,G47857,G47856,G47855);
  xor GNAME47868(G47868,G47869,G46253);
  xor GNAME47869(G47869,G46178,G46158);
  and GNAME47870(G47870,G46178,G46253);
  and GNAME47871(G47871,G46158,G46253);
  and GNAME47872(G47872,G46178,G46158);
  or GNAME47873(G47873,G47872,G47871,G47870);
  xor GNAME47883(G47883,G47884,G46268);
  xor GNAME47884(G47884,G46433,G46173);
  and GNAME47885(G47885,G46433,G46268);
  and GNAME47886(G47886,G46173,G46268);
  and GNAME47887(G47887,G46433,G46173);
  or GNAME47888(G47888,G47887,G47886,G47885);
  xor GNAME47898(G47898,G47899,G46283);
  xor GNAME47899(G47899,G46223,G46188);
  and GNAME47900(G47900,G46223,G46283);
  and GNAME47901(G47901,G46188,G46283);
  and GNAME47902(G47902,G46223,G46188);
  or GNAME47903(G47903,G47902,G47901,G47900);
  xor GNAME47913(G47913,G47914,G46298);
  xor GNAME47914(G47914,G46448,G46218);
  and GNAME47915(G47915,G46448,G46298);
  and GNAME47916(G47916,G46218,G46298);
  and GNAME47917(G47917,G46448,G46218);
  or GNAME47918(G47918,G47917,G47916,G47915);
  xor GNAME47928(G47928,G47929,G46313);
  xor GNAME47929(G47929,G46238,G46203);
  and GNAME47930(G47930,G46238,G46313);
  and GNAME47931(G47931,G46203,G46313);
  and GNAME47932(G47932,G46238,G46203);
  or GNAME47933(G47933,G47932,G47931,G47930);
  xor GNAME47943(G47943,G47944,G46328);
  xor GNAME47944(G47944,G46463,G46233);
  and GNAME47945(G47945,G46463,G46328);
  and GNAME47946(G47946,G46233,G46328);
  and GNAME47947(G47947,G46463,G46233);
  or GNAME47948(G47948,G47947,G47946,G47945);
  xor GNAME47958(G47958,G47959,G47868);
  xor GNAME47959(G47959,G46083,G47888);
  and GNAME47960(G47960,G46083,G47868);
  and GNAME47961(G47961,G47888,G47868);
  and GNAME47962(G47962,G46083,G47888);
  or GNAME47963(G47963,G47962,G47961,G47960);
  xor GNAME47973(G47973,G47974,G47883);
  xor GNAME47974(G47974,G46248,G46343);
  and GNAME47975(G47975,G46248,G47883);
  and GNAME47976(G47976,G46343,G47883);
  and GNAME47977(G47977,G46248,G46343);
  or GNAME47978(G47978,G47977,G47976,G47975);
  xor GNAME47988(G47988,G47989,G47898);
  xor GNAME47989(G47989,G46113,G47918);
  and GNAME47990(G47990,G46113,G47898);
  and GNAME47991(G47991,G47918,G47898);
  and GNAME47992(G47992,G46113,G47918);
  or GNAME47993(G47993,G47992,G47991,G47990);
  xor GNAME48003(G48003,G48004,G47928);
  xor GNAME48004(G48004,G46143,G47948);
  and GNAME48005(G48005,G46143,G47928);
  and GNAME48006(G48006,G47948,G47928);
  and GNAME48007(G48007,G46143,G47948);
  or GNAME48008(G48008,G48007,G48006,G48005);
  xor GNAME48018(G48018,G48019,G47913);
  xor GNAME48019(G48019,G46278,G46373);
  and GNAME48020(G48020,G46278,G47913);
  and GNAME48021(G48021,G46373,G47913);
  and GNAME48022(G48022,G46278,G46373);
  or GNAME48023(G48023,G48022,G48021,G48020);
  xor GNAME48033(G48033,G48034,G47943);
  xor GNAME48034(G48034,G46308,G46403);
  and GNAME48035(G48035,G46308,G47943);
  and GNAME48036(G48036,G46403,G47943);
  and GNAME48037(G48037,G46308,G46403);
  or GNAME48038(G48038,G48037,G48036,G48035);
  xor GNAME48048(G48048,G48049,G46338);
  xor GNAME48049(G48049,G46263,G46358);
  and GNAME48050(G48050,G46263,G46338);
  and GNAME48051(G48051,G46358,G46338);
  and GNAME48052(G48052,G46263,G46358);
  or GNAME48053(G48053,G48052,G48051,G48050);
  xor GNAME48063(G48063,G48064,G46353);
  xor GNAME48064(G48064,G46473,G46523);
  and GNAME48065(G48065,G46473,G46353);
  and GNAME48066(G48066,G46523,G46353);
  and GNAME48067(G48067,G46473,G46523);
  or GNAME48068(G48068,G48067,G48066,G48065);
  xor GNAME48078(G48078,G48079,G46368);
  xor GNAME48079(G48079,G46293,G46388);
  and GNAME48080(G48080,G46293,G46368);
  and GNAME48081(G48081,G46388,G46368);
  and GNAME48082(G48082,G46293,G46388);
  or GNAME48083(G48083,G48082,G48081,G48080);
  xor GNAME48093(G48093,G48094,G46398);
  xor GNAME48094(G48094,G46323,G46418);
  and GNAME48095(G48095,G46323,G46398);
  and GNAME48096(G48096,G46418,G46398);
  and GNAME48097(G48097,G46323,G46418);
  or GNAME48098(G48098,G48097,G48096,G48095);
  xor GNAME48108(G48108,G48109,G46383);
  xor GNAME48109(G48109,G46488,G46553);
  and GNAME48110(G48110,G46488,G46383);
  and GNAME48111(G48111,G46553,G46383);
  and GNAME48112(G48112,G46488,G46553);
  or GNAME48113(G48113,G48112,G48111,G48110);
  xor GNAME48123(G48123,G48124,G46413);
  xor GNAME48124(G48124,G46503,G46583);
  and GNAME48125(G48125,G46503,G46413);
  and GNAME48126(G48126,G46583,G46413);
  and GNAME48127(G48127,G46503,G46583);
  or GNAME48128(G48128,G48127,G48126,G48125);
  xor GNAME48138(G48138,G48139,G46533);
  xor GNAME48139(G48139,G46653,G46703);
  and GNAME48140(G48140,G46653,G46533);
  and GNAME48141(G48141,G46703,G46533);
  and GNAME48142(G48142,G46653,G46703);
  or GNAME48143(G48143,G48142,G48141,G48140);
  xor GNAME48153(G48153,G48154,G46563);
  xor GNAME48154(G48154,G46668,G46733);
  and GNAME48155(G48155,G46668,G46563);
  and GNAME48156(G48156,G46733,G46563);
  and GNAME48157(G48157,G46668,G46733);
  or GNAME48158(G48158,G48157,G48156,G48155);
  xor GNAME48168(G48168,G48169,G46593);
  xor GNAME48169(G48169,G46683,G46763);
  and GNAME48170(G48170,G46683,G46593);
  and GNAME48171(G48171,G46763,G46593);
  and GNAME48172(G48172,G46683,G46763);
  or GNAME48173(G48173,G48172,G48171,G48170);
  xor GNAME48183(G48183,G48184,G48203);
  xor GNAME48184(G48184,G44988,G45038);
  and GNAME48185(G48185,G44988,G48203);
  and GNAME48186(G48186,G45038,G48203);
  and GNAME48187(G48187,G44988,G45038);
  or GNAME48188(G48188,G48187,G48186,G48185);
  xor GNAME48198(G48198,G48199,G48218);
  xor GNAME48199(G48199,G45033,G45128);
  and GNAME48200(G48200,G45033,G48218);
  and GNAME48201(G48201,G45128,G48218);
  and GNAME48202(G48202,G45033,G45128);
  or GNAME48203(G48203,G48202,G48201,G48200);
  xor GNAME48213(G48213,G48214,G48233);
  xor GNAME48214(G48214,G45143,G45123);
  and GNAME48215(G48215,G45143,G48233);
  and GNAME48216(G48216,G45123,G48233);
  and GNAME48217(G48217,G45143,G45123);
  or GNAME48218(G48218,G48217,G48216,G48215);
  xor GNAME48228(G48228,G48229,G48248);
  xor GNAME48229(G48229,G45308,G45138);
  and GNAME48230(G48230,G45308,G48248);
  and GNAME48231(G48231,G45138,G48248);
  and GNAME48232(G48232,G45308,G45138);
  or GNAME48233(G48233,G48232,G48231,G48230);
  xor GNAME48243(G48243,G48244,G48263);
  xor GNAME48244(G48244,G45323,G45303);
  and GNAME48245(G48245,G45323,G48263);
  and GNAME48246(G48246,G45303,G48263);
  and GNAME48247(G48247,G45323,G45303);
  or GNAME48248(G48248,G48247,G48246,G48245);
  xor GNAME48258(G48258,G48259,G48278);
  xor GNAME48259(G48259,G47333,G45318);
  and GNAME48260(G48260,G47333,G48278);
  and GNAME48261(G48261,G45318,G48278);
  and GNAME48262(G48262,G47333,G45318);
  or GNAME48263(G48263,G48262,G48261,G48260);
  xor GNAME48273(G48273,G48274,G48293);
  xor GNAME48274(G48274,G45533,G47328);
  and GNAME48275(G48275,G45533,G48293);
  and GNAME48276(G48276,G47328,G48293);
  and GNAME48277(G48277,G45533,G47328);
  or GNAME48278(G48278,G48277,G48276,G48275);
  xor GNAME48288(G48288,G48289,G48308);
  xor GNAME48289(G48289,G45623,G45528);
  and GNAME48290(G48290,G45623,G48308);
  and GNAME48291(G48291,G45528,G48308);
  and GNAME48292(G48292,G45623,G45528);
  or GNAME48293(G48293,G48292,G48291,G48290);
  xor GNAME48303(G48303,G48304,G48953);
  xor GNAME48304(G48304,G47468,G45618);
  and GNAME48305(G48305,G47468,G48953);
  and GNAME48306(G48306,G45618,G48953);
  and GNAME48307(G48307,G47468,G45618);
  or GNAME48308(G48308,G48307,G48306,G48305);
  xor GNAME48318(G48318,G48319,G48338);
  xor GNAME48319(G48319,G45003,G45053);
  and GNAME48320(G48320,G45003,G48338);
  and GNAME48321(G48321,G45053,G48338);
  and GNAME48322(G48322,G45003,G45053);
  or GNAME48323(G48323,G48322,G48321,G48320);
  xor GNAME48333(G48333,G48334,G48383);
  xor GNAME48334(G48334,G45048,G45158);
  and GNAME48335(G48335,G45048,G48383);
  and GNAME48336(G48336,G45158,G48383);
  and GNAME48337(G48337,G45048,G45158);
  or GNAME48338(G48338,G48337,G48336,G48335);
  xor GNAME48348(G48348,G48349,G48368);
  xor GNAME48349(G48349,G45018,G45068);
  and GNAME48350(G48350,G45018,G48368);
  and GNAME48351(G48351,G45068,G48368);
  and GNAME48352(G48352,G45018,G45068);
  or GNAME48353(G48353,G48352,G48351,G48350);
  xor GNAME48363(G48363,G48364,G48428);
  xor GNAME48364(G48364,G45063,G45173);
  and GNAME48365(G48365,G45063,G48428);
  and GNAME48366(G48366,G45173,G48428);
  and GNAME48367(G48367,G45063,G45173);
  or GNAME48368(G48368,G48367,G48366,G48365);
  xor GNAME48378(G48378,G48379,G48398);
  xor GNAME48379(G48379,G45188,G45153);
  and GNAME48380(G48380,G45188,G48398);
  and GNAME48381(G48381,G45153,G48398);
  and GNAME48382(G48382,G45188,G45153);
  or GNAME48383(G48383,G48382,G48381,G48380);
  xor GNAME48393(G48393,G48394,G48458);
  xor GNAME48394(G48394,G45338,G45183);
  and GNAME48395(G48395,G45338,G48458);
  and GNAME48396(G48396,G45183,G48458);
  and GNAME48397(G48397,G45338,G45183);
  or GNAME48398(G48398,G48397,G48396,G48395);
  xor GNAME48408(G48408,G48409,G48488);
  xor GNAME48409(G48409,G46613,G48063);
  and GNAME48410(G48410,G46613,G48488);
  and GNAME48411(G48411,G48063,G48488);
  and GNAME48412(G48412,G46613,G48063);
  or GNAME48413(G48413,G48412,G48411,G48410);
  xor GNAME48423(G48423,G48424,G48443);
  xor GNAME48424(G48424,G45203,G45168);
  and GNAME48425(G48425,G45203,G48443);
  and GNAME48426(G48426,G45168,G48443);
  and GNAME48427(G48427,G45203,G45168);
  or GNAME48428(G48428,G48427,G48426,G48425);
  xor GNAME48438(G48438,G48439,G48548);
  xor GNAME48439(G48439,G45353,G45198);
  and GNAME48440(G48440,G45353,G48548);
  and GNAME48441(G48441,G45198,G48548);
  and GNAME48442(G48442,G45353,G45198);
  or GNAME48443(G48443,G48442,G48441,G48440);
  xor GNAME48453(G48453,G48454,G48473);
  xor GNAME48454(G48454,G45368,G45333);
  and GNAME48455(G48455,G45368,G48473);
  and GNAME48456(G48456,G45333,G48473);
  and GNAME48457(G48457,G45368,G45333);
  or GNAME48458(G48458,G48457,G48456,G48455);
  xor GNAME48468(G48468,G48469,G48578);
  xor GNAME48469(G48469,G47348,G45363);
  and GNAME48470(G48470,G47348,G48578);
  and GNAME48471(G48471,G45363,G48578);
  and GNAME48472(G48472,G47348,G45363);
  or GNAME48473(G48473,G48472,G48471,G48470);
  xor GNAME48483(G48483,G48484,G48503);
  xor GNAME48484(G48484,G48143,G46608);
  and GNAME48485(G48485,G48143,G48503);
  and GNAME48486(G48486,G46608,G48503);
  and GNAME48487(G48487,G48143,G46608);
  or GNAME48488(G48488,G48487,G48486,G48485);
  xor GNAME48498(G48498,G48499,G48518);
  xor GNAME48499(G48499,G46793,G48138);
  and GNAME48500(G48500,G46793,G48518);
  and GNAME48501(G48501,G48138,G48518);
  and GNAME48502(G48502,G46793,G48138);
  or GNAME48503(G48503,G48502,G48501,G48500);
  xor GNAME48513(G48513,G48514,G48533);
  xor GNAME48514(G48514,G46808,G46788);
  and GNAME48515(G48515,G46808,G48533);
  and GNAME48516(G48516,G46788,G48533);
  and GNAME48517(G48517,G46808,G46788);
  or GNAME48518(G48518,G48517,G48516,G48515);
  xor GNAME48528(G48528,G48529,G48608);
  xor GNAME48529(G48529,G46823,G46803);
  and GNAME48530(G48530,G46823,G48608);
  and GNAME48531(G48531,G46803,G48608);
  and GNAME48532(G48532,G46823,G46803);
  or GNAME48533(G48533,G48532,G48531,G48530);
  xor GNAME48543(G48543,G48544,G48563);
  xor GNAME48544(G48544,G45383,G45348);
  and GNAME48545(G48545,G45383,G48563);
  and GNAME48546(G48546,G45348,G48563);
  and GNAME48547(G48547,G45383,G45348);
  or GNAME48548(G48548,G48547,G48546,G48545);
  xor GNAME48558(G48558,G48559,G48653);
  xor GNAME48559(G48559,G47363,G45378);
  and GNAME48560(G48560,G47363,G48653);
  and GNAME48561(G48561,G45378,G48653);
  and GNAME48562(G48562,G47363,G45378);
  or GNAME48563(G48563,G48562,G48561,G48560);
  xor GNAME48573(G48573,G48574,G48593);
  xor GNAME48574(G48574,G45548,G47343);
  and GNAME48575(G48575,G45548,G48593);
  and GNAME48576(G48576,G47343,G48593);
  and GNAME48577(G48577,G45548,G47343);
  or GNAME48578(G48578,G48577,G48576,G48575);
  xor GNAME48588(G48588,G48589,G48683);
  xor GNAME48589(G48589,G45638,G45543);
  and GNAME48590(G48590,G45638,G48683);
  and GNAME48591(G48591,G45543,G48683);
  and GNAME48592(G48592,G45638,G45543);
  or GNAME48593(G48593,G48592,G48591,G48590);
  xor GNAME48603(G48603,G48604,G48623);
  xor GNAME48604(G48604,G46928,G46818);
  and GNAME48605(G48605,G46928,G48623);
  and GNAME48606(G48606,G46818,G48623);
  and GNAME48607(G48607,G46928,G46818);
  or GNAME48608(G48608,G48607,G48606,G48605);
  xor GNAME48618(G48618,G48619,G48638);
  xor GNAME48619(G48619,G46943,G46923);
  and GNAME48620(G48620,G46943,G48638);
  and GNAME48621(G48621,G46923,G48638);
  and GNAME48622(G48622,G46943,G46923);
  or GNAME48623(G48623,G48622,G48621,G48620);
  xor GNAME48633(G48633,G48634,G47198);
  xor GNAME48634(G48634,G47018,G46938);
  and GNAME48635(G48635,G47018,G47198);
  and GNAME48636(G48636,G46938,G47198);
  and GNAME48637(G48637,G47018,G46938);
  or GNAME48638(G48638,G48637,G48636,G48635);
  xor GNAME48648(G48648,G48649,G48668);
  xor GNAME48649(G48649,G45563,G47358);
  and GNAME48650(G48650,G45563,G48668);
  and GNAME48651(G48651,G47358,G48668);
  and GNAME48652(G48652,G45563,G47358);
  or GNAME48653(G48653,G48652,G48651,G48650);
  xor GNAME48663(G48663,G48664,G48698);
  xor GNAME48664(G48664,G45653,G45558);
  and GNAME48665(G48665,G45653,G48698);
  and GNAME48666(G48666,G45558,G48698);
  and GNAME48667(G48667,G45653,G45558);
  or GNAME48668(G48668,G48667,G48666,G48665);
  xor GNAME48678(G48678,G48679,G49073);
  xor GNAME48679(G48679,G47483,G45633);
  and GNAME48680(G48680,G47483,G49073);
  and GNAME48681(G48681,G45633,G49073);
  and GNAME48682(G48682,G47483,G45633);
  or GNAME48683(G48683,G48682,G48681,G48680);
  xor GNAME48693(G48693,G48694,G49088);
  xor GNAME48694(G48694,G47498,G45648);
  and GNAME48695(G48695,G47498,G49088);
  and GNAME48696(G48696,G45648,G49088);
  and GNAME48697(G48697,G47498,G45648);
  or GNAME48698(G48698,G48697,G48696,G48695);
  xor GNAME48708(G48708,G48709,G48743);
  xor GNAME48709(G48709,G46628,G48108);
  and GNAME48710(G48710,G46628,G48743);
  and GNAME48711(G48711,G48108,G48743);
  and GNAME48712(G48712,G46628,G48108);
  or GNAME48713(G48713,G48712,G48711,G48710);
  xor GNAME48723(G48723,G48724,G48773);
  xor GNAME48724(G48724,G46643,G48123);
  and GNAME48725(G48725,G46643,G48773);
  and GNAME48726(G48726,G48123,G48773);
  and GNAME48727(G48727,G46643,G48123);
  or GNAME48728(G48728,G48727,G48726,G48725);
  xor GNAME48738(G48738,G48739,G48758);
  xor GNAME48739(G48739,G48158,G46623);
  and GNAME48740(G48740,G48158,G48758);
  and GNAME48741(G48741,G46623,G48758);
  and GNAME48742(G48742,G48158,G46623);
  or GNAME48743(G48743,G48742,G48741,G48740);
  xor GNAME48753(G48753,G48754,G48803);
  xor GNAME48754(G48754,G46838,G48153);
  and GNAME48755(G48755,G46838,G48803);
  and GNAME48756(G48756,G48153,G48803);
  and GNAME48757(G48757,G46838,G48153);
  or GNAME48758(G48758,G48757,G48756,G48755);
  xor GNAME48768(G48768,G48769,G48788);
  xor GNAME48769(G48769,G48173,G46638);
  and GNAME48770(G48770,G48173,G48788);
  and GNAME48771(G48771,G46638,G48788);
  and GNAME48772(G48772,G48173,G46638);
  or GNAME48773(G48773,G48772,G48771,G48770);
  xor GNAME48783(G48783,G48784,G48833);
  xor GNAME48784(G48784,G46853,G48168);
  and GNAME48785(G48785,G46853,G48833);
  and GNAME48786(G48786,G48168,G48833);
  and GNAME48787(G48787,G46853,G48168);
  or GNAME48788(G48788,G48787,G48786,G48785);
  xor GNAME48798(G48798,G48799,G48818);
  xor GNAME48799(G48799,G46868,G46833);
  and GNAME48800(G48800,G46868,G48818);
  and GNAME48801(G48801,G46833,G48818);
  and GNAME48802(G48802,G46868,G46833);
  or GNAME48803(G48803,G48802,G48801,G48800);
  xor GNAME48813(G48813,G48814,G48863);
  xor GNAME48814(G48814,G46883,G46863);
  and GNAME48815(G48815,G46883,G48863);
  and GNAME48816(G48816,G46863,G48863);
  and GNAME48817(G48817,G46883,G46863);
  or GNAME48818(G48818,G48817,G48816,G48815);
  xor GNAME48828(G48828,G48829,G48848);
  xor GNAME48829(G48829,G46898,G46848);
  and GNAME48830(G48830,G46898,G48848);
  and GNAME48831(G48831,G46848,G48848);
  and GNAME48832(G48832,G46898,G46848);
  or GNAME48833(G48833,G48832,G48831,G48830);
  xor GNAME48843(G48843,G48844,G48893);
  xor GNAME48844(G48844,G46913,G46893);
  and GNAME48845(G48845,G46913,G48893);
  and GNAME48846(G48846,G46893,G48893);
  and GNAME48847(G48847,G46913,G46893);
  or GNAME48848(G48848,G48847,G48846,G48845);
  xor GNAME48858(G48858,G48859,G48878);
  xor GNAME48859(G48859,G46958,G46878);
  and GNAME48860(G48860,G46958,G48878);
  and GNAME48861(G48861,G46878,G48878);
  and GNAME48862(G48862,G46958,G46878);
  or GNAME48863(G48863,G48862,G48861,G48860);
  xor GNAME48873(G48873,G48874,G48923);
  xor GNAME48874(G48874,G46973,G46953);
  and GNAME48875(G48875,G46973,G48923);
  and GNAME48876(G48876,G46953,G48923);
  and GNAME48877(G48877,G46973,G46953);
  or GNAME48878(G48878,G48877,G48876,G48875);
  xor GNAME48888(G48888,G48889,G48908);
  xor GNAME48889(G48889,G46988,G46908);
  and GNAME48890(G48890,G46988,G48908);
  and GNAME48891(G48891,G46908,G48908);
  and GNAME48892(G48892,G46988,G46908);
  or GNAME48893(G48893,G48892,G48891,G48890);
  xor GNAME48903(G48903,G48904,G48938);
  xor GNAME48904(G48904,G47003,G46983);
  and GNAME48905(G48905,G47003,G48938);
  and GNAME48906(G48906,G46983,G48938);
  and GNAME48907(G48907,G47003,G46983);
  or GNAME48908(G48908,G48907,G48906,G48905);
  xor GNAME48918(G48918,G48919,G47228);
  xor GNAME48919(G48919,G47033,G46968);
  and GNAME48920(G48920,G47033,G47228);
  and GNAME48921(G48921,G46968,G47228);
  and GNAME48922(G48922,G47033,G46968);
  or GNAME48923(G48923,G48922,G48921,G48920);
  xor GNAME48933(G48933,G48934,G47243);
  xor GNAME48934(G48934,G47048,G46998);
  and GNAME48935(G48935,G47048,G47243);
  and GNAME48936(G48936,G46998,G47243);
  and GNAME48937(G48937,G47048,G46998);
  or GNAME48938(G48938,G48937,G48936,G48935);
  xor GNAME48948(G48948,G48949,G48968);
  xor GNAME48949(G48949,G47603,G47463);
  and GNAME48950(G48950,G47603,G48968);
  and GNAME48951(G48951,G47463,G48968);
  and GNAME48952(G48952,G47603,G47463);
  or GNAME48953(G48953,G48952,G48951,G48950);
  xor GNAME48963(G48963,G48964,G48983);
  xor GNAME48964(G48964,G47618,G47598);
  and GNAME48965(G48965,G47618,G48983);
  and GNAME48966(G48966,G47598,G48983);
  and GNAME48967(G48967,G47618,G47598);
  or GNAME48968(G48968,G48967,G48966,G48965);
  xor GNAME48978(G48978,G48979,G48998);
  xor GNAME48979(G48979,G47783,G47613);
  and GNAME48980(G48980,G47783,G48998);
  and GNAME48981(G48981,G47613,G48998);
  and GNAME48982(G48982,G47783,G47613);
  or GNAME48983(G48983,G48982,G48981,G48980);
  xor GNAME48993(G48993,G48994,G49013);
  xor GNAME48994(G48994,G47798,G47778);
  and GNAME48995(G48995,G47798,G49013);
  and GNAME48996(G48996,G47778,G49013);
  and GNAME48997(G48997,G47798,G47778);
  or GNAME48998(G48998,G48997,G48996,G48995);
  xor GNAME49008(G49008,G49009,G49028);
  xor GNAME49009(G49009,G47963,G47793);
  and GNAME49010(G49010,G47963,G49028);
  and GNAME49011(G49011,G47793,G49028);
  and GNAME49012(G49012,G47963,G47793);
  or GNAME49013(G49013,G49012,G49011,G49010);
  xor GNAME49023(G49023,G49024,G49043);
  xor GNAME49024(G49024,G47978,G47958);
  and GNAME49025(G49025,G47978,G49043);
  and GNAME49026(G49026,G47958,G49043);
  and GNAME49027(G49027,G47978,G47958);
  or GNAME49028(G49028,G49027,G49026,G49025);
  xor GNAME49038(G49038,G49039,G49058);
  xor GNAME49039(G49039,G48053,G47973);
  and GNAME49040(G49040,G48053,G49058);
  and GNAME49041(G49041,G47973,G49058);
  and GNAME49042(G49042,G48053,G47973);
  or GNAME49043(G49043,G49042,G49041,G49040);
  xor GNAME49053(G49053,G49054,G48413);
  xor GNAME49054(G49054,G48068,G48048);
  and GNAME49055(G49055,G48068,G48413);
  and GNAME49056(G49056,G48048,G48413);
  and GNAME49057(G49057,G48068,G48048);
  or GNAME49058(G49058,G49057,G49056,G49055);
  xor GNAME49068(G49068,G49069,G49103);
  xor GNAME49069(G49069,G47633,G47478);
  and GNAME49070(G49070,G47633,G49103);
  and GNAME49071(G49071,G47478,G49103);
  and GNAME49072(G49072,G47633,G47478);
  or GNAME49073(G49073,G49072,G49071,G49070);
  xor GNAME49083(G49083,G49084,G49133);
  xor GNAME49084(G49084,G47648,G47493);
  and GNAME49085(G49085,G47648,G49133);
  and GNAME49086(G49086,G47493,G49133);
  and GNAME49087(G49087,G47648,G47493);
  or GNAME49088(G49088,G49087,G49086,G49085);
  xor GNAME49098(G49098,G49099,G49118);
  xor GNAME49099(G49099,G47663,G47628);
  and GNAME49100(G49100,G47663,G49118);
  and GNAME49101(G49101,G47628,G49118);
  and GNAME49102(G49102,G47663,G47628);
  or GNAME49103(G49103,G49102,G49101,G49100);
  xor GNAME49113(G49113,G49114,G49163);
  xor GNAME49114(G49114,G47813,G47658);
  and GNAME49115(G49115,G47813,G49163);
  and GNAME49116(G49116,G47658,G49163);
  and GNAME49117(G49117,G47813,G47658);
  or GNAME49118(G49118,G49117,G49116,G49115);
  xor GNAME49128(G49128,G49129,G49148);
  xor GNAME49129(G49129,G47678,G47643);
  and GNAME49130(G49130,G47678,G49148);
  and GNAME49131(G49131,G47643,G49148);
  and GNAME49132(G49132,G47678,G47643);
  or GNAME49133(G49133,G49132,G49131,G49130);
  xor GNAME49143(G49143,G49144,G49193);
  xor GNAME49144(G49144,G47828,G47673);
  and GNAME49145(G49145,G47828,G49193);
  and GNAME49146(G49146,G47673,G49193);
  and GNAME49147(G49147,G47828,G47673);
  or GNAME49148(G49148,G49147,G49146,G49145);
  xor GNAME49158(G49158,G49159,G49178);
  xor GNAME49159(G49159,G47843,G47808);
  and GNAME49160(G49160,G47843,G49178);
  and GNAME49161(G49161,G47808,G49178);
  and GNAME49162(G49162,G47843,G47808);
  or GNAME49163(G49163,G49162,G49161,G49160);
  xor GNAME49173(G49173,G49174,G49223);
  xor GNAME49174(G49174,G47993,G47838);
  and GNAME49175(G49175,G47993,G49223);
  and GNAME49176(G49176,G47838,G49223);
  and GNAME49177(G49177,G47993,G47838);
  or GNAME49178(G49178,G49177,G49176,G49175);
  xor GNAME49188(G49188,G49189,G49208);
  xor GNAME49189(G49189,G47858,G47823);
  and GNAME49190(G49190,G47858,G49208);
  and GNAME49191(G49191,G47823,G49208);
  and GNAME49192(G49192,G47858,G47823);
  or GNAME49193(G49193,G49192,G49191,G49190);
  xor GNAME49203(G49203,G49204,G49253);
  xor GNAME49204(G49204,G48008,G47853);
  and GNAME49205(G49205,G48008,G49253);
  and GNAME49206(G49206,G47853,G49253);
  and GNAME49207(G49207,G48008,G47853);
  or GNAME49208(G49208,G49207,G49206,G49205);
  xor GNAME49218(G49218,G49219,G49238);
  xor GNAME49219(G49219,G48023,G47988);
  and GNAME49220(G49220,G48023,G49238);
  and GNAME49221(G49221,G47988,G49238);
  and GNAME49222(G49222,G48023,G47988);
  or GNAME49223(G49223,G49222,G49221,G49220);
  xor GNAME49233(G49233,G49234,G49283);
  xor GNAME49234(G49234,G48083,G48018);
  and GNAME49235(G49235,G48083,G49283);
  and GNAME49236(G49236,G48018,G49283);
  and GNAME49237(G49237,G48083,G48018);
  or GNAME49238(G49238,G49237,G49236,G49235);
  xor GNAME49248(G49248,G49249,G49268);
  xor GNAME49249(G49249,G48038,G48003);
  and GNAME49250(G49250,G48038,G49268);
  and GNAME49251(G49251,G48003,G49268);
  and GNAME49252(G49252,G48038,G48003);
  or GNAME49253(G49253,G49252,G49251,G49250);
  xor GNAME49263(G49263,G49264,G49298);
  xor GNAME49264(G49264,G48098,G48033);
  and GNAME49265(G49265,G48098,G49298);
  and GNAME49266(G49266,G48033,G49298);
  and GNAME49267(G49267,G48098,G48033);
  or GNAME49268(G49268,G49267,G49266,G49265);
  xor GNAME49278(G49278,G49279,G48713);
  xor GNAME49279(G49279,G48113,G48078);
  and GNAME49280(G49280,G48113,G48713);
  and GNAME49281(G49281,G48078,G48713);
  and GNAME49282(G49282,G48113,G48078);
  or GNAME49283(G49283,G49282,G49281,G49280);
  xor GNAME49293(G49293,G49294,G48728);
  xor GNAME49294(G49294,G48128,G48093);
  and GNAME49295(G49295,G48128,G48728);
  and GNAME49296(G49296,G48093,G48728);
  and GNAME49297(G49297,G48128,G48093);
  or GNAME49298(G49298,G49297,G49296,G49295);
  xor GNAME49308(G49308,G49309,G49808);
  xor GNAME49309(G49309,G57069,G4384);
  and GNAME49310(G49310,G57069,G49808);
  and GNAME49311(G49311,G4384,G49808);
  and GNAME49312(G49312,G57069,G4384);
  or GNAME49313(G49313,G49312,G49311,G49310);
  xor GNAME49323(G49323,G49324,G50633);
  xor GNAME49324(G49324,G57667,G57693);
  and GNAME49325(G49325,G57667,G50633);
  and GNAME49326(G49326,G57693,G50633);
  and GNAME49327(G49327,G57667,G57693);
  or GNAME49328(G49328,G49327,G49326,G49325);
  xor GNAME49338(G49338,G49339,G50696);
  xor GNAME49339(G49339,G54898,G3634);
  and GNAME49340(G49340,G54898,G50696);
  and GNAME49341(G49341,G3634,G50696);
  and GNAME49342(G49342,G54898,G3634);
  or GNAME49343(G49343,G49342,G49341,G49340);
  xor GNAME49353(G49353,G49354,G50695);
  xor GNAME49354(G49354,G54924,G54937);
  and GNAME49355(G49355,G54924,G50695);
  and GNAME49356(G49356,G54937,G50695);
  and GNAME49357(G49357,G54924,G54937);
  or GNAME49358(G49358,G49357,G49356,G49355);
  xor GNAME49368(G49368,G49369,G50694);
  xor GNAME49369(G49369,G50978,G50981);
  and GNAME49370(G49370,G50978,G50694);
  and GNAME49371(G49371,G50981,G50694);
  and GNAME49372(G49372,G50978,G50981);
  or GNAME49373(G49373,G49372,G49371,G49370);
  xor GNAME49383(G49383,G49384,G49343);
  xor GNAME49384(G49384,G54911,G3655);
  and GNAME49385(G49385,G54911,G49343);
  and GNAME49386(G49386,G3655,G49343);
  and GNAME49387(G49387,G54911,G3655);
  or GNAME49388(G49388,G49387,G49386,G49385);
  xor GNAME49398(G49398,G49399,G49388);
  xor GNAME49399(G49399,G55002,G3676);
  and GNAME49400(G49400,G55002,G49388);
  and GNAME49401(G49401,G3676,G49388);
  and GNAME49402(G49402,G55002,G3676);
  or GNAME49403(G49403,G49402,G49401,G49400);
  xor GNAME49413(G49413,G49414,G49403);
  xor GNAME49414(G49414,G55015,G3697);
  and GNAME49415(G49415,G55015,G49403);
  and GNAME49416(G49416,G3697,G49403);
  and GNAME49417(G49417,G55015,G3697);
  or GNAME49418(G49418,G49417,G49416,G49415);
  xor GNAME49428(G49428,G49429,G49418);
  xor GNAME49429(G49429,G55132,G3718);
  and GNAME49430(G49430,G55132,G49418);
  and GNAME49431(G49431,G3718,G49418);
  and GNAME49432(G49432,G55132,G3718);
  or GNAME49433(G49433,G49432,G49431,G49430);
  xor GNAME49443(G49443,G49444,G49433);
  xor GNAME49444(G49444,G55145,G3739);
  and GNAME49445(G49445,G55145,G49433);
  and GNAME49446(G49446,G3739,G49433);
  and GNAME49447(G49447,G55145,G3739);
  or GNAME49448(G49448,G49447,G49446,G49445);
  xor GNAME49458(G49458,G49459,G49448);
  xor GNAME49459(G49459,G55262,G3760);
  and GNAME49460(G49460,G55262,G49448);
  and GNAME49461(G49461,G3760,G49448);
  and GNAME49462(G49462,G55262,G3760);
  or GNAME49463(G49463,G49462,G49461,G49460);
  xor GNAME49473(G49473,G49474,G49463);
  xor GNAME49474(G49474,G55275,G3821);
  and GNAME49475(G49475,G55275,G49463);
  and GNAME49476(G49476,G3821,G49463);
  and GNAME49477(G49477,G55275,G3821);
  or GNAME49478(G49478,G49477,G49476,G49475);
  xor GNAME49488(G49488,G49489,G49478);
  xor GNAME49489(G49489,G55392,G3842);
  and GNAME49490(G49490,G55392,G49478);
  and GNAME49491(G49491,G3842,G49478);
  and GNAME49492(G49492,G55392,G3842);
  or GNAME49493(G49493,G49492,G49491,G49490);
  xor GNAME49503(G49503,G49504,G49493);
  xor GNAME49504(G49504,G55405,G3863);
  and GNAME49505(G49505,G55405,G49493);
  and GNAME49506(G49506,G3863,G49493);
  and GNAME49507(G49507,G55405,G3863);
  or GNAME49508(G49508,G49507,G49506,G49505);
  xor GNAME49518(G49518,G49519,G49508);
  xor GNAME49519(G49519,G55522,G3884);
  and GNAME49520(G49520,G55522,G49508);
  and GNAME49521(G49521,G3884,G49508);
  and GNAME49522(G49522,G55522,G3884);
  or GNAME49523(G49523,G49522,G49521,G49520);
  xor GNAME49533(G49533,G49534,G49523);
  xor GNAME49534(G49534,G55535,G3905);
  and GNAME49535(G49535,G55535,G49523);
  and GNAME49536(G49536,G3905,G49523);
  and GNAME49537(G49537,G55535,G3905);
  or GNAME49538(G49538,G49537,G49536,G49535);
  xor GNAME49548(G49548,G49549,G49538);
  xor GNAME49549(G49549,G55652,G3926);
  and GNAME49550(G49550,G55652,G49538);
  and GNAME49551(G49551,G3926,G49538);
  and GNAME49552(G49552,G55652,G3926);
  or GNAME49553(G49553,G49552,G49551,G49550);
  xor GNAME49563(G49563,G49564,G49553);
  xor GNAME49564(G49564,G55665,G3947);
  and GNAME49565(G49565,G55665,G49553);
  and GNAME49566(G49566,G3947,G49553);
  and GNAME49567(G49567,G55665,G3947);
  or GNAME49568(G49568,G49567,G49566,G49565);
  xor GNAME49578(G49578,G49579,G49568);
  xor GNAME49579(G49579,G55782,G3968);
  and GNAME49580(G49580,G55782,G49568);
  and GNAME49581(G49581,G3968,G49568);
  and GNAME49582(G49582,G55782,G3968);
  or GNAME49583(G49583,G49582,G49581,G49580);
  xor GNAME49593(G49593,G49594,G49583);
  xor GNAME49594(G49594,G55795,G4029);
  and GNAME49595(G49595,G55795,G49583);
  and GNAME49596(G49596,G4029,G49583);
  and GNAME49597(G49597,G55795,G4029);
  or GNAME49598(G49598,G49597,G49596,G49595);
  xor GNAME49608(G49608,G49609,G49598);
  xor GNAME49609(G49609,G55912,G4050);
  and GNAME49610(G49610,G55912,G49598);
  and GNAME49611(G49611,G4050,G49598);
  and GNAME49612(G49612,G55912,G4050);
  or GNAME49613(G49613,G49612,G49611,G49610);
  xor GNAME49623(G49623,G49624,G49613);
  xor GNAME49624(G49624,G55925,G4071);
  and GNAME49625(G49625,G55925,G49613);
  and GNAME49626(G49626,G4071,G49613);
  and GNAME49627(G49627,G55925,G4071);
  or GNAME49628(G49628,G49627,G49626,G49625);
  xor GNAME49638(G49638,G49639,G49628);
  xor GNAME49639(G49639,G56107,G4092);
  and GNAME49640(G49640,G56107,G49628);
  and GNAME49641(G49641,G4092,G49628);
  and GNAME49642(G49642,G56107,G4092);
  or GNAME49643(G49643,G49642,G49641,G49640);
  xor GNAME49653(G49653,G49654,G49643);
  xor GNAME49654(G49654,G56120,G4113);
  and GNAME49655(G49655,G56120,G49643);
  and GNAME49656(G49656,G4113,G49643);
  and GNAME49657(G49657,G56120,G4113);
  or GNAME49658(G49658,G49657,G49656,G49655);
  xor GNAME49668(G49668,G49669,G49658);
  xor GNAME49669(G49669,G56289,G4134);
  and GNAME49670(G49670,G56289,G49658);
  and GNAME49671(G49671,G4134,G49658);
  and GNAME49672(G49672,G56289,G4134);
  or GNAME49673(G49673,G49672,G49671,G49670);
  xor GNAME49683(G49683,G49684,G49673);
  xor GNAME49684(G49684,G56302,G4155);
  and GNAME49685(G49685,G56302,G49673);
  and GNAME49686(G49686,G4155,G49673);
  and GNAME49687(G49687,G56302,G4155);
  or GNAME49688(G49688,G49687,G49686,G49685);
  xor GNAME49698(G49698,G49699,G49688);
  xor GNAME49699(G49699,G56315,G4176);
  and GNAME49700(G49700,G56315,G49688);
  and GNAME49701(G49701,G4176,G49688);
  and GNAME49702(G49702,G56315,G4176);
  or GNAME49703(G49703,G49702,G49701,G49700);
  xor GNAME49713(G49713,G49714,G49703);
  xor GNAME49714(G49714,G56497,G4237);
  and GNAME49715(G49715,G56497,G49703);
  and GNAME49716(G49716,G4237,G49703);
  and GNAME49717(G49717,G56497,G4237);
  or GNAME49718(G49718,G49717,G49716,G49715);
  xor GNAME49728(G49728,G49729,G49718);
  xor GNAME49729(G49729,G56510,G4258);
  and GNAME49730(G49730,G56510,G49718);
  and GNAME49731(G49731,G4258,G49718);
  and GNAME49732(G49732,G56510,G4258);
  or GNAME49733(G49733,G49732,G49731,G49730);
  xor GNAME49743(G49743,G49744,G49733);
  xor GNAME49744(G49744,G56679,G4279);
  and GNAME49745(G49745,G56679,G49733);
  and GNAME49746(G49746,G4279,G49733);
  and GNAME49747(G49747,G56679,G4279);
  or GNAME49748(G49748,G49747,G49746,G49745);
  xor GNAME49758(G49758,G49759,G49748);
  xor GNAME49759(G49759,G56692,G4300);
  and GNAME49760(G49760,G56692,G49748);
  and GNAME49761(G49761,G4300,G49748);
  and GNAME49762(G49762,G56692,G4300);
  or GNAME49763(G49763,G49762,G49761,G49760);
  xor GNAME49773(G49773,G49774,G49763);
  xor GNAME49774(G49774,G56874,G4321);
  and GNAME49775(G49775,G56874,G49763);
  and GNAME49776(G49776,G4321,G49763);
  and GNAME49777(G49777,G56874,G4321);
  or GNAME49778(G49778,G49777,G49776,G49775);
  xor GNAME49788(G49788,G49789,G49778);
  xor GNAME49789(G49789,G56887,G4342);
  and GNAME49790(G49790,G56887,G49778);
  and GNAME49791(G49791,G4342,G49778);
  and GNAME49792(G49792,G56887,G4342);
  or GNAME49793(G49793,G49792,G49791,G49790);
  xor GNAME49803(G49803,G49804,G49793);
  xor GNAME49804(G49804,G57056,G4363);
  and GNAME49805(G49805,G57056,G49793);
  and GNAME49806(G49806,G4363,G49793);
  and GNAME49807(G49807,G57056,G4363);
  or GNAME49808(G49808,G49807,G49806,G49805);
  xor GNAME49818(G49818,G49819,G49358);
  xor GNAME49819(G49819,G55028,G55054);
  and GNAME49820(G49820,G55028,G49358);
  and GNAME49821(G49821,G55054,G49358);
  and GNAME49822(G49822,G55028,G55054);
  or GNAME49823(G49823,G49822,G49821,G49820);
  xor GNAME49833(G49833,G49834,G49823);
  xor GNAME49834(G49834,G55041,G55067);
  and GNAME49835(G49835,G55041,G49823);
  and GNAME49836(G49836,G55067,G49823);
  and GNAME49837(G49837,G55041,G55067);
  or GNAME49838(G49838,G49837,G49836,G49835);
  xor GNAME49848(G49848,G49849,G49838);
  xor GNAME49849(G49849,G55158,G55184);
  and GNAME49850(G49850,G55158,G49838);
  and GNAME49851(G49851,G55184,G49838);
  and GNAME49852(G49852,G55158,G55184);
  or GNAME49853(G49853,G49852,G49851,G49850);
  xor GNAME49863(G49863,G49864,G49373);
  xor GNAME49864(G49864,G50972,G50975);
  and GNAME49865(G49865,G50972,G49373);
  and GNAME49866(G49866,G50975,G49373);
  and GNAME49867(G49867,G50972,G50975);
  or GNAME49868(G49868,G49867,G49866,G49865);
  xor GNAME49878(G49878,G49879,G49853);
  xor GNAME49879(G49879,G55171,G55197);
  and GNAME49880(G49880,G55171,G49853);
  and GNAME49881(G49881,G55197,G49853);
  and GNAME49882(G49882,G55171,G55197);
  or GNAME49883(G49883,G49882,G49881,G49880);
  xor GNAME49893(G49893,G49894,G49883);
  xor GNAME49894(G49894,G55288,G55314);
  and GNAME49895(G49895,G55288,G49883);
  and GNAME49896(G49896,G55314,G49883);
  and GNAME49897(G49897,G55288,G55314);
  or GNAME49898(G49898,G49897,G49896,G49895);
  xor GNAME49908(G49908,G49909,G49868);
  xor GNAME49909(G49909,G50966,G50969);
  and GNAME49910(G49910,G50966,G49868);
  and GNAME49911(G49911,G50969,G49868);
  and GNAME49912(G49912,G50966,G50969);
  or GNAME49913(G49913,G49912,G49911,G49910);
  xor GNAME49923(G49923,G49924,G49913);
  xor GNAME49924(G49924,G50960,G50963);
  and GNAME49925(G49925,G50960,G49913);
  and GNAME49926(G49926,G50963,G49913);
  and GNAME49927(G49927,G50960,G50963);
  or GNAME49928(G49928,G49927,G49926,G49925);
  xor GNAME49938(G49938,G49939,G49898);
  xor GNAME49939(G49939,G55301,G55327);
  and GNAME49940(G49940,G55301,G49898);
  and GNAME49941(G49941,G55327,G49898);
  and GNAME49942(G49942,G55301,G55327);
  or GNAME49943(G49943,G49942,G49941,G49940);
  xor GNAME49953(G49953,G49954,G49943);
  xor GNAME49954(G49954,G55418,G55444);
  and GNAME49955(G49955,G55418,G49943);
  and GNAME49956(G49956,G55444,G49943);
  and GNAME49957(G49957,G55418,G55444);
  or GNAME49958(G49958,G49957,G49956,G49955);
  xor GNAME49968(G49968,G49969,G49928);
  xor GNAME49969(G49969,G50954,G50957);
  and GNAME49970(G49970,G50954,G49928);
  and GNAME49971(G49971,G50957,G49928);
  and GNAME49972(G49972,G50954,G50957);
  or GNAME49973(G49973,G49972,G49971,G49970);
  xor GNAME49983(G49983,G49984,G49973);
  xor GNAME49984(G49984,G50948,G50951);
  and GNAME49985(G49985,G50948,G49973);
  and GNAME49986(G49986,G50951,G49973);
  and GNAME49987(G49987,G50948,G50951);
  or GNAME49988(G49988,G49987,G49986,G49985);
  xor GNAME49998(G49998,G49999,G49958);
  xor GNAME49999(G49999,G55431,G55457);
  and GNAME50000(G50000,G55431,G49958);
  and GNAME50001(G50001,G55457,G49958);
  and GNAME50002(G50002,G55431,G55457);
  or GNAME50003(G50003,G50002,G50001,G50000);
  xor GNAME50013(G50013,G50014,G50003);
  xor GNAME50014(G50014,G55548,G55574);
  and GNAME50015(G50015,G55548,G50003);
  and GNAME50016(G50016,G55574,G50003);
  and GNAME50017(G50017,G55548,G55574);
  or GNAME50018(G50018,G50017,G50016,G50015);
  xor GNAME50028(G50028,G50029,G49988);
  xor GNAME50029(G50029,G50942,G50945);
  and GNAME50030(G50030,G50942,G49988);
  and GNAME50031(G50031,G50945,G49988);
  and GNAME50032(G50032,G50942,G50945);
  or GNAME50033(G50033,G50032,G50031,G50030);
  xor GNAME50043(G50043,G50044,G50033);
  xor GNAME50044(G50044,G50936,G50939);
  and GNAME50045(G50045,G50936,G50033);
  and GNAME50046(G50046,G50939,G50033);
  and GNAME50047(G50047,G50936,G50939);
  or GNAME50048(G50048,G50047,G50046,G50045);
  xor GNAME50058(G50058,G50059,G50048);
  xor GNAME50059(G50059,G50930,G50933);
  and GNAME50060(G50060,G50930,G50048);
  and GNAME50061(G50061,G50933,G50048);
  and GNAME50062(G50062,G50930,G50933);
  or GNAME50063(G50063,G50062,G50061,G50060);
  xor GNAME50073(G50073,G50074,G50018);
  xor GNAME50074(G50074,G55561,G55587);
  and GNAME50075(G50075,G55561,G50018);
  and GNAME50076(G50076,G55587,G50018);
  and GNAME50077(G50077,G55561,G55587);
  or GNAME50078(G50078,G50077,G50076,G50075);
  xor GNAME50088(G50088,G50089,G50078);
  xor GNAME50089(G50089,G55678,G55704);
  and GNAME50090(G50090,G55678,G50078);
  and GNAME50091(G50091,G55704,G50078);
  and GNAME50092(G50092,G55678,G55704);
  or GNAME50093(G50093,G50092,G50091,G50090);
  xor GNAME50103(G50103,G50104,G50063);
  xor GNAME50104(G50104,G50924,G50927);
  and GNAME50105(G50105,G50924,G50063);
  and GNAME50106(G50106,G50927,G50063);
  and GNAME50107(G50107,G50924,G50927);
  or GNAME50108(G50108,G50107,G50106,G50105);
  xor GNAME50118(G50118,G50119,G50108);
  xor GNAME50119(G50119,G50918,G50921);
  and GNAME50120(G50120,G50918,G50108);
  and GNAME50121(G50121,G50921,G50108);
  and GNAME50122(G50122,G50918,G50921);
  or GNAME50123(G50123,G50122,G50121,G50120);
  xor GNAME50133(G50133,G50134,G50093);
  xor GNAME50134(G50134,G55691,G55717);
  and GNAME50135(G50135,G55691,G50093);
  and GNAME50136(G50136,G55717,G50093);
  and GNAME50137(G50137,G55691,G55717);
  or GNAME50138(G50138,G50137,G50136,G50135);
  xor GNAME50148(G50148,G50149,G50138);
  xor GNAME50149(G50149,G55808,G55834);
  and GNAME50150(G50150,G55808,G50138);
  and GNAME50151(G50151,G55834,G50138);
  and GNAME50152(G50152,G55808,G55834);
  or GNAME50153(G50153,G50152,G50151,G50150);
  xor GNAME50163(G50163,G50164,G50123);
  xor GNAME50164(G50164,G50912,G50915);
  and GNAME50165(G50165,G50912,G50123);
  and GNAME50166(G50166,G50915,G50123);
  and GNAME50167(G50167,G50912,G50915);
  or GNAME50168(G50168,G50167,G50166,G50165);
  xor GNAME50178(G50178,G50179,G50168);
  xor GNAME50179(G50179,G50906,G50909);
  and GNAME50180(G50180,G50906,G50168);
  and GNAME50181(G50181,G50909,G50168);
  and GNAME50182(G50182,G50906,G50909);
  or GNAME50183(G50183,G50182,G50181,G50180);
  xor GNAME50193(G50193,G50194,G50153);
  xor GNAME50194(G50194,G55821,G55847);
  and GNAME50195(G50195,G55821,G50153);
  and GNAME50196(G50196,G55847,G50153);
  and GNAME50197(G50197,G55821,G55847);
  or GNAME50198(G50198,G50197,G50196,G50195);
  xor GNAME50208(G50208,G50209,G50198);
  xor GNAME50209(G50209,G55938,G55964);
  and GNAME50210(G50210,G55938,G50198);
  and GNAME50211(G50211,G55964,G50198);
  and GNAME50212(G50212,G55938,G55964);
  or GNAME50213(G50213,G50212,G50211,G50210);
  xor GNAME50223(G50223,G50224,G50183);
  xor GNAME50224(G50224,G50900,G50903);
  and GNAME50225(G50225,G50900,G50183);
  and GNAME50226(G50226,G50903,G50183);
  and GNAME50227(G50227,G50900,G50903);
  or GNAME50228(G50228,G50227,G50226,G50225);
  xor GNAME50238(G50238,G50239,G50228);
  xor GNAME50239(G50239,G50894,G50897);
  and GNAME50240(G50240,G50894,G50228);
  and GNAME50241(G50241,G50897,G50228);
  and GNAME50242(G50242,G50894,G50897);
  or GNAME50243(G50243,G50242,G50241,G50240);
  xor GNAME50253(G50253,G50254,G50213);
  xor GNAME50254(G50254,G55951,G55977);
  and GNAME50255(G50255,G55951,G50213);
  and GNAME50256(G50256,G55977,G50213);
  and GNAME50257(G50257,G55951,G55977);
  or GNAME50258(G50258,G50257,G50256,G50255);
  xor GNAME50268(G50268,G50269,G50258);
  xor GNAME50269(G50269,G56133,G56159);
  and GNAME50270(G50270,G56133,G50258);
  and GNAME50271(G50271,G56159,G50258);
  and GNAME50272(G50272,G56133,G56159);
  or GNAME50273(G50273,G50272,G50271,G50270);
  xor GNAME50283(G50283,G50284,G50243);
  xor GNAME50284(G50284,G50888,G50891);
  and GNAME50285(G50285,G50888,G50243);
  and GNAME50286(G50286,G50891,G50243);
  and GNAME50287(G50287,G50888,G50891);
  or GNAME50288(G50288,G50287,G50286,G50285);
  xor GNAME50298(G50298,G50299,G50288);
  xor GNAME50299(G50299,G50882,G50885);
  and GNAME50300(G50300,G50882,G50288);
  and GNAME50301(G50301,G50885,G50288);
  and GNAME50302(G50302,G50882,G50885);
  or GNAME50303(G50303,G50302,G50301,G50300);
  xor GNAME50313(G50313,G50314,G50273);
  xor GNAME50314(G50314,G56146,G56172);
  and GNAME50315(G50315,G56146,G50273);
  and GNAME50316(G50316,G56172,G50273);
  and GNAME50317(G50317,G56146,G56172);
  or GNAME50318(G50318,G50317,G50316,G50315);
  xor GNAME50328(G50328,G50329,G50318);
  xor GNAME50329(G50329,G56328,G56354);
  and GNAME50330(G50330,G56328,G50318);
  and GNAME50331(G50331,G56354,G50318);
  and GNAME50332(G50332,G56328,G56354);
  or GNAME50333(G50333,G50332,G50331,G50330);
  xor GNAME50343(G50343,G50344,G50333);
  xor GNAME50344(G50344,G56341,G56367);
  and GNAME50345(G50345,G56341,G50333);
  and GNAME50346(G50346,G56367,G50333);
  and GNAME50347(G50347,G56341,G56367);
  or GNAME50348(G50348,G50347,G50346,G50345);
  xor GNAME50358(G50358,G50359,G50303);
  xor GNAME50359(G50359,G50876,G50879);
  and GNAME50360(G50360,G50876,G50303);
  and GNAME50361(G50361,G50879,G50303);
  and GNAME50362(G50362,G50876,G50879);
  or GNAME50363(G50363,G50362,G50361,G50360);
  xor GNAME50373(G50373,G50374,G50363);
  xor GNAME50374(G50374,G50870,G50873);
  and GNAME50375(G50375,G50870,G50363);
  and GNAME50376(G50376,G50873,G50363);
  and GNAME50377(G50377,G50870,G50873);
  or GNAME50378(G50378,G50377,G50376,G50375);
  xor GNAME50388(G50388,G50389,G50348);
  xor GNAME50389(G50389,G56523,G56549);
  and GNAME50390(G50390,G56523,G50348);
  and GNAME50391(G50391,G56549,G50348);
  and GNAME50392(G50392,G56523,G56549);
  or GNAME50393(G50393,G50392,G50391,G50390);
  xor GNAME50403(G50403,G50404,G50393);
  xor GNAME50404(G50404,G56536,G56562);
  and GNAME50405(G50405,G56536,G50393);
  and GNAME50406(G50406,G56562,G50393);
  and GNAME50407(G50407,G56536,G56562);
  or GNAME50408(G50408,G50407,G50406,G50405);
  xor GNAME50418(G50418,G50419,G50378);
  xor GNAME50419(G50419,G50864,G50867);
  and GNAME50420(G50420,G50864,G50378);
  and GNAME50421(G50421,G50867,G50378);
  and GNAME50422(G50422,G50864,G50867);
  or GNAME50423(G50423,G50422,G50421,G50420);
  xor GNAME50433(G50433,G50434,G50423);
  xor GNAME50434(G50434,G50858,G50861);
  and GNAME50435(G50435,G50858,G50423);
  and GNAME50436(G50436,G50861,G50423);
  and GNAME50437(G50437,G50858,G50861);
  or GNAME50438(G50438,G50437,G50436,G50435);
  xor GNAME50448(G50448,G50449,G50408);
  xor GNAME50449(G50449,G56705,G56731);
  and GNAME50450(G50450,G56705,G50408);
  and GNAME50451(G50451,G56731,G50408);
  and GNAME50452(G50452,G56705,G56731);
  or GNAME50453(G50453,G50452,G50451,G50450);
  xor GNAME50463(G50463,G50464,G50453);
  xor GNAME50464(G50464,G56718,G56744);
  and GNAME50465(G50465,G56718,G50453);
  and GNAME50466(G50466,G56744,G50453);
  and GNAME50467(G50467,G56718,G56744);
  or GNAME50468(G50468,G50467,G50466,G50465);
  xor GNAME50478(G50478,G50479,G50438);
  xor GNAME50479(G50479,G50852,G50855);
  and GNAME50480(G50480,G50852,G50438);
  and GNAME50481(G50481,G50855,G50438);
  and GNAME50482(G50482,G50852,G50855);
  or GNAME50483(G50483,G50482,G50481,G50480);
  xor GNAME50493(G50493,G50494,G50483);
  xor GNAME50494(G50494,G50846,G50849);
  and GNAME50495(G50495,G50846,G50483);
  and GNAME50496(G50496,G50849,G50483);
  and GNAME50497(G50497,G50846,G50849);
  or GNAME50498(G50498,G50497,G50496,G50495);
  xor GNAME50508(G50508,G50509,G50468);
  xor GNAME50509(G50509,G56900,G56926);
  and GNAME50510(G50510,G56900,G50468);
  and GNAME50511(G50511,G56926,G50468);
  and GNAME50512(G50512,G56900,G56926);
  or GNAME50513(G50513,G50512,G50511,G50510);
  xor GNAME50523(G50523,G50524,G50513);
  xor GNAME50524(G50524,G56913,G56939);
  and GNAME50525(G50525,G56913,G50513);
  and GNAME50526(G50526,G56939,G50513);
  and GNAME50527(G50527,G56913,G56939);
  or GNAME50528(G50528,G50527,G50526,G50525);
  xor GNAME50538(G50538,G50539,G50498);
  xor GNAME50539(G50539,G50840,G50843);
  and GNAME50540(G50540,G50840,G50498);
  and GNAME50541(G50541,G50843,G50498);
  and GNAME50542(G50542,G50840,G50843);
  or GNAME50543(G50543,G50542,G50541,G50540);
  xor GNAME50553(G50553,G50554,G50543);
  xor GNAME50554(G50554,G50834,G50837);
  and GNAME50555(G50555,G50834,G50543);
  and GNAME50556(G50556,G50837,G50543);
  and GNAME50557(G50557,G50834,G50837);
  or GNAME50558(G50558,G50557,G50556,G50555);
  xor GNAME50568(G50568,G50569,G50528);
  xor GNAME50569(G50569,G57082,G57108);
  and GNAME50570(G50570,G57082,G50528);
  and GNAME50571(G50571,G57108,G50528);
  and GNAME50572(G50572,G57082,G57108);
  or GNAME50573(G50573,G50572,G50571,G50570);
  xor GNAME50583(G50583,G50584,G50573);
  xor GNAME50584(G50584,G57095,G57121);
  and GNAME50585(G50585,G57095,G50573);
  and GNAME50586(G50586,G57121,G50573);
  and GNAME50587(G50587,G57095,G57121);
  or GNAME50588(G50588,G50587,G50586,G50585);
  xor GNAME50598(G50598,G50599,G50558);
  xor GNAME50599(G50599,G50828,G50831);
  and GNAME50600(G50600,G50828,G50558);
  and GNAME50601(G50601,G50831,G50558);
  and GNAME50602(G50602,G50828,G50831);
  or GNAME50603(G50603,G50602,G50601,G50600);
  xor GNAME50613(G50613,G50614,G50603);
  xor GNAME50614(G50614,G50822,G50825);
  and GNAME50615(G50615,G50822,G50603);
  and GNAME50616(G50616,G50825,G50603);
  and GNAME50617(G50617,G50822,G50825);
  or GNAME50618(G50618,G50617,G50616,G50615);
  xor GNAME50628(G50628,G50629,G50588);
  xor GNAME50629(G50629,G57654,G57680);
  and GNAME50630(G50630,G57654,G50588);
  and GNAME50631(G50631,G57680,G50588);
  and GNAME50632(G50632,G57654,G57680);
  or GNAME50633(G50633,G50632,G50631,G50630);
  xor GNAME50643(G50643,G50644,G50618);
  xor GNAME50644(G50644,G50816,G50819);
  and GNAME50645(G50645,G50816,G50618);
  and GNAME50646(G50646,G50819,G50618);
  and GNAME50647(G50647,G50816,G50819);
  or GNAME50648(G50648,G50647,G50646,G50645);
  xor GNAME50658(G50658,G50659,G50648);
  xor GNAME50659(G50659,G50810,G50813);
  and GNAME50660(G50660,G50810,G50648);
  and GNAME50661(G50661,G50813,G50648);
  and GNAME50662(G50662,G50810,G50813);
  or GNAME50663(G50663,G50662,G50661,G50660);
  xor GNAME50673(G50673,G50674,G50663);
  xor GNAME50674(G50674,G50804,G50807);
  and GNAME50675(G50675,G50804,G50663);
  and GNAME50676(G50676,G50807,G50663);
  and GNAME50677(G50677,G50804,G50807);
  or GNAME50678(G50678,G50677,G50676,G50675);
  xor GNAME50688(G50688,G50689,G50678);
  xor GNAME50689(G50689,G50798,G50801);
  and GNAME50690(G50690,G50798,G50678);
  and GNAME50691(G50691,G50801,G50678);
  and GNAME50692(G50692,G50798,G50801);
  or GNAME50693(G50693,G50692,G50691,G50690);
  and GNAME50694(G50694,G50987,G50984);
  and GNAME50695(G50695,G54807,G54833);
  and GNAME50696(G50696,G3613,G54820);
  and GNAME50697(G50697,G53071,G53080);
  and GNAME50698(G50698,G53074,G53083);
  and GNAME50699(G50699,G53077,G53086);
  and GNAME50700(G50700,G51745,G57723);
  and GNAME50701(G50701,G56068,G54569);
  or GNAME50702(G50702,G50701,G50700);
  and GNAME50703(G50703,G51739,G57723);
  and GNAME50704(G50704,G56055,G54569);
  or GNAME50705(G50705,G50704,G50703);
  and GNAME50706(G50706,G51733,G57723);
  and GNAME50707(G50707,G56042,G54569);
  or GNAME50708(G50708,G50707,G50706);
  and GNAME50709(G50709,G51721,G57723);
  and GNAME50710(G50710,G56029,G54569);
  or GNAME50711(G50711,G50710,G50709);
  and GNAME50712(G50712,G54563,G57723);
  and GNAME50713(G50713,G55990,G54569);
  or GNAME50714(G50714,G50713,G50712);
  and GNAME50715(G50715,G51763,G57723);
  and GNAME50716(G50716,G56237,G54569);
  or GNAME50717(G50717,G50716,G50715);
  and GNAME50718(G50718,G51757,G57723);
  and GNAME50719(G50719,G56224,G54569);
  or GNAME50720(G50720,G50719,G50718);
  and GNAME50721(G50721,G51751,G57723);
  and GNAME50722(G50722,G56211,G54569);
  or GNAME50723(G50723,G50722,G50721);
  and GNAME50724(G50724,G51769,G57724);
  and GNAME50725(G50725,G56250,G54569);
  or GNAME50726(G50726,G50725,G50724);
  and GNAME50727(G50727,G57724,G51775);
  and GNAME50728(G50728,G56406,G54569);
  or GNAME50729(G50729,G50728,G50727);
  and GNAME50730(G50730,G51799,G57723);
  and GNAME50731(G50731,G56458,G54569);
  or GNAME50732(G50732,G50731,G50730);
  and GNAME50733(G50733,G51793,G57723);
  and GNAME50734(G50734,G56445,G54569);
  or GNAME50735(G50735,G50734,G50733);
  and GNAME50736(G50736,G51787,G57723);
  and GNAME50737(G50737,G56432,G54569);
  or GNAME50738(G50738,G50737,G50736);
  and GNAME50739(G50739,G51781,G57723);
  and GNAME50740(G50740,G56419,G54569);
  or GNAME50741(G50741,G50740,G50739);
  and GNAME50742(G50742,G51829,G57723);
  and GNAME50743(G50743,G56783,G54569);
  or GNAME50744(G50744,G50743,G50742);
  and GNAME50745(G50745,G51823,G57723);
  and GNAME50746(G50746,G56640,G54569);
  or GNAME50747(G50747,G50746,G50745);
  and GNAME50748(G50748,G51817,G57723);
  and GNAME50749(G50749,G56627,G54569);
  or GNAME50750(G50750,G50749,G50748);
  and GNAME50751(G50751,G51811,G57723);
  and GNAME50752(G50752,G56614,G54569);
  or GNAME50753(G50753,G50752,G50751);
  and GNAME50754(G50754,G51805,G57723);
  and GNAME50755(G50755,G56601,G54569);
  or GNAME50756(G50756,G50755,G50754);
  and GNAME50757(G50757,G51853,G57723);
  and GNAME50758(G50758,G56835,G54569);
  or GNAME50759(G50759,G50758,G50757);
  and GNAME50760(G50760,G51847,G57723);
  and GNAME50761(G50761,G56822,G54569);
  or GNAME50762(G50762,G50761,G50760);
  and GNAME50763(G50763,G51841,G57723);
  and GNAME50764(G50764,G56809,G54569);
  or GNAME50765(G50765,G50764,G50763);
  and GNAME50766(G50766,G51835,G57723);
  and GNAME50767(G50767,G56796,G54569);
  or GNAME50768(G50768,G50767,G50766);
  and GNAME50769(G50769,G51883,G57723);
  and GNAME50770(G50770,G57602,G54569);
  or GNAME50771(G50771,G50770,G50769);
  and GNAME50772(G50772,G51877,G57723);
  and GNAME50773(G50773,G57017,G54569);
  or GNAME50774(G50774,G50773,G50772);
  and GNAME50775(G50775,G51871,G57723);
  and GNAME50776(G50776,G57004,G54569);
  or GNAME50777(G50777,G50776,G50775);
  and GNAME50778(G50778,G51865,G57723);
  and GNAME50779(G50779,G56991,G54569);
  or GNAME50780(G50780,G50779,G50778);
  and GNAME50781(G50781,G51859,G57723);
  and GNAME50782(G50782,G56978,G54569);
  or GNAME50783(G50783,G50782,G50781);
  and GNAME50784(G50784,G54711,G57723);
  and GNAME50785(G50785,G57576,G54569);
  or GNAME50786(G50786,G50785,G50784);
  and GNAME50787(G50787,G51727,G57723);
  and GNAME50788(G50788,G57641,G54569);
  or GNAME50789(G50789,G50788,G50787);
  and GNAME50790(G50790,G51895,G57723);
  and GNAME50791(G50791,G57628,G54569);
  or GNAME50792(G50792,G50791,G50790);
  and GNAME50793(G50793,G51889,G57723);
  and GNAME50794(G50794,G57615,G54569);
  or GNAME50795(G50795,G50794,G50793);
  and GNAME50796(G50796,G54712,G57780);
  and GNAME50797(G50797,G57563,G54646);
  or GNAME50798(G50798,G50797,G50796);
  and GNAME50799(G50799,G54713,G57779);
  and GNAME50800(G50800,G57589,G54645);
  or GNAME50801(G50801,G50800,G50799);
  and GNAME50802(G50802,G51709,G57780);
  and GNAME50803(G50803,G56965,G54646);
  or GNAME50804(G50804,G50803,G50802);
  and GNAME50805(G50805,G51715,G57779);
  and GNAME50806(G50806,G57043,G54645);
  or GNAME50807(G50807,G50806,G50805);
  and GNAME50808(G50808,G51697,G57780);
  and GNAME50809(G50809,G56952,G54646);
  or GNAME50810(G50810,G50809,G50808);
  and GNAME50811(G50811,G51703,G57779);
  and GNAME50812(G50812,G57030,G54645);
  or GNAME50813(G50813,G50812,G50811);
  and GNAME50814(G50814,G51685,G57780);
  and GNAME50815(G50815,G56770,G54646);
  or GNAME50816(G50816,G50815,G50814);
  and GNAME50817(G50817,G51691,G57779);
  and GNAME50818(G50818,G56861,G54645);
  or GNAME50819(G50819,G50818,G50817);
  and GNAME50820(G50820,G51673,G57780);
  and GNAME50821(G50821,G56757,G54646);
  or GNAME50822(G50822,G50821,G50820);
  and GNAME50823(G50823,G51679,G57779);
  and GNAME50824(G50824,G56848,G54645);
  or GNAME50825(G50825,G50824,G50823);
  and GNAME50826(G50826,G51661,G57780);
  and GNAME50827(G50827,G56588,G54646);
  or GNAME50828(G50828,G50827,G50826);
  and GNAME50829(G50829,G51667,G57779);
  and GNAME50830(G50830,G56666,G54645);
  or GNAME50831(G50831,G50830,G50829);
  and GNAME50832(G50832,G51649,G57780);
  and GNAME50833(G50833,G56575,G54646);
  or GNAME50834(G50834,G50833,G50832);
  and GNAME50835(G50835,G51655,G57779);
  and GNAME50836(G50836,G56653,G54645);
  or GNAME50837(G50837,G50836,G50835);
  and GNAME50838(G50838,G51637,G57780);
  and GNAME50839(G50839,G56393,G54646);
  or GNAME50840(G50840,G50839,G50838);
  and GNAME50841(G50841,G51643,G57779);
  and GNAME50842(G50842,G56484,G54645);
  or GNAME50843(G50843,G50842,G50841);
  and GNAME50844(G50844,G51625,G57780);
  and GNAME50845(G50845,G56380,G54646);
  or GNAME50846(G50846,G50845,G50844);
  and GNAME50847(G50847,G51631,G57779);
  and GNAME50848(G50848,G56471,G54645);
  or GNAME50849(G50849,G50848,G50847);
  and GNAME50850(G50850,G51613,G57780);
  and GNAME50851(G50851,G56198,G54646);
  or GNAME50852(G50852,G50851,G50850);
  and GNAME50853(G50853,G51619,G57779);
  and GNAME50854(G50854,G56276,G54645);
  or GNAME50855(G50855,G50854,G50853);
  and GNAME50856(G50856,G51601,G57780);
  and GNAME50857(G50857,G56185,G54646);
  or GNAME50858(G50858,G50857,G50856);
  and GNAME50859(G50859,G51607,G57779);
  and GNAME50860(G50860,G56263,G54645);
  or GNAME50861(G50861,G50860,G50859);
  and GNAME50862(G50862,G51589,G57780);
  and GNAME50863(G50863,G56016,G54646);
  or GNAME50864(G50864,G50863,G50862);
  and GNAME50865(G50865,G51595,G57779);
  and GNAME50866(G50866,G56094,G54645);
  or GNAME50867(G50867,G50866,G50865);
  and GNAME50868(G50868,G51577,G57780);
  and GNAME50869(G50869,G56003,G54646);
  or GNAME50870(G50870,G50869,G50868);
  and GNAME50871(G50871,G51583,G57779);
  and GNAME50872(G50872,G56081,G54645);
  or GNAME50873(G50873,G50872,G50871);
  and GNAME50874(G50874,G51565,G57780);
  and GNAME50875(G50875,G55873,G54646);
  or GNAME50876(G50876,G50875,G50874);
  and GNAME50877(G50877,G51571,G57779);
  and GNAME50878(G50878,G55899,G54645);
  or GNAME50879(G50879,G50878,G50877);
  and GNAME50880(G50880,G51553,G57780);
  and GNAME50881(G50881,G55860,G54646);
  or GNAME50882(G50882,G50881,G50880);
  and GNAME50883(G50883,G51559,G57779);
  and GNAME50884(G50884,G55886,G54645);
  or GNAME50885(G50885,G50884,G50883);
  and GNAME50886(G50886,G51541,G57780);
  and GNAME50887(G50887,G55743,G54646);
  or GNAME50888(G50888,G50887,G50886);
  and GNAME50889(G50889,G51547,G57779);
  and GNAME50890(G50890,G55769,G54645);
  or GNAME50891(G50891,G50890,G50889);
  and GNAME50892(G50892,G51529,G57780);
  and GNAME50893(G50893,G55730,G54646);
  or GNAME50894(G50894,G50893,G50892);
  and GNAME50895(G50895,G51535,G57779);
  and GNAME50896(G50896,G55756,G54645);
  or GNAME50897(G50897,G50896,G50895);
  and GNAME50898(G50898,G51517,G57780);
  and GNAME50899(G50899,G55613,G54646);
  or GNAME50900(G50900,G50899,G50898);
  and GNAME50901(G50901,G51523,G57779);
  and GNAME50902(G50902,G55639,G54645);
  or GNAME50903(G50903,G50902,G50901);
  and GNAME50904(G50904,G51505,G57780);
  and GNAME50905(G50905,G55600,G54646);
  or GNAME50906(G50906,G50905,G50904);
  and GNAME50907(G50907,G51511,G57779);
  and GNAME50908(G50908,G55626,G54645);
  or GNAME50909(G50909,G50908,G50907);
  and GNAME50910(G50910,G51493,G57780);
  and GNAME50911(G50911,G55483,G54646);
  or GNAME50912(G50912,G50911,G50910);
  and GNAME50913(G50913,G51499,G57779);
  and GNAME50914(G50914,G55509,G54645);
  or GNAME50915(G50915,G50914,G50913);
  and GNAME50916(G50916,G51469,G57780);
  and GNAME50917(G50917,G55470,G54646);
  or GNAME50918(G50918,G50917,G50916);
  and GNAME50919(G50919,G51475,G57779);
  and GNAME50920(G50920,G55496,G54645);
  or GNAME50921(G50921,G50920,G50919);
  and GNAME50922(G50922,G51457,G57780);
  and GNAME50923(G50923,G55353,G54646);
  or GNAME50924(G50924,G50923,G50922);
  and GNAME50925(G50925,G51463,G57779);
  and GNAME50926(G50926,G55379,G54645);
  or GNAME50927(G50927,G50926,G50925);
  and GNAME50928(G50928,G57788,G51481);
  and GNAME50929(G50929,G55340,G54646);
  or GNAME50930(G50930,G50929,G50928);
  and GNAME50931(G50931,G57787,G51487);
  and GNAME50932(G50932,G55366,G54645);
  or GNAME50933(G50933,G50932,G50931);
  and GNAME50934(G50934,G51445,G57788);
  and GNAME50935(G50935,G55223,G54646);
  or GNAME50936(G50936,G50935,G50934);
  and GNAME50937(G50937,G51451,G57787);
  and GNAME50938(G50938,G55249,G54645);
  or GNAME50939(G50939,G50938,G50937);
  and GNAME50940(G50940,G51433,G57780);
  and GNAME50941(G50941,G55210,G54646);
  or GNAME50942(G50942,G50941,G50940);
  and GNAME50943(G50943,G51439,G57779);
  and GNAME50944(G50944,G55236,G54645);
  or GNAME50945(G50945,G50944,G50943);
  and GNAME50946(G50946,G51421,G57780);
  and GNAME50947(G50947,G55093,G54646);
  or GNAME50948(G50948,G50947,G50946);
  and GNAME50949(G50949,G51427,G57779);
  and GNAME50950(G50950,G55119,G54645);
  or GNAME50951(G50951,G50950,G50949);
  and GNAME50952(G50952,G51409,G57780);
  and GNAME50953(G50953,G55080,G54646);
  or GNAME50954(G50954,G50953,G50952);
  and GNAME50955(G50955,G51415,G57779);
  and GNAME50956(G50956,G55106,G54645);
  or GNAME50957(G50957,G50956,G50955);
  and GNAME50958(G50958,G51397,G57780);
  and GNAME50959(G50959,G54963,G54646);
  or GNAME50960(G50960,G50959,G50958);
  and GNAME50961(G50961,G51403,G57779);
  and GNAME50962(G50962,G54989,G54645);
  or GNAME50963(G50963,G50962,G50961);
  and GNAME50964(G50964,G51385,G57780);
  and GNAME50965(G50965,G54950,G54646);
  or GNAME50966(G50966,G50965,G50964);
  and GNAME50967(G50967,G51391,G57779);
  and GNAME50968(G50968,G54976,G54645);
  or GNAME50969(G50969,G50968,G50967);
  and GNAME50970(G50970,G51373,G57780);
  and GNAME50971(G50971,G54859,G54646);
  or GNAME50972(G50972,G50971,G50970);
  and GNAME50973(G50973,G51379,G57779);
  and GNAME50974(G50974,G54885,G54645);
  or GNAME50975(G50975,G50974,G50973);
  and GNAME50976(G50976,G51361,G57780);
  and GNAME50977(G50977,G54846,G54646);
  or GNAME50978(G50978,G50977,G50976);
  and GNAME50979(G50979,G51367,G57779);
  and GNAME50980(G50980,G54872,G54645);
  or GNAME50981(G50981,G50980,G50979);
  and GNAME50982(G50982,G54564,G57780);
  and GNAME50983(G50983,G54755,G54646);
  or GNAME50984(G50984,G50983,G50982);
  and GNAME50985(G50985,G54565,G57779);
  and GNAME50986(G50986,G54768,G54645);
  or GNAME50987(G50987,G50986,G50985);
  not GNAME50988(G50988,G50990);
  not GNAME50989(G50989,G57804);
  and GNAME50990(G50990,G57781,G50989);
  not GNAME50991(G50991,G50993);
  not GNAME50992(G50992,G57805);
  and GNAME50993(G50993,G57782,G50992);
  not GNAME50994(G50994,G50996);
  not GNAME50995(G50995,G57806);
  and GNAME50996(G50996,G57783,G50995);
  not GNAME50997(G50997,G50999);
  not GNAME50998(G50998,G57804);
  and GNAME50999(G50999,G57784,G50998);
  not GNAME51000(G51000,G51002);
  not GNAME51001(G51001,G57805);
  and GNAME51002(G51002,G57785,G51001);
  not GNAME51003(G51003,G51005);
  not GNAME51004(G51004,G57806);
  and GNAME51005(G51005,G57786,G51004);
  not GNAME51006(G51006,G51008);
  not GNAME51007(G51007,G57804);
  and GNAME51008(G51008,G57801,G51007);
  not GNAME51009(G51009,G51011);
  not GNAME51010(G51010,G57805);
  and GNAME51011(G51011,G57802,G51010);
  not GNAME51012(G51012,G51014);
  not GNAME51013(G51013,G57806);
  and GNAME51014(G51014,G57803,G51013);
  not GNAME51015(G51015,G51017);
  not GNAME51016(G51016,G57837);
  and GNAME51017(G51017,G57816,G51016);
  not GNAME51018(G51018,G51020);
  not GNAME51019(G51019,G57838);
  and GNAME51020(G51020,G57817,G51019);
  not GNAME51021(G51021,G51023);
  not GNAME51022(G51022,G57839);
  and GNAME51023(G51023,G57818,G51022);
  not GNAME51024(G51024,G51026);
  not GNAME51025(G51025,G57837);
  and GNAME51026(G51026,G57831,G51025);
  not GNAME51027(G51027,G51029);
  not GNAME51028(G51028,G57838);
  and GNAME51029(G51029,G57832,G51028);
  not GNAME51030(G51030,G51032);
  not GNAME51031(G51031,G57839);
  and GNAME51032(G51032,G57833,G51031);
  not GNAME51033(G51033,G51035);
  not GNAME51034(G51034,G57837);
  and GNAME51035(G51035,G57846,G51034);
  not GNAME51036(G51036,G51038);
  not GNAME51037(G51037,G57838);
  and GNAME51038(G51038,G57847,G51037);
  not GNAME51039(G51039,G51041);
  not GNAME51040(G51040,G57839);
  and GNAME51041(G51041,G57848,G51040);
  not GNAME51042(G51042,G51044);
  not GNAME51043(G51043,G57837);
  and GNAME51044(G51044,G57834,G51043);
  not GNAME51045(G51045,G51047);
  not GNAME51046(G51046,G57838);
  and GNAME51047(G51047,G57835,G51046);
  not GNAME51048(G51048,G51050);
  not GNAME51049(G51049,G57839);
  and GNAME51050(G51050,G57836,G51049);
  not GNAME51051(G51051,G51053);
  not GNAME51052(G51052,G57837);
  and GNAME51053(G51053,G57849,G51052);
  not GNAME51054(G51054,G51056);
  not GNAME51055(G51055,G57838);
  and GNAME51056(G51056,G57850,G51055);
  not GNAME51057(G51057,G51059);
  not GNAME51058(G51058,G57839);
  and GNAME51059(G51059,G57851,G51058);
  xor GNAME51060(G51060,G51061,G52048);
  xor GNAME51061(G51061,G52716,G52114);
  xor GNAME51062(G51062,G51063,G52049);
  xor GNAME51063(G51063,G52718,G52115);
  xor GNAME51064(G51064,G51065,G52050);
  xor GNAME51065(G51065,G52720,G52116);
  xor GNAME51066(G51066,G51067,G49313);
  xor GNAME51067(G51067,G57706,G4405);
  not GNAME51068(G51068,G51070);
  not GNAME51069(G51069,G57804);
  or GNAME51070(G51070,G57912,G51069);
  not GNAME51071(G51071,G51073);
  not GNAME51072(G51072,G57805);
  or GNAME51073(G51073,G57913,G51072);
  not GNAME51074(G51074,G51076);
  not GNAME51075(G51075,G57806);
  or GNAME51076(G51076,G57914,G51075);
  not GNAME51077(G51077,G51079);
  not GNAME51078(G51078,G57804);
  or GNAME51079(G51079,G57858,G51078);
  not GNAME51080(G51080,G51082);
  not GNAME51081(G51081,G57805);
  or GNAME51082(G51082,G57859,G51081);
  not GNAME51083(G51083,G51085);
  not GNAME51084(G51084,G57806);
  or GNAME51085(G51085,G57860,G51084);
  not GNAME51086(G51086,G51088);
  not GNAME51087(G51087,G49698);
  or GNAME51088(G51088,G57856,G51087);
  not GNAME51089(G51089,G51091);
  not GNAME51090(G51090,G49683);
  or GNAME51091(G51091,G57856,G51090);
  not GNAME51092(G51092,G51094);
  not GNAME51093(G51093,G49668);
  or GNAME51094(G51094,G57856,G51093);
  not GNAME51095(G51095,G51097);
  not GNAME51096(G51096,G49653);
  or GNAME51097(G51097,G57856,G51096);
  not GNAME51098(G51098,G51100);
  not GNAME51099(G51099,G49638);
  or GNAME51100(G51100,G57856,G51099);
  not GNAME51101(G51101,G51103);
  not GNAME51102(G51102,G49623);
  or GNAME51103(G51103,G57856,G51102);
  not GNAME51104(G51104,G51106);
  not GNAME51105(G51105,G49608);
  or GNAME51106(G51106,G57856,G51105);
  not GNAME51107(G51107,G51109);
  not GNAME51108(G51108,G49593);
  or GNAME51109(G51109,G57856,G51108);
  not GNAME51110(G51110,G51112);
  not GNAME51111(G51111,G49803);
  or GNAME51112(G51112,G57857,G51111);
  not GNAME51113(G51113,G51115);
  not GNAME51114(G51114,G49788);
  or GNAME51115(G51115,G57857,G51114);
  not GNAME51116(G51116,G51118);
  not GNAME51117(G51117,G49773);
  or GNAME51118(G51118,G57857,G51117);
  not GNAME51119(G51119,G51121);
  not GNAME51120(G51120,G49758);
  or GNAME51121(G51121,G57857,G51120);
  not GNAME51122(G51122,G51124);
  not GNAME51123(G51123,G49743);
  or GNAME51124(G51124,G57856,G51123);
  not GNAME51125(G51125,G51127);
  not GNAME51126(G51126,G49728);
  or GNAME51127(G51127,G57856,G51126);
  not GNAME51128(G51128,G51130);
  not GNAME51129(G51129,G49713);
  or GNAME51130(G51130,G57856,G51129);
  not GNAME51131(G51131,G51133);
  not GNAME51132(G51132,G49458);
  or GNAME51133(G51133,G57857,G51132);
  not GNAME51134(G51134,G51136);
  not GNAME51135(G51135,G49443);
  or GNAME51136(G51136,G57857,G51135);
  not GNAME51137(G51137,G51139);
  not GNAME51138(G51138,G49428);
  or GNAME51139(G51139,G57857,G51138);
  not GNAME51140(G51140,G51142);
  not GNAME51141(G51141,G49413);
  or GNAME51142(G51142,G57857,G51141);
  not GNAME51143(G51143,G51145);
  not GNAME51144(G51144,G49398);
  or GNAME51145(G51145,G57857,G51144);
  not GNAME51146(G51146,G51148);
  not GNAME51147(G51147,G49383);
  or GNAME51148(G51148,G57857,G51147);
  not GNAME51149(G51149,G51151);
  not GNAME51150(G51150,G49338);
  or GNAME51151(G51151,G57856,G51150);
  not GNAME51152(G51152,G51154);
  not GNAME51153(G51153,G49578);
  or GNAME51154(G51154,G57852,G51153);
  not GNAME51155(G51155,G51157);
  not GNAME51156(G51156,G49563);
  or GNAME51157(G51157,G57852,G51156);
  not GNAME51158(G51158,G51160);
  not GNAME51159(G51159,G49548);
  or GNAME51160(G51160,G57852,G51159);
  not GNAME51161(G51161,G51163);
  not GNAME51162(G51162,G49533);
  or GNAME51163(G51163,G57852,G51162);
  not GNAME51164(G51164,G51166);
  not GNAME51165(G51165,G49518);
  or GNAME51166(G51166,G57852,G51165);
  not GNAME51167(G51167,G51169);
  not GNAME51168(G51168,G49503);
  or GNAME51169(G51169,G57852,G51168);
  not GNAME51170(G51170,G51172);
  not GNAME51171(G51171,G49488);
  or GNAME51172(G51172,G57857,G51171);
  not GNAME51173(G51173,G51175);
  not GNAME51174(G51174,G49473);
  or GNAME51175(G51175,G57857,G51174);
  not GNAME51176(G51176,G51178);
  not GNAME51177(G51177,G57804);
  or GNAME51178(G51178,G57864,G51177);
  not GNAME51179(G51179,G51181);
  not GNAME51180(G51180,G57805);
  or GNAME51181(G51181,G57865,G51180);
  not GNAME51182(G51182,G51184);
  not GNAME51183(G51183,G57806);
  or GNAME51184(G51184,G57866,G51183);
  not GNAME51185(G51185,G51187);
  not GNAME51186(G51186,G57804);
  or GNAME51187(G51187,G57873,G51186);
  not GNAME51188(G51188,G51190);
  not GNAME51189(G51189,G57805);
  or GNAME51190(G51190,G57874,G51189);
  not GNAME51191(G51191,G51193);
  not GNAME51192(G51192,G57806);
  or GNAME51193(G51193,G57875,G51192);
  not GNAME51194(G51194,G51196);
  not GNAME51195(G51195,G57804);
  or GNAME51196(G51196,G57936,G51195);
  not GNAME51197(G51197,G51199);
  not GNAME51198(G51198,G57805);
  or GNAME51199(G51199,G57937,G51198);
  not GNAME51200(G51200,G51202);
  not GNAME51201(G51201,G57806);
  or GNAME51202(G51202,G57938,G51201);
  not GNAME51203(G51203,G51205);
  not GNAME51204(G51204,G57837);
  or GNAME51205(G51205,G57939,G51204);
  not GNAME51206(G51206,G51208);
  not GNAME51207(G51207,G57838);
  or GNAME51208(G51208,G57940,G51207);
  not GNAME51209(G51209,G51211);
  not GNAME51210(G51210,G57839);
  or GNAME51211(G51211,G57941,G51210);
  not GNAME51212(G51212,G51214);
  not GNAME51213(G51213,G57837);
  or GNAME51214(G51214,G57900,G51213);
  not GNAME51215(G51215,G51217);
  not GNAME51216(G51216,G57838);
  or GNAME51217(G51217,G57902,G51216);
  not GNAME51218(G51218,G51220);
  not GNAME51219(G51219,G57839);
  or GNAME51220(G51220,G57904,G51219);
  not GNAME51221(G51221,G51223);
  not GNAME51222(G51222,G57837);
  or GNAME51223(G51223,G57901,G51222);
  not GNAME51224(G51224,G51226);
  not GNAME51225(G51225,G57838);
  or GNAME51226(G51226,G57903,G51225);
  not GNAME51227(G51227,G51229);
  not GNAME51228(G51228,G57839);
  or GNAME51229(G51229,G57905,G51228);
  or GNAME51230(G51230,G49308,G51066);
  xor GNAME51235(G51235,G52864,G52867);
  and GNAME51236(G51236,G52864,G52867);
  xor GNAME51241(G51241,G52870,G52873);
  and GNAME51242(G51242,G52870,G52873);
  xor GNAME51247(G51247,G52876,G52879);
  and GNAME51248(G51248,G52876,G52879);
  xor GNAME51253(G51253,G52882,G52885);
  and GNAME51254(G51254,G52882,G52885);
  xor GNAME51259(G51259,G52888,G52891);
  and GNAME51260(G51260,G52888,G52891);
  xor GNAME51265(G51265,G52894,G52897);
  and GNAME51266(G51266,G52894,G52897);
  xor GNAME51271(G51271,G52918,G52921);
  and GNAME51272(G51272,G52918,G52921);
  xor GNAME51277(G51277,G52924,G52927);
  and GNAME51278(G51278,G52924,G52927);
  xor GNAME51283(G51283,G52930,G52933);
  and GNAME51284(G51284,G52930,G52933);
  xor GNAME51289(G51289,G52954,G52957);
  and GNAME51290(G51290,G52954,G52957);
  xor GNAME51295(G51295,G52960,G52963);
  and GNAME51296(G51296,G52960,G52963);
  xor GNAME51301(G51301,G52966,G52969);
  and GNAME51302(G51302,G52966,G52969);
  xor GNAME51307(G51307,G52990,G52993);
  and GNAME51308(G51308,G52990,G52993);
  xor GNAME51313(G51313,G52996,G52999);
  and GNAME51314(G51314,G52996,G52999);
  xor GNAME51319(G51319,G53002,G53005);
  and GNAME51320(G51320,G53002,G53005);
  xor GNAME51325(G51325,G53089,G54556);
  and GNAME51326(G51326,G53089,G54556);
  xor GNAME51331(G51331,G53092,G54559);
  and GNAME51332(G51332,G53092,G54559);
  xor GNAME51337(G51337,G53095,G54562);
  and GNAME51338(G51338,G53095,G54562);
  xor GNAME51343(G51343,G54538,G54541);
  and GNAME51344(G51344,G54538,G54541);
  xor GNAME51349(G51349,G54544,G54547);
  and GNAME51350(G51350,G54544,G54547);
  xor GNAME51355(G51355,G54550,G54553);
  and GNAME51356(G51356,G54550,G54553);
  xor GNAME51361(G51361,G54846,G54755);
  and GNAME51362(G51362,G54846,G54755);
  xor GNAME51367(G51367,G54872,G54768);
  and GNAME51368(G51368,G54872,G54768);
  xor GNAME51373(G51373,G54859,G51362);
  and GNAME51374(G51374,G54859,G51362);
  xor GNAME51379(G51379,G54885,G51368);
  and GNAME51380(G51380,G54885,G51368);
  xor GNAME51385(G51385,G54950,G51374);
  and GNAME51386(G51386,G54950,G51374);
  xor GNAME51391(G51391,G54976,G51380);
  and GNAME51392(G51392,G54976,G51380);
  xor GNAME51397(G51397,G54963,G51386);
  and GNAME51398(G51398,G54963,G51386);
  xor GNAME51403(G51403,G54989,G51392);
  and GNAME51404(G51404,G54989,G51392);
  xor GNAME51409(G51409,G55080,G51398);
  and GNAME51410(G51410,G55080,G51398);
  xor GNAME51415(G51415,G55106,G51404);
  and GNAME51416(G51416,G55106,G51404);
  xor GNAME51421(G51421,G55093,G51410);
  and GNAME51422(G51422,G55093,G51410);
  xor GNAME51427(G51427,G55119,G51416);
  and GNAME51428(G51428,G55119,G51416);
  xor GNAME51433(G51433,G55210,G51422);
  and GNAME51434(G51434,G55210,G51422);
  xor GNAME51439(G51439,G55236,G51428);
  and GNAME51440(G51440,G55236,G51428);
  xor GNAME51445(G51445,G55223,G51434);
  and GNAME51446(G51446,G55223,G51434);
  xor GNAME51451(G51451,G55249,G51440);
  and GNAME51452(G51452,G55249,G51440);
  xor GNAME51457(G51457,G55353,G51482);
  and GNAME51458(G51458,G55353,G51482);
  xor GNAME51463(G51463,G55379,G51488);
  and GNAME51464(G51464,G55379,G51488);
  xor GNAME51469(G51469,G55470,G51458);
  and GNAME51470(G51470,G55470,G51458);
  xor GNAME51475(G51475,G55496,G51464);
  and GNAME51476(G51476,G55496,G51464);
  xor GNAME51481(G51481,G55340,G51446);
  and GNAME51482(G51482,G55340,G51446);
  xor GNAME51487(G51487,G55366,G51452);
  and GNAME51488(G51488,G55366,G51452);
  xor GNAME51493(G51493,G55483,G51470);
  and GNAME51494(G51494,G55483,G51470);
  xor GNAME51499(G51499,G55509,G51476);
  and GNAME51500(G51500,G55509,G51476);
  xor GNAME51505(G51505,G55600,G51494);
  and GNAME51506(G51506,G55600,G51494);
  xor GNAME51511(G51511,G55626,G51500);
  and GNAME51512(G51512,G55626,G51500);
  xor GNAME51517(G51517,G55613,G51506);
  and GNAME51518(G51518,G55613,G51506);
  xor GNAME51523(G51523,G55639,G51512);
  and GNAME51524(G51524,G55639,G51512);
  xor GNAME51529(G51529,G55730,G51518);
  and GNAME51530(G51530,G55730,G51518);
  xor GNAME51535(G51535,G55756,G51524);
  and GNAME51536(G51536,G55756,G51524);
  xor GNAME51541(G51541,G55743,G51530);
  and GNAME51542(G51542,G55743,G51530);
  xor GNAME51547(G51547,G55769,G51536);
  and GNAME51548(G51548,G55769,G51536);
  xor GNAME51553(G51553,G55860,G51542);
  and GNAME51554(G51554,G55860,G51542);
  xor GNAME51559(G51559,G55886,G51548);
  and GNAME51560(G51560,G55886,G51548);
  xor GNAME51565(G51565,G55873,G51554);
  and GNAME51566(G51566,G55873,G51554);
  xor GNAME51571(G51571,G55899,G51560);
  and GNAME51572(G51572,G55899,G51560);
  xor GNAME51577(G51577,G56003,G51566);
  and GNAME51578(G51578,G56003,G51566);
  xor GNAME51583(G51583,G56081,G51572);
  and GNAME51584(G51584,G56081,G51572);
  xor GNAME51589(G51589,G56016,G51578);
  and GNAME51590(G51590,G56016,G51578);
  xor GNAME51595(G51595,G56094,G51584);
  and GNAME51596(G51596,G56094,G51584);
  xor GNAME51601(G51601,G56185,G51590);
  and GNAME51602(G51602,G56185,G51590);
  xor GNAME51607(G51607,G56263,G51596);
  and GNAME51608(G51608,G56263,G51596);
  xor GNAME51613(G51613,G56198,G51602);
  and GNAME51614(G51614,G56198,G51602);
  xor GNAME51619(G51619,G56276,G51608);
  and GNAME51620(G51620,G56276,G51608);
  xor GNAME51625(G51625,G56380,G51614);
  and GNAME51626(G51626,G56380,G51614);
  xor GNAME51631(G51631,G56471,G51620);
  and GNAME51632(G51632,G56471,G51620);
  xor GNAME51637(G51637,G56393,G51626);
  and GNAME51638(G51638,G56393,G51626);
  xor GNAME51643(G51643,G56484,G51632);
  and GNAME51644(G51644,G56484,G51632);
  xor GNAME51649(G51649,G56575,G51638);
  and GNAME51650(G51650,G56575,G51638);
  xor GNAME51655(G51655,G56653,G51644);
  and GNAME51656(G51656,G56653,G51644);
  xor GNAME51661(G51661,G56588,G51650);
  and GNAME51662(G51662,G56588,G51650);
  xor GNAME51667(G51667,G56666,G51656);
  and GNAME51668(G51668,G56666,G51656);
  xor GNAME51673(G51673,G56757,G51662);
  and GNAME51674(G51674,G56757,G51662);
  xor GNAME51679(G51679,G56848,G51668);
  and GNAME51680(G51680,G56848,G51668);
  xor GNAME51685(G51685,G56770,G51674);
  and GNAME51686(G51686,G56770,G51674);
  xor GNAME51691(G51691,G56861,G51680);
  and GNAME51692(G51692,G56861,G51680);
  xor GNAME51697(G51697,G56952,G51686);
  and GNAME51698(G51698,G56952,G51686);
  xor GNAME51703(G51703,G57030,G51692);
  and GNAME51704(G51704,G57030,G51692);
  xor GNAME51709(G51709,G56965,G51698);
  and GNAME51710(G51710,G56965,G51698);
  xor GNAME51715(G51715,G57043,G51704);
  and GNAME51716(G51716,G57043,G51704);
  xor GNAME51721(G51721,G56029,G55990);
  and GNAME51722(G51722,G56029,G55990);
  xor GNAME51727(G51727,G57641,G51896);
  and GNAME51728(G51728,G57641,G51896);
  xor GNAME51733(G51733,G56042,G51722);
  and GNAME51734(G51734,G56042,G51722);
  xor GNAME51739(G51739,G56055,G51734);
  and GNAME51740(G51740,G56055,G51734);
  xor GNAME51745(G51745,G56068,G51740);
  and GNAME51746(G51746,G56068,G51740);
  xor GNAME51751(G51751,G56211,G51746);
  and GNAME51752(G51752,G56211,G51746);
  xor GNAME51757(G51757,G56224,G51752);
  and GNAME51758(G51758,G56224,G51752);
  xor GNAME51763(G51763,G56237,G51758);
  and GNAME51764(G51764,G56237,G51758);
  xor GNAME51769(G51769,G56250,G51764);
  and GNAME51770(G51770,G56250,G51764);
  xor GNAME51775(G51775,G56406,G51770);
  and GNAME51776(G51776,G56406,G51770);
  xor GNAME51781(G51781,G56419,G51776);
  and GNAME51782(G51782,G56419,G51776);
  xor GNAME51787(G51787,G56432,G51782);
  and GNAME51788(G51788,G56432,G51782);
  xor GNAME51793(G51793,G56445,G51788);
  and GNAME51794(G51794,G56445,G51788);
  xor GNAME51799(G51799,G56458,G51794);
  and GNAME51800(G51800,G56458,G51794);
  xor GNAME51805(G51805,G56601,G51800);
  and GNAME51806(G51806,G56601,G51800);
  xor GNAME51811(G51811,G56614,G51806);
  and GNAME51812(G51812,G56614,G51806);
  xor GNAME51817(G51817,G56627,G51812);
  and GNAME51818(G51818,G56627,G51812);
  xor GNAME51823(G51823,G56640,G51818);
  and GNAME51824(G51824,G56640,G51818);
  xor GNAME51829(G51829,G56783,G51824);
  and GNAME51830(G51830,G56783,G51824);
  xor GNAME51835(G51835,G56796,G51830);
  and GNAME51836(G51836,G56796,G51830);
  xor GNAME51841(G51841,G56809,G51836);
  and GNAME51842(G51842,G56809,G51836);
  xor GNAME51847(G51847,G56822,G51842);
  and GNAME51848(G51848,G56822,G51842);
  xor GNAME51853(G51853,G56835,G51848);
  and GNAME51854(G51854,G56835,G51848);
  xor GNAME51859(G51859,G56978,G51854);
  and GNAME51860(G51860,G56978,G51854);
  xor GNAME51865(G51865,G56991,G51860);
  and GNAME51866(G51866,G56991,G51860);
  xor GNAME51871(G51871,G57004,G51866);
  and GNAME51872(G51872,G57004,G51866);
  xor GNAME51877(G51877,G57017,G51872);
  and GNAME51878(G51878,G57017,G51872);
  xor GNAME51883(G51883,G57602,G51878);
  and GNAME51884(G51884,G57602,G51878);
  xor GNAME51889(G51889,G57615,G51884);
  and GNAME51890(G51890,G57615,G51884);
  xor GNAME51895(G51895,G57628,G51890);
  and GNAME51896(G51896,G57628,G51890);
  and GNAME51903(G51903,G50697,G51221);
  and GNAME51904(G51904,G53062,G50697);
  and GNAME51905(G51905,G51221,G53062);
  or GNAME51906(G51906,G51905,G51904,G51903);
  and GNAME51913(G51913,G50698,G51224);
  and GNAME51914(G51914,G53065,G50698);
  and GNAME51915(G51915,G51224,G53065);
  or GNAME51916(G51916,G51915,G51914,G51913);
  and GNAME51923(G51923,G50699,G51227);
  and GNAME51924(G51924,G53068,G50699);
  and GNAME51925(G51925,G51227,G53068);
  or GNAME51926(G51926,G51925,G51924,G51923);
  and GNAME51933(G51933,G51906,G54529);
  and GNAME51934(G51934,G51325,G51906);
  and GNAME51935(G51935,G54529,G51325);
  or GNAME51936(G51936,G51935,G51934,G51933);
  and GNAME51943(G51943,G51936,G51326);
  and GNAME51944(G51944,G40983,G51936);
  and GNAME51945(G51945,G51326,G40983);
  or GNAME51946(G51946,G51945,G51944,G51943);
  and GNAME51953(G51953,G51916,G54532);
  and GNAME51954(G51954,G51331,G51916);
  and GNAME51955(G51955,G54532,G51331);
  or GNAME51956(G51956,G51955,G51954,G51953);
  and GNAME51963(G51963,G51956,G51332);
  and GNAME51964(G51964,G40998,G51956);
  and GNAME51965(G51965,G51332,G40998);
  or GNAME51966(G51966,G51965,G51964,G51963);
  and GNAME51973(G51973,G51926,G54535);
  and GNAME51974(G51974,G51337,G51926);
  and GNAME51975(G51975,G54535,G51337);
  or GNAME51976(G51976,G51975,G51974,G51973);
  and GNAME51983(G51983,G51976,G51338);
  and GNAME51984(G51984,G41013,G51976);
  and GNAME51985(G51985,G51338,G41013);
  or GNAME51986(G51986,G51985,G51984,G51983);
  and GNAME51993(G51993,G51946,G40988);
  and GNAME51994(G51994,G40938,G51946);
  and GNAME51995(G51995,G40988,G40938);
  or GNAME51996(G51996,G51995,G51994,G51993);
  and GNAME52003(G52003,G51996,G40943);
  and GNAME52004(G52004,G44898,G51996);
  and GNAME52005(G52005,G40943,G44898);
  or GNAME52006(G52006,G52005,G52004,G52003);
  and GNAME52013(G52013,G51966,G41003);
  and GNAME52014(G52014,G40953,G51966);
  and GNAME52015(G52015,G41003,G40953);
  or GNAME52016(G52016,G52015,G52014,G52013);
  and GNAME52023(G52023,G52016,G40958);
  and GNAME52024(G52024,G44928,G52016);
  and GNAME52025(G52025,G40958,G44928);
  or GNAME52026(G52026,G52025,G52024,G52023);
  and GNAME52033(G52033,G51986,G41018);
  and GNAME52034(G52034,G40968,G51986);
  and GNAME52035(G52035,G41018,G40968);
  or GNAME52036(G52036,G52035,G52034,G52033);
  and GNAME52043(G52043,G52036,G40973);
  and GNAME52044(G52044,G44958,G52036);
  and GNAME52045(G52045,G40973,G44958);
  or GNAME52046(G52046,G52045,G52044,G52043);
  nor GNAME52047(G52047,G52117,G57852);
  nor GNAME52048(G52048,G57909,G54573);
  nor GNAME52049(G52049,G57910,G54574);
  nor GNAME52050(G52050,G57911,G54575);
  nor GNAME52051(G52051,G57910,G54576);
  nor GNAME52052(G52052,G57909,G54577);
  nor GNAME52053(G52053,G57911,G54578);
  nor GNAME52054(G52054,G57910,G54579);
  nor GNAME52055(G52055,G57909,G54580);
  nor GNAME52056(G52056,G57911,G54581);
  nor GNAME52057(G52057,G57910,G54582);
  nor GNAME52058(G52058,G57909,G54583);
  nor GNAME52059(G52059,G57911,G54584);
  nor GNAME52060(G52060,G57910,G54585);
  nor GNAME52061(G52061,G57909,G54586);
  nor GNAME52062(G52062,G57911,G54587);
  nor GNAME52063(G52063,G57910,G54588);
  nor GNAME52064(G52064,G57909,G54589);
  nor GNAME52065(G52065,G57911,G54590);
  nor GNAME52066(G52066,G57910,G54591);
  nor GNAME52067(G52067,G57909,G54592);
  nor GNAME52068(G52068,G57911,G54593);
  nor GNAME52069(G52069,G57910,G54594);
  nor GNAME52070(G52070,G57909,G54595);
  nor GNAME52071(G52071,G57911,G54596);
  nor GNAME52072(G52072,G57910,G54597);
  nor GNAME52073(G52073,G57909,G54598);
  nor GNAME52074(G52074,G57911,G54599);
  nor GNAME52075(G52075,G57910,G54600);
  nor GNAME52076(G52076,G57909,G54601);
  nor GNAME52077(G52077,G57911,G54602);
  nor GNAME52078(G52078,G57910,G54603);
  nor GNAME52079(G52079,G57909,G54604);
  nor GNAME52080(G52080,G57911,G54605);
  nor GNAME52081(G52081,G57912,G54609);
  nor GNAME52082(G52082,G57913,G54610);
  nor GNAME52083(G52083,G57914,G54611);
  nor GNAME52084(G52084,G57912,G54612);
  nor GNAME52085(G52085,G57913,G54613);
  nor GNAME52086(G52086,G57914,G54614);
  nor GNAME52087(G52087,G57912,G54615);
  nor GNAME52088(G52088,G57913,G54616);
  nor GNAME52089(G52089,G57914,G54617);
  nor GNAME52090(G52090,G57912,G54606);
  nor GNAME52091(G52091,G57913,G54607);
  nor GNAME52092(G52092,G57914,G54608);
  nor GNAME52093(G52093,G57912,G54618);
  nor GNAME52094(G52094,G57912,G54619);
  nor GNAME52095(G52095,G57913,G54620);
  nor GNAME52096(G52096,G57914,G54621);
  nor GNAME52097(G52097,G57913,G54622);
  nor GNAME52098(G52098,G57914,G54623);
  nor GNAME52099(G52099,G57912,G54624);
  nor GNAME52100(G52100,G57912,G54625);
  nor GNAME52101(G52101,G57913,G54626);
  nor GNAME52102(G52102,G57914,G54627);
  nor GNAME52103(G52103,G57913,G54628);
  nor GNAME52104(G52104,G57914,G54629);
  nor GNAME52105(G52105,G57912,G54630);
  nor GNAME52106(G52106,G57912,G54631);
  nor GNAME52107(G52107,G57913,G54632);
  nor GNAME52108(G52108,G57914,G54633);
  nor GNAME52109(G52109,G57913,G54634);
  nor GNAME52110(G52110,G57914,G54635);
  nor GNAME52111(G52111,G57912,G54636);
  nor GNAME52112(G52112,G57913,G54637);
  nor GNAME52113(G52113,G57914,G54638);
  nor GNAME52114(G52114,G57909,G54570);
  nor GNAME52115(G52115,G57910,G54571);
  nor GNAME52116(G52116,G57911,G54572);
  xnor GNAME52117(G52117,G54820,G3613);
  xnor GNAME52118(G52118,G2678,G2657);
  xnor GNAME52119(G52119,G2262,G2241);
  xnor GNAME52120(G52120,G1846,G1825);
  xnor GNAME52121(G52121,G2636,G2615);
  xnor GNAME52122(G52122,G2220,G2199);
  xnor GNAME52123(G52123,G1804,G1783);
  xnor GNAME52124(G52124,G2552,G2491);
  xnor GNAME52125(G52125,G2136,G2075);
  xnor GNAME52126(G52126,G1720,G1659);
  xnor GNAME52127(G52127,G2594,G2573);
  xnor GNAME52128(G52128,G2178,G2157);
  xnor GNAME52129(G52129,G1762,G1741);
  xnor GNAME52130(G52130,G2470,G2449);
  xnor GNAME52131(G52131,G2054,G2033);
  xnor GNAME52132(G52132,G1638,G1617);
  xnor GNAME52133(G52133,G2428,G2407);
  xnor GNAME52134(G52134,G2012,G1991);
  xnor GNAME52135(G52135,G1596,G1575);
  xnor GNAME52136(G52136,G2386,G2365);
  xnor GNAME52137(G52137,G1970,G1949);
  xnor GNAME52138(G52138,G1554,G1533);
  xnor GNAME52139(G52139,G57725,G57728);
  xnor GNAME52140(G52140,G57725,G57737);
  xnor GNAME52141(G52141,G57726,G57729);
  xnor GNAME52142(G52142,G57726,G57738);
  xnor GNAME52143(G52143,G57727,G57730);
  xnor GNAME52144(G52144,G57727,G57739);
  xnor GNAME52145(G52145,G57725,G57734);
  xnor GNAME52146(G52146,G57731,G57728);
  xnor GNAME52147(G52147,G57731,G57737);
  xnor GNAME52148(G52148,G57725,G57746);
  xnor GNAME52149(G52149,G57726,G57735);
  xnor GNAME52150(G52150,G57732,G57729);
  xnor GNAME52151(G52151,G57732,G57738);
  xnor GNAME52152(G52152,G57726,G57747);
  xnor GNAME52153(G52153,G57727,G57736);
  xnor GNAME52154(G52154,G57733,G57730);
  xnor GNAME52155(G52155,G57733,G57739);
  xnor GNAME52156(G52156,G57727,G57748);
  xnor GNAME52157(G52157,G57725,G57755);
  xnor GNAME52158(G52158,G57731,G57746);
  xnor GNAME52159(G52159,G57726,G57756);
  xnor GNAME52160(G52160,G57732,G57747);
  xnor GNAME52161(G52161,G57727,G57757);
  xnor GNAME52162(G52162,G57733,G57748);
  xnor GNAME52163(G52163,G57731,G57734);
  xnor GNAME52164(G52164,G57740,G57728);
  xnor GNAME52165(G52165,G57725,G57743);
  xnor GNAME52166(G52166,G57732,G57735);
  xnor GNAME52167(G52167,G57741,G57729);
  xnor GNAME52168(G52168,G57733,G57736);
  xnor GNAME52169(G52169,G57742,G57730);
  xnor GNAME52170(G52170,G57726,G57744);
  xnor GNAME52171(G52171,G57727,G57745);
  xnor GNAME52172(G52172,G57740,G57737);
  xnor GNAME52173(G52173,G57740,G57734);
  xnor GNAME52174(G52174,G57749,G57728);
  xnor GNAME52175(G52175,G57725,G57752);
  xnor GNAME52176(G52176,G57731,G57743);
  xnor GNAME52177(G52177,G57741,G57738);
  xnor GNAME52178(G52178,G57741,G57735);
  xnor GNAME52179(G52179,G57750,G57729);
  xnor GNAME52180(G52180,G57742,G57739);
  xnor GNAME52181(G52181,G57742,G57736);
  xnor GNAME52182(G52182,G57751,G57730);
  xnor GNAME52183(G52183,G57726,G57753);
  xnor GNAME52184(G52184,G57732,G57744);
  xnor GNAME52185(G52185,G57727,G57754);
  xnor GNAME52186(G52186,G57733,G57745);
  xnor GNAME52187(G52187,G57740,G57746);
  xnor GNAME52188(G52188,G57725,G57764);
  xnor GNAME52189(G52189,G57731,G57755);
  xnor GNAME52190(G52190,G57731,G57752);
  xnor GNAME52191(G52191,G57758,G57728);
  xnor GNAME52192(G52192,G57741,G57747);
  xnor GNAME52193(G52193,G57726,G57765);
  xnor GNAME52194(G52194,G57732,G57756);
  xnor GNAME52195(G52195,G57742,G57748);
  xnor GNAME52196(G52196,G57727,G57766);
  xnor GNAME52197(G52197,G57733,G57757);
  xnor GNAME52198(G52198,G57732,G57753);
  xnor GNAME52199(G52199,G57759,G57729);
  xnor GNAME52200(G52200,G57733,G57754);
  xnor GNAME52201(G52201,G57760,G57730);
  xnor GNAME52202(G52202,G57740,G57743);
  xnor GNAME52203(G52203,G57725,G57761);
  xnor GNAME52204(G52204,G57749,G57737);
  xnor GNAME52205(G52205,G57749,G57734);
  xnor GNAME52206(G52206,G57741,G57744);
  xnor GNAME52207(G52207,G57726,G57762);
  xnor GNAME52208(G52208,G57750,G57738);
  xnor GNAME52209(G52209,G57750,G57735);
  xnor GNAME52210(G52210,G57742,G57745);
  xnor GNAME52211(G52211,G57727,G57763);
  xnor GNAME52212(G52212,G57751,G57739);
  xnor GNAME52213(G52213,G57751,G57736);
  xnor GNAME52214(G52214,G57731,G57764);
  xnor GNAME52215(G52215,G57732,G57765);
  xnor GNAME52216(G52216,G57733,G57766);
  xnor GNAME52217(G52217,G57749,G57746);
  xnor GNAME52218(G52218,G57725,G57771);
  xnor GNAME52219(G52219,G57740,G57755);
  xnor GNAME52220(G52220,G57758,G57737);
  xnor GNAME52221(G52221,G57758,G57734);
  xnor GNAME52222(G52222,G57767,G57728);
  xnor GNAME52223(G52223,G57740,G57752);
  xnor GNAME52224(G52224,G57725,G57770);
  xnor GNAME52225(G52225,G57749,G57743);
  xnor GNAME52226(G52226,G57731,G57761);
  xnor GNAME52227(G52227,G57750,G57747);
  xnor GNAME52228(G52228,G57726,G57773);
  xnor GNAME52229(G52229,G57741,G57756);
  xnor GNAME52230(G52230,G57751,G57748);
  xnor GNAME52231(G52231,G57727,G57775);
  xnor GNAME52232(G52232,G57742,G57757);
  xnor GNAME52233(G52233,G57759,G57738);
  xnor GNAME52234(G52234,G57759,G57735);
  xnor GNAME52235(G52235,G57768,G57729);
  xnor GNAME52236(G52236,G57741,G57753);
  xnor GNAME52237(G52237,G57726,G57772);
  xnor GNAME52238(G52238,G57750,G57744);
  xnor GNAME52239(G52239,G57732,G57762);
  xnor GNAME52240(G52240,G57760,G57739);
  xnor GNAME52241(G52241,G57760,G57736);
  xnor GNAME52242(G52242,G57769,G57730);
  xnor GNAME52243(G52243,G57742,G57754);
  xnor GNAME52244(G52244,G57727,G57774);
  xnor GNAME52245(G52245,G57751,G57745);
  xnor GNAME52246(G52246,G57733,G57763);
  xnor GNAME52247(G52247,G57758,G57746);
  xnor GNAME52248(G52248,G57725,G57789);
  xnor GNAME52249(G52249,G57767,G57737);
  xnor GNAME52250(G52250,G57749,G57755);
  xnor GNAME52251(G52251,G57731,G57771);
  xnor GNAME52252(G52252,G57740,G57764);
  xnor GNAME52253(G52253,G57749,G57752);
  xnor GNAME52254(G52254,G57740,G57761);
  xnor GNAME52255(G52255,G57758,G57743);
  xnor GNAME52256(G52256,G57731,G57770);
  xnor GNAME52257(G52257,G57725,G57790);
  xnor GNAME52258(G52258,G57767,G57734);
  xnor GNAME52259(G52259,G57776,G57728);
  xnor GNAME52260(G52260,G57759,G57747);
  xnor GNAME52261(G52261,G57726,G57792);
  xnor GNAME52262(G52262,G57768,G57738);
  xnor GNAME52263(G52263,G57750,G57756);
  xnor GNAME52264(G52264,G57732,G57773);
  xnor GNAME52265(G52265,G57741,G57765);
  xnor GNAME52266(G52266,G57760,G57748);
  xnor GNAME52267(G52267,G57727,G57794);
  xnor GNAME52268(G52268,G57769,G57739);
  xnor GNAME52269(G52269,G57751,G57757);
  xnor GNAME52270(G52270,G57733,G57775);
  xnor GNAME52271(G52271,G57742,G57766);
  xnor GNAME52272(G52272,G57750,G57753);
  xnor GNAME52273(G52273,G57741,G57762);
  xnor GNAME52274(G52274,G57759,G57744);
  xnor GNAME52275(G52275,G57732,G57772);
  xnor GNAME52276(G52276,G57726,G57793);
  xnor GNAME52277(G52277,G57768,G57735);
  xnor GNAME52278(G52278,G57777,G57729);
  xnor GNAME52279(G52279,G57751,G57754);
  xnor GNAME52280(G52280,G57742,G57763);
  xnor GNAME52281(G52281,G57760,G57745);
  xnor GNAME52282(G52282,G57733,G57774);
  xnor GNAME52283(G52283,G57727,G57795);
  xnor GNAME52284(G52284,G57769,G57736);
  xnor GNAME52285(G52285,G57778,G57730);
  xnor GNAME52286(G52286,G57781,G57791);
  xnor GNAME52287(G52287,G57749,G57764);
  xnor GNAME52288(G52288,G57767,G57746);
  xnor GNAME52289(G52289,G57740,G57771);
  xnor GNAME52290(G52290,G57776,G57737);
  xnor GNAME52291(G52291,G57758,G57755);
  xnor GNAME52292(G52292,G57731,G57789);
  xnor GNAME52293(G52293,G57749,G57761);
  xnor GNAME52294(G52294,G57740,G57770);
  xnor GNAME52295(G52295,G57758,G57752);
  xnor GNAME52296(G52296,G57731,G57790);
  xnor GNAME52297(G52297,G57781,G57813);
  xnor GNAME52298(G52298,G57767,G57743);
  xnor GNAME52299(G52299,G57776,G57734);
  xnor GNAME52300(G52300,G57782,G57796);
  xnor GNAME52301(G52301,G57750,G57765);
  xnor GNAME52302(G52302,G57768,G57747);
  xnor GNAME52303(G52303,G57741,G57773);
  xnor GNAME52304(G52304,G57777,G57738);
  xnor GNAME52305(G52305,G57759,G57756);
  xnor GNAME52306(G52306,G57732,G57792);
  xnor GNAME52307(G52307,G57783,G57797);
  xnor GNAME52308(G52308,G57751,G57766);
  xnor GNAME52309(G52309,G57769,G57748);
  xnor GNAME52310(G52310,G57742,G57775);
  xnor GNAME52311(G52311,G57778,G57739);
  xnor GNAME52312(G52312,G57760,G57757);
  xnor GNAME52313(G52313,G57733,G57794);
  xnor GNAME52314(G52314,G57750,G57762);
  xnor GNAME52315(G52315,G57741,G57772);
  xnor GNAME52316(G52316,G57759,G57753);
  xnor GNAME52317(G52317,G57732,G57793);
  xnor GNAME52318(G52318,G57782,G57814);
  xnor GNAME52319(G52319,G57768,G57744);
  xnor GNAME52320(G52320,G57777,G57735);
  xnor GNAME52321(G52321,G57751,G57763);
  xnor GNAME52322(G52322,G57742,G57774);
  xnor GNAME52323(G52323,G57760,G57754);
  xnor GNAME52324(G52324,G57733,G57795);
  xnor GNAME52325(G52325,G57783,G57815);
  xnor GNAME52326(G52326,G57769,G57745);
  xnor GNAME52327(G52327,G57778,G57736);
  xnor GNAME52328(G52328,G57798,G57728);
  xnor GNAME52329(G52329,G57799,G57729);
  xnor GNAME52330(G52330,G57800,G57730);
  xnor GNAME52331(G52331,G57749,G57771);
  xnor GNAME52332(G52332,G57740,G57789);
  xnor GNAME52333(G52333,G57758,G57764);
  xnor GNAME52334(G52334,G57784,G57791);
  xnor GNAME52335(G52335,G57781,G57808);
  xnor GNAME52336(G52336,G57767,G57755);
  xnor GNAME52337(G52337,G57776,G57746);
  xnor GNAME52338(G52338,G57749,G57770);
  xnor GNAME52339(G52339,G57740,G57790);
  xnor GNAME52340(G52340,G57758,G57761);
  xnor GNAME52341(G52341,G57784,G57813);
  xnor GNAME52342(G52342,G57781,G57807);
  xnor GNAME52343(G52343,G57767,G57752);
  xnor GNAME52344(G52344,G57776,G57743);
  xnor GNAME52345(G52345,G57750,G57773);
  xnor GNAME52346(G52346,G57741,G57792);
  xnor GNAME52347(G52347,G57759,G57765);
  xnor GNAME52348(G52348,G57785,G57796);
  xnor GNAME52349(G52349,G57782,G57810);
  xnor GNAME52350(G52350,G57768,G57756);
  xnor GNAME52351(G52351,G57777,G57747);
  xnor GNAME52352(G52352,G57751,G57775);
  xnor GNAME52353(G52353,G57742,G57794);
  xnor GNAME52354(G52354,G57760,G57766);
  xnor GNAME52355(G52355,G57786,G57797);
  xnor GNAME52356(G52356,G57783,G57812);
  xnor GNAME52357(G52357,G57769,G57757);
  xnor GNAME52358(G52358,G57778,G57748);
  xnor GNAME52359(G52359,G57750,G57772);
  xnor GNAME52360(G52360,G57741,G57793);
  xnor GNAME52361(G52361,G57759,G57762);
  xnor GNAME52362(G52362,G57785,G57814);
  xnor GNAME52363(G52363,G57782,G57809);
  xnor GNAME52364(G52364,G57768,G57753);
  xnor GNAME52365(G52365,G57777,G57744);
  xnor GNAME52366(G52366,G57751,G57774);
  xnor GNAME52367(G52367,G57742,G57795);
  xnor GNAME52368(G52368,G57760,G57763);
  xnor GNAME52369(G52369,G57786,G57815);
  xnor GNAME52370(G52370,G57783,G57811);
  xnor GNAME52371(G52371,G57769,G57754);
  xnor GNAME52372(G52372,G57778,G57745);
  xnor GNAME52373(G52373,G57798,G57737);
  xnor GNAME52374(G52374,G57798,G57734);
  xnor GNAME52375(G52375,G57799,G57738);
  xnor GNAME52376(G52376,G57800,G57739);
  xnor GNAME52377(G52377,G57799,G57735);
  xnor GNAME52378(G52378,G57800,G57736);
  xnor GNAME52379(G52379,G57749,G57789);
  xnor GNAME52380(G52380,G57801,G57791);
  xnor GNAME52381(G52381,G57758,G57771);
  xnor GNAME52382(G52382,G57784,G57808);
  xnor GNAME52383(G52383,G57781,G57822);
  xnor GNAME52384(G52384,G57767,G57764);
  xnor GNAME52385(G52385,G57776,G57755);
  xnor GNAME52386(G52386,G57749,G57790);
  xnor GNAME52387(G52387,G57801,G57813);
  xnor GNAME52388(G52388,G57758,G57770);
  xnor GNAME52389(G52389,G57784,G57807);
  xnor GNAME52390(G52390,G57781,G57819);
  xnor GNAME52391(G52391,G57767,G57761);
  xnor GNAME52392(G52392,G57776,G57752);
  xnor GNAME52393(G52393,G57750,G57792);
  xnor GNAME52394(G52394,G57802,G57796);
  xnor GNAME52395(G52395,G57759,G57773);
  xnor GNAME52396(G52396,G57785,G57810);
  xnor GNAME52397(G52397,G57782,G57823);
  xnor GNAME52398(G52398,G57768,G57765);
  xnor GNAME52399(G52399,G57777,G57756);
  xnor GNAME52400(G52400,G57751,G57794);
  xnor GNAME52401(G52401,G57803,G57797);
  xnor GNAME52402(G52402,G57760,G57775);
  xnor GNAME52403(G52403,G57786,G57812);
  xnor GNAME52404(G52404,G57783,G57824);
  xnor GNAME52405(G52405,G57769,G57766);
  xnor GNAME52406(G52406,G57778,G57757);
  xnor GNAME52407(G52407,G57750,G57793);
  xnor GNAME52408(G52408,G57802,G57814);
  xnor GNAME52409(G52409,G57759,G57772);
  xnor GNAME52410(G52410,G57785,G57809);
  xnor GNAME52411(G52411,G57782,G57827);
  xnor GNAME52412(G52412,G57768,G57762);
  xnor GNAME52413(G52413,G57777,G57753);
  xnor GNAME52414(G52414,G57751,G57795);
  xnor GNAME52415(G52415,G57803,G57815);
  xnor GNAME52416(G52416,G57760,G57774);
  xnor GNAME52417(G52417,G57786,G57811);
  xnor GNAME52418(G52418,G57783,G57830);
  xnor GNAME52419(G52419,G57769,G57763);
  xnor GNAME52420(G52420,G57778,G57754);
  xnor GNAME52421(G52421,G57798,G57746);
  xnor GNAME52422(G52422,G57798,G57743);
  xnor GNAME52423(G52423,G57799,G57747);
  xnor GNAME52424(G52424,G57800,G57748);
  xnor GNAME52425(G52425,G57799,G57744);
  xnor GNAME52426(G52426,G57800,G57745);
  xnor GNAME52427(G52427,G57816,G57791);
  xnor GNAME52428(G52428,G57801,G57808);
  xnor GNAME52429(G52429,G57758,G57789);
  xnor GNAME52430(G52430,G57784,G57822);
  xnor GNAME52431(G52431,G57781,G57820);
  xnor GNAME52432(G52432,G57767,G57771);
  xnor GNAME52433(G52433,G57776,G57764);
  xnor GNAME52434(G52434,G57816,G57813);
  xnor GNAME52435(G52435,G57801,G57807);
  xnor GNAME52436(G52436,G57758,G57790);
  xnor GNAME52437(G52437,G57784,G57819);
  xnor GNAME52438(G52438,G57781,G57821);
  xnor GNAME52439(G52439,G57767,G57770);
  xnor GNAME52440(G52440,G57776,G57761);
  xnor GNAME52441(G52441,G57817,G57796);
  xnor GNAME52442(G52442,G57802,G57810);
  xnor GNAME52443(G52443,G57759,G57792);
  xnor GNAME52444(G52444,G57785,G57823);
  xnor GNAME52445(G52445,G57782,G57826);
  xnor GNAME52446(G52446,G57768,G57773);
  xnor GNAME52447(G52447,G57777,G57765);
  xnor GNAME52448(G52448,G57818,G57797);
  xnor GNAME52449(G52449,G57803,G57812);
  xnor GNAME52450(G52450,G57760,G57794);
  xnor GNAME52451(G52451,G57786,G57824);
  xnor GNAME52452(G52452,G57783,G57829);
  xnor GNAME52453(G52453,G57769,G57775);
  xnor GNAME52454(G52454,G57778,G57766);
  xnor GNAME52455(G52455,G57817,G57814);
  xnor GNAME52456(G52456,G57802,G57809);
  xnor GNAME52457(G52457,G57759,G57793);
  xnor GNAME52458(G52458,G57785,G57827);
  xnor GNAME52459(G52459,G57782,G57825);
  xnor GNAME52460(G52460,G57768,G57772);
  xnor GNAME52461(G52461,G57777,G57762);
  xnor GNAME52462(G52462,G57818,G57815);
  xnor GNAME52463(G52463,G57803,G57811);
  xnor GNAME52464(G52464,G57760,G57795);
  xnor GNAME52465(G52465,G57786,G57830);
  xnor GNAME52466(G52466,G57783,G57828);
  xnor GNAME52467(G52467,G57769,G57774);
  xnor GNAME52468(G52468,G57778,G57763);
  xnor GNAME52469(G52469,G57798,G57755);
  xnor GNAME52470(G52470,G57798,G57752);
  xnor GNAME52471(G52471,G57799,G57756);
  xnor GNAME52472(G52472,G57800,G57757);
  xnor GNAME52473(G52473,G57799,G57753);
  xnor GNAME52474(G52474,G57800,G57754);
  xnor GNAME52475(G52475,G57767,G57790);
  xnor GNAME52476(G52476,G57768,G57793);
  xnor GNAME52477(G52477,G57769,G57795);
  xnor GNAME52478(G52478,G57816,G57808);
  xnor GNAME52479(G52479,G57801,G57822);
  xnor GNAME52480(G52480,G57831,G57791);
  xnor GNAME52481(G52481,G57784,G57820);
  xnor GNAME52482(G52482,G57781,G57840);
  xnor GNAME52483(G52483,G57767,G57789);
  xnor GNAME52484(G52484,G57776,G57771);
  xnor GNAME52485(G52485,G57816,G57807);
  xnor GNAME52486(G52486,G57801,G57819);
  xnor GNAME52487(G52487,G57831,G57813);
  xnor GNAME52488(G52488,G57784,G57821);
  xnor GNAME52489(G52489,G57776,G57770);
  xnor GNAME52490(G52490,G57817,G57810);
  xnor GNAME52491(G52491,G57802,G57823);
  xnor GNAME52492(G52492,G57832,G57796);
  xnor GNAME52493(G52493,G57785,G57826);
  xnor GNAME52494(G52494,G57782,G57842);
  xnor GNAME52495(G52495,G57768,G57792);
  xnor GNAME52496(G52496,G57777,G57773);
  xnor GNAME52497(G52497,G57818,G57812);
  xnor GNAME52498(G52498,G57803,G57824);
  xnor GNAME52499(G52499,G57833,G57797);
  xnor GNAME52500(G52500,G57786,G57829);
  xnor GNAME52501(G52501,G57783,G57844);
  xnor GNAME52502(G52502,G57769,G57794);
  xnor GNAME52503(G52503,G57778,G57775);
  xnor GNAME52504(G52504,G57817,G57809);
  xnor GNAME52505(G52505,G57802,G57827);
  xnor GNAME52506(G52506,G57832,G57814);
  xnor GNAME52507(G52507,G57785,G57825);
  xnor GNAME52508(G52508,G57777,G57772);
  xnor GNAME52509(G52509,G57818,G57811);
  xnor GNAME52510(G52510,G57803,G57830);
  xnor GNAME52511(G52511,G57833,G57815);
  xnor GNAME52512(G52512,G57786,G57828);
  xnor GNAME52513(G52513,G57778,G57774);
  xnor GNAME52514(G52514,G57798,G57764);
  xnor GNAME52515(G52515,G57799,G57765);
  xnor GNAME52516(G52516,G57800,G57766);
  xnor GNAME52517(G52517,G57784,G57804);
  xnor GNAME52518(G52518,G57785,G57805);
  xnor GNAME52519(G52519,G57786,G57806);
  xnor GNAME52520(G52520,G57781,G57804);
  xnor GNAME52521(G52521,G57782,G57805);
  xnor GNAME52522(G52522,G57783,G57806);
  xnor GNAME52523(G52523,G57831,G57822);
  xnor GNAME52524(G52524,G57832,G57823);
  xnor GNAME52525(G52525,G57833,G57824);
  xnor GNAME52526(G52526,G57781,G57841);
  xnor GNAME52527(G52527,G57831,G57808);
  xnor GNAME52528(G52528,G57776,G57789);
  xnor GNAME52529(G52529,G57801,G57820);
  xnor GNAME52530(G52530,G57784,G57840);
  xnor GNAME52531(G52531,G57816,G57822);
  xnor GNAME52532(G52532,G57776,G57790);
  xnor GNAME52533(G52533,G57801,G57821);
  xnor GNAME52534(G52534,G57784,G57841);
  xnor GNAME52535(G52535,G57834,G57791);
  xnor GNAME52536(G52536,G57834,G57813);
  xnor GNAME52537(G52537,G57816,G57819);
  xnor GNAME52538(G52538,G57831,G57807);
  xnor GNAME52539(G52539,G57782,G57843);
  xnor GNAME52540(G52540,G57832,G57810);
  xnor GNAME52541(G52541,G57777,G57792);
  xnor GNAME52542(G52542,G57802,G57826);
  xnor GNAME52543(G52543,G57785,G57842);
  xnor GNAME52544(G52544,G57817,G57823);
  xnor GNAME52545(G52545,G57783,G57845);
  xnor GNAME52546(G52546,G57833,G57812);
  xnor GNAME52547(G52547,G57778,G57794);
  xnor GNAME52548(G52548,G57803,G57829);
  xnor GNAME52549(G52549,G57786,G57844);
  xnor GNAME52550(G52550,G57818,G57824);
  xnor GNAME52551(G52551,G57777,G57793);
  xnor GNAME52552(G52552,G57802,G57825);
  xnor GNAME52553(G52553,G57785,G57843);
  xnor GNAME52554(G52554,G57835,G57796);
  xnor GNAME52555(G52555,G57835,G57814);
  xnor GNAME52556(G52556,G57817,G57827);
  xnor GNAME52557(G52557,G57832,G57809);
  xnor GNAME52558(G52558,G57778,G57795);
  xnor GNAME52559(G52559,G57803,G57828);
  xnor GNAME52560(G52560,G57786,G57845);
  xnor GNAME52561(G52561,G57836,G57797);
  xnor GNAME52562(G52562,G57836,G57815);
  xnor GNAME52563(G52563,G57818,G57830);
  xnor GNAME52564(G52564,G57833,G57811);
  xnor GNAME52565(G52565,G57798,G57761);
  xnor GNAME52566(G52566,G57798,G57771);
  xnor GNAME52567(G52567,G57798,G57770);
  xnor GNAME52568(G52568,G57799,G57762);
  xnor GNAME52569(G52569,G57799,G57773);
  xnor GNAME52570(G52570,G57800,G57763);
  xnor GNAME52571(G52571,G57800,G57775);
  xnor GNAME52572(G52572,G57799,G57772);
  xnor GNAME52573(G52573,G57800,G57774);
  xnor GNAME52574(G52574,G57816,G57821);
  xnor GNAME52575(G52575,G57816,G57840);
  xnor GNAME52576(G52576,G57834,G57807);
  xnor GNAME52577(G52577,G57834,G57822);
  xnor GNAME52578(G52578,G57831,G57820);
  xnor GNAME52579(G52579,G57817,G57825);
  xnor GNAME52580(G52580,G57817,G57842);
  xnor GNAME52581(G52581,G57835,G57809);
  xnor GNAME52582(G52582,G57835,G57823);
  xnor GNAME52583(G52583,G57832,G57826);
  xnor GNAME52584(G52584,G57818,G57828);
  xnor GNAME52585(G52585,G57818,G57844);
  xnor GNAME52586(G52586,G57836,G57811);
  xnor GNAME52587(G52587,G57836,G57824);
  xnor GNAME52588(G52588,G57833,G57829);
  xnor GNAME52589(G52589,G57801,G57840);
  xnor GNAME52590(G52590,G57834,G57808);
  xnor GNAME52591(G52591,G57846,G57791);
  xnor GNAME52592(G52592,G57816,G57820);
  xnor GNAME52593(G52593,G57801,G57841);
  xnor GNAME52594(G52594,G57846,G57813);
  xnor GNAME52595(G52595,G57831,G57819);
  xnor GNAME52596(G52596,G57802,G57842);
  xnor GNAME52597(G52597,G57835,G57810);
  xnor GNAME52598(G52598,G57847,G57796);
  xnor GNAME52599(G52599,G57817,G57826);
  xnor GNAME52600(G52600,G57803,G57844);
  xnor GNAME52601(G52601,G57836,G57812);
  xnor GNAME52602(G52602,G57848,G57797);
  xnor GNAME52603(G52603,G57818,G57829);
  xnor GNAME52604(G52604,G57802,G57843);
  xnor GNAME52605(G52605,G57847,G57814);
  xnor GNAME52606(G52606,G57832,G57827);
  xnor GNAME52607(G52607,G57803,G57845);
  xnor GNAME52608(G52608,G57848,G57815);
  xnor GNAME52609(G52609,G57833,G57830);
  xnor GNAME52610(G52610,G57798,G57789);
  xnor GNAME52611(G52611,G57798,G57790);
  xnor GNAME52612(G52612,G57799,G57792);
  xnor GNAME52613(G52613,G57799,G57793);
  xnor GNAME52614(G52614,G57800,G57794);
  xnor GNAME52615(G52615,G57800,G57795);
  xnor GNAME52616(G52616,G57801,G57804);
  xnor GNAME52617(G52617,G57802,G57805);
  xnor GNAME52618(G52618,G57803,G57806);
  xnor GNAME52619(G52619,G57816,G57804);
  xnor GNAME52620(G52620,G57817,G57805);
  xnor GNAME52621(G52621,G57818,G57806);
  xnor GNAME52622(G52622,G57846,G57807);
  xnor GNAME52623(G52623,G57831,G57840);
  xnor GNAME52624(G52624,G57834,G57820);
  xnor GNAME52625(G52625,G57847,G57809);
  xnor GNAME52626(G52626,G57848,G57811);
  xnor GNAME52627(G52627,G57832,G57842);
  xnor GNAME52628(G52628,G57835,G57826);
  xnor GNAME52629(G52629,G57833,G57844);
  xnor GNAME52630(G52630,G57836,G57829);
  xnor GNAME52631(G52631,G57831,G57821);
  xnor GNAME52632(G52632,G57816,G57841);
  xnor GNAME52633(G52633,G57834,G57819);
  xnor GNAME52634(G52634,G57846,G57808);
  xnor GNAME52635(G52635,G57846,G57822);
  xnor GNAME52636(G52636,G57831,G57841);
  xnor GNAME52637(G52637,G57832,G57825);
  xnor GNAME52638(G52638,G57817,G57843);
  xnor GNAME52639(G52639,G57835,G57827);
  xnor GNAME52640(G52640,G57847,G57810);
  xnor GNAME52641(G52641,G57833,G57828);
  xnor GNAME52642(G52642,G57818,G57845);
  xnor GNAME52643(G52643,G57836,G57830);
  xnor GNAME52644(G52644,G57848,G57812);
  xnor GNAME52645(G52645,G57847,G57823);
  xnor GNAME52646(G52646,G57848,G57824);
  xnor GNAME52647(G52647,G57832,G57843);
  xnor GNAME52648(G52648,G57833,G57845);
  xnor GNAME52649(G52649,G57849,G57791);
  xnor GNAME52650(G52650,G57849,G57813);
  xnor GNAME52651(G52651,G57849,G57808);
  xnor GNAME52652(G52652,G57849,G57807);
  xnor GNAME52653(G52653,G57850,G57796);
  xnor GNAME52654(G52654,G57850,G57814);
  xnor GNAME52655(G52655,G57851,G57797);
  xnor GNAME52656(G52656,G57851,G57815);
  xnor GNAME52657(G52657,G57850,G57810);
  xnor GNAME52658(G52658,G57850,G57809);
  xnor GNAME52659(G52659,G57851,G57812);
  xnor GNAME52660(G52660,G57851,G57811);
  xnor GNAME52661(G52661,G57831,G57837);
  xnor GNAME52662(G52662,G57832,G57838);
  xnor GNAME52663(G52663,G57833,G57839);
  xnor GNAME52664(G52664,G57834,G57837);
  xnor GNAME52665(G52665,G57835,G57838);
  xnor GNAME52666(G52666,G57836,G57839);
  xnor GNAME52667(G52667,G57834,G57840);
  xnor GNAME52668(G52668,G57834,G57821);
  xnor GNAME52669(G52669,G57846,G57819);
  xnor GNAME52670(G52670,G57846,G57820);
  xnor GNAME52671(G52671,G57835,G57825);
  xnor GNAME52672(G52672,G57835,G57842);
  xnor GNAME52673(G52673,G57847,G57827);
  xnor GNAME52674(G52674,G57847,G57826);
  xnor GNAME52675(G52675,G57836,G57828);
  xnor GNAME52676(G52676,G57836,G57844);
  xnor GNAME52677(G52677,G57848,G57830);
  xnor GNAME52678(G52678,G57848,G57829);
  xnor GNAME52679(G52679,G57846,G57821);
  xnor GNAME52680(G52680,G57834,G57841);
  xnor GNAME52681(G52681,G57847,G57825);
  xnor GNAME52682(G52682,G57835,G57843);
  xnor GNAME52683(G52683,G57848,G57828);
  xnor GNAME52684(G52684,G57836,G57845);
  xnor GNAME52685(G52685,G57849,G57819);
  xnor GNAME52686(G52686,G57849,G57822);
  xnor GNAME52687(G52687,G57850,G57823);
  xnor GNAME52688(G52688,G57851,G57824);
  xnor GNAME52689(G52689,G57850,G57827);
  xnor GNAME52690(G52690,G57851,G57830);
  xnor GNAME52691(G52691,G57846,G57840);
  xnor GNAME52692(G52692,G57846,G57841);
  xnor GNAME52693(G52693,G57847,G57842);
  xnor GNAME52694(G52694,G57847,G57843);
  xnor GNAME52695(G52695,G57848,G57844);
  xnor GNAME52696(G52696,G57848,G57845);
  xnor GNAME52697(G52697,G57849,G57820);
  xnor GNAME52698(G52698,G57849,G57821);
  xnor GNAME52699(G52699,G57850,G57826);
  xnor GNAME52700(G52700,G57850,G57825);
  xnor GNAME52701(G52701,G57851,G57829);
  xnor GNAME52702(G52702,G57851,G57828);
  xnor GNAME52703(G52703,G57849,G57840);
  xnor GNAME52704(G52704,G57849,G57841);
  xnor GNAME52705(G52705,G57850,G57842);
  xnor GNAME52706(G52706,G57850,G57843);
  xnor GNAME52707(G52707,G57851,G57844);
  xnor GNAME52708(G52708,G57851,G57845);
  xnor GNAME52709(G52709,G57849,G57837);
  xnor GNAME52710(G52710,G57850,G57838);
  xnor GNAME52711(G52711,G57851,G57839);
  xnor GNAME52712(G52712,G57846,G57837);
  xnor GNAME52713(G52713,G57847,G57838);
  xnor GNAME52714(G52714,G57848,G57839);
  and GNAME52715(G52715,G57922,G57854);
  or GNAME52716(G52716,G54639,G52715);
  and GNAME52717(G52717,G57921,G57853);
  or GNAME52718(G52718,G54640,G52717);
  and GNAME52719(G52719,G57923,G57855);
  or GNAME52720(G52720,G54641,G52719);
  and GNAME52721(G52721,G57927,G57861);
  or GNAME52722(G52722,G54642,G52721);
  and GNAME52723(G52723,G57928,G57862);
  or GNAME52724(G52724,G54643,G52723);
  and GNAME52725(G52725,G57929,G57863);
  or GNAME52726(G52726,G54644,G52725);
  and GNAME52727(G52727,G57876,G57867);
  or GNAME52728(G52728,G54647,G52727);
  and GNAME52729(G52729,G57878,G57869);
  or GNAME52730(G52730,G54649,G52729);
  and GNAME52731(G52731,G57879,G57870);
  or GNAME52732(G52732,G54650,G52731);
  and GNAME52733(G52733,G57877,G57868);
  or GNAME52734(G52734,G54648,G52733);
  and GNAME52735(G52735,G57880,G57871);
  or GNAME52736(G52736,G54651,G52735);
  and GNAME52737(G52737,G57881,G57872);
  or GNAME52738(G52738,G54652,G52737);
  and GNAME52739(G52739,G57954,G57930);
  or GNAME52740(G52740,G54653,G52739);
  and GNAME52741(G52741,G57955,G57931);
  or GNAME52742(G52742,G54654,G52741);
  and GNAME52743(G52743,G57956,G57932);
  or GNAME52744(G52744,G54655,G52743);
  and GNAME52745(G52745,G57951,G57933);
  or GNAME52746(G52746,G54659,G52745);
  and GNAME52747(G52747,G57952,G57934);
  or GNAME52748(G52748,G54656,G52747);
  and GNAME52749(G52749,G57953,G57935);
  or GNAME52750(G52750,G54657,G52749);
  and GNAME52751(G52751,G57906,G57888);
  or GNAME52752(G52752,G54658,G52751);
  and GNAME52753(G52753,G57907,G57889);
  or GNAME52754(G52754,G54660,G52753);
  and GNAME52755(G52755,G57908,G57890);
  or GNAME52756(G52756,G54661,G52755);
  and GNAME52757(G52757,G57891,G57885);
  or GNAME52758(G52758,G54662,G52757);
  and GNAME52759(G52759,G57892,G57886);
  or GNAME52760(G52760,G54663,G52759);
  and GNAME52761(G52761,G57893,G57887);
  or GNAME52762(G52762,G54664,G52761);
  or GNAME52763(G52763,G57921,G52139);
  or GNAME52764(G52764,G57853,G52140);
  nand GNAME52765(G52765,G52764,G52763);
  or GNAME52766(G52766,G57922,G52141);
  or GNAME52767(G52767,G57854,G52142);
  nand GNAME52768(G52768,G52767,G52766);
  or GNAME52769(G52769,G57923,G52143);
  or GNAME52770(G52770,G57855,G52144);
  nand GNAME52771(G52771,G52770,G52769);
  or GNAME52772(G52772,G57927,G52146);
  or GNAME52773(G52773,G57861,G52147);
  nand GNAME52774(G52774,G52773,G52772);
  or GNAME52775(G52775,G57928,G52150);
  or GNAME52776(G52776,G57862,G52151);
  nand GNAME52777(G52777,G52776,G52775);
  or GNAME52778(G52778,G57929,G52154);
  or GNAME52779(G52779,G57863,G52155);
  nand GNAME52780(G52780,G52779,G52778);
  or GNAME52781(G52781,G57876,G52164);
  or GNAME52782(G52782,G57867,G52172);
  nand GNAME52783(G52783,G52782,G52781);
  or GNAME52784(G52784,G57878,G52167);
  or GNAME52785(G52785,G57869,G52177);
  nand GNAME52786(G52786,G52785,G52784);
  or GNAME52787(G52787,G57879,G52169);
  or GNAME52788(G52788,G57870,G52180);
  nand GNAME52789(G52789,G52788,G52787);
  or GNAME52790(G52790,G57876,G52173);
  or GNAME52791(G52791,G57867,G52187);
  nand GNAME52792(G52792,G52791,G52790);
  or GNAME52793(G52793,G57878,G52178);
  or GNAME52794(G52794,G57869,G52192);
  nand GNAME52795(G52795,G52794,G52793);
  or GNAME52796(G52796,G57879,G52181);
  or GNAME52797(G52797,G57870,G52195);
  nand GNAME52798(G52798,G52797,G52796);
  or GNAME52799(G52799,G57877,G52205);
  or GNAME52800(G52800,G57868,G52217);
  nand GNAME52801(G52801,G52800,G52799);
  or GNAME52802(G52802,G57880,G52209);
  or GNAME52803(G52803,G57871,G52227);
  nand GNAME52804(G52804,G52803,G52802);
  or GNAME52805(G52805,G57881,G52213);
  or GNAME52806(G52806,G57872,G52230);
  nand GNAME52807(G52807,G52806,G52805);
  or GNAME52808(G52808,G57877,G52225);
  or GNAME52809(G52809,G57868,G52250);
  nand GNAME52810(G52810,G52809,G52808);
  or GNAME52811(G52811,G57880,G52238);
  or GNAME52812(G52812,G57871,G52263);
  nand GNAME52813(G52813,G52812,G52811);
  or GNAME52814(G52814,G57881,G52245);
  or GNAME52815(G52815,G57872,G52269);
  nand GNAME52816(G52816,G52815,G52814);
  or GNAME52817(G52817,G57906,G54658);
  or GNAME52818(G52818,G57888,G52259);
  nand GNAME52819(G52819,G52818,G52817);
  or GNAME52820(G52820,G57907,G54660);
  or GNAME52821(G52821,G57889,G52278);
  nand GNAME52822(G52822,G52821,G52820);
  or GNAME52823(G52823,G57908,G54661);
  or GNAME52824(G52824,G57890,G52285);
  nand GNAME52825(G52825,G52824,G52823);
  or GNAME52826(G52826,G57906,G52484);
  or GNAME52827(G52827,G57888,G52489);
  nand GNAME52828(G52828,G52827,G52826);
  or GNAME52829(G52829,G52514,G57891);
  or GNAME52830(G52830,G57885,G52565);
  nand GNAME52831(G52831,G52830,G52829);
  or GNAME52832(G52832,G57907,G52496);
  or GNAME52833(G52833,G57889,G52508);
  nand GNAME52834(G52834,G52833,G52832);
  or GNAME52835(G52835,G52515,G57892);
  or GNAME52836(G52836,G57886,G52568);
  nand GNAME52837(G52837,G52836,G52835);
  or GNAME52838(G52838,G57908,G52503);
  or GNAME52839(G52839,G57890,G52513);
  nand GNAME52840(G52840,G52839,G52838);
  or GNAME52841(G52841,G52516,G57893);
  or GNAME52842(G52842,G57887,G52570);
  nand GNAME52843(G52843,G52842,G52841);
  or GNAME52844(G52844,G57901,G52528);
  or GNAME52845(G52845,G57897,G52532);
  nand GNAME52846(G52846,G52845,G52844);
  or GNAME52847(G52847,G52566,G57891);
  or GNAME52848(G52848,G57885,G52567);
  nand GNAME52849(G52849,G52848,G52847);
  or GNAME52850(G52850,G57903,G52541);
  or GNAME52851(G52851,G57898,G52551);
  nand GNAME52852(G52852,G52851,G52850);
  or GNAME52853(G52853,G52569,G57892);
  or GNAME52854(G52854,G57886,G52572);
  nand GNAME52855(G52855,G52854,G52853);
  or GNAME52856(G52856,G57905,G52547);
  or GNAME52857(G52857,G57899,G52558);
  nand GNAME52858(G52858,G52857,G52856);
  or GNAME52859(G52859,G52571,G57893);
  or GNAME52860(G52860,G57887,G52573);
  nand GNAME52861(G52861,G52860,G52859);
  or GNAME52862(G52862,G57864,G52534);
  or GNAME52863(G52863,G57916,G52517);
  nand GNAME52864(G52864,G52863,G52862);
  or GNAME52865(G52865,G52567,G57891);
  or GNAME52866(G52866,G57894,G52610);
  nand GNAME52867(G52867,G52866,G52865);
  or GNAME52868(G52868,G57865,G52553);
  or GNAME52869(G52869,G57919,G52518);
  nand GNAME52870(G52870,G52869,G52868);
  or GNAME52871(G52871,G52572,G57892);
  or GNAME52872(G52872,G57895,G52612);
  nand GNAME52873(G52873,G52872,G52871);
  or GNAME52874(G52874,G57866,G52560);
  or GNAME52875(G52875,G57920,G52519);
  nand GNAME52876(G52876,G52875,G52874);
  or GNAME52877(G52877,G52573,G57893);
  or GNAME52878(G52878,G57896,G52614);
  nand GNAME52879(G52879,G52878,G52877);
  or GNAME52880(G52880,G57858,G52526);
  or GNAME52881(G52881,G57915,G52520);
  nand GNAME52882(G52882,G52881,G52880);
  or GNAME52883(G52883,G52565,G57891);
  or GNAME52884(G52884,G57885,G52566);
  nand GNAME52885(G52885,G52884,G52883);
  or GNAME52886(G52886,G57859,G52539);
  or GNAME52887(G52887,G57917,G52521);
  nand GNAME52888(G52888,G52887,G52886);
  or GNAME52889(G52889,G52568,G57892);
  or GNAME52890(G52890,G57886,G52569);
  nand GNAME52891(G52891,G52890,G52889);
  or GNAME52892(G52892,G57860,G52545);
  or GNAME52893(G52893,G57918,G52522);
  nand GNAME52894(G52894,G52893,G52892);
  or GNAME52895(G52895,G52570,G57893);
  or GNAME52896(G52896,G57887,G52571);
  nand GNAME52897(G52897,G52896,G52895);
  or GNAME52898(G52898,G57901,G52591);
  or GNAME52899(G52899,G57897,G52594);
  nand GNAME52900(G52900,G52899,G52898);
  or GNAME52901(G52901,G52610,G57882);
  or GNAME52902(G52902,G57894,G52611);
  nand GNAME52903(G52903,G52902,G52901);
  or GNAME52904(G52904,G57903,G52598);
  or GNAME52905(G52905,G57898,G52605);
  nand GNAME52906(G52906,G52905,G52904);
  or GNAME52907(G52907,G52612,G57883);
  or GNAME52908(G52908,G57895,G52613);
  nand GNAME52909(G52909,G52908,G52907);
  or GNAME52910(G52910,G57905,G52602);
  or GNAME52911(G52911,G57899,G52608);
  nand GNAME52912(G52912,G52911,G52910);
  or GNAME52913(G52913,G52614,G57884);
  or GNAME52914(G52914,G57896,G52615);
  nand GNAME52915(G52915,G52914,G52913);
  or GNAME52916(G52916,G57873,G52593);
  or GNAME52917(G52917,G57924,G52616);
  nand GNAME52918(G52918,G52917,G52916);
  or GNAME52919(G52919,G52611,G57882);
  or GNAME52920(G52920,G57894,G52649);
  nand GNAME52921(G52921,G52920,G52919);
  or GNAME52922(G52922,G57874,G52604);
  or GNAME52923(G52923,G57925,G52617);
  nand GNAME52924(G52924,G52923,G52922);
  or GNAME52925(G52925,G52613,G57883);
  or GNAME52926(G52926,G57895,G52653);
  nand GNAME52927(G52927,G52926,G52925);
  or GNAME52928(G52928,G57875,G52607);
  or GNAME52929(G52929,G57926,G52618);
  nand GNAME52930(G52930,G52929,G52928);
  or GNAME52931(G52931,G52615,G57884);
  or GNAME52932(G52932,G57896,G52655);
  nand GNAME52933(G52933,G52932,G52931);
  or GNAME52934(G52934,G57901,G52634);
  or GNAME52935(G52935,G57897,G52622);
  nand GNAME52936(G52936,G52935,G52934);
  or GNAME52937(G52937,G52649,G57882);
  or GNAME52938(G52938,G57894,G52650);
  nand GNAME52939(G52939,G52938,G52937);
  or GNAME52940(G52940,G57903,G52640);
  or GNAME52941(G52941,G57898,G52625);
  nand GNAME52942(G52942,G52941,G52940);
  or GNAME52943(G52943,G52653,G57883);
  or GNAME52944(G52944,G57895,G52654);
  nand GNAME52945(G52945,G52944,G52943);
  or GNAME52946(G52946,G57905,G52644);
  or GNAME52947(G52947,G57899,G52626);
  nand GNAME52948(G52948,G52947,G52946);
  or GNAME52949(G52949,G52655,G57884);
  or GNAME52950(G52950,G57896,G52656);
  nand GNAME52951(G52951,G52950,G52949);
  or GNAME52952(G52952,G57936,G52632);
  or GNAME52953(G52953,G57942,G52619);
  nand GNAME52954(G52954,G52953,G52952);
  or GNAME52955(G52955,G52650,G57882);
  or GNAME52956(G52956,G57894,G52651);
  nand GNAME52957(G52957,G52956,G52955);
  or GNAME52958(G52958,G57937,G52638);
  or GNAME52959(G52959,G57943,G52620);
  nand GNAME52960(G52960,G52959,G52958);
  or GNAME52961(G52961,G52654,G57883);
  or GNAME52962(G52962,G57895,G52657);
  nand GNAME52963(G52963,G52962,G52961);
  or GNAME52964(G52964,G57938,G52642);
  or GNAME52965(G52965,G57944,G52621);
  nand GNAME52966(G52966,G52965,G52964);
  or GNAME52967(G52967,G52656,G57884);
  or GNAME52968(G52968,G57896,G52659);
  nand GNAME52969(G52969,G52968,G52967);
  or GNAME52970(G52970,G57901,G52635);
  or GNAME52971(G52971,G57897,G52669);
  nand GNAME52972(G52972,G52971,G52970);
  or GNAME52973(G52973,G52651,G57882);
  or GNAME52974(G52974,G57894,G52652);
  nand GNAME52975(G52975,G52974,G52973);
  or GNAME52976(G52976,G57903,G52645);
  or GNAME52977(G52977,G57898,G52673);
  nand GNAME52978(G52978,G52977,G52976);
  or GNAME52979(G52979,G52657,G57883);
  or GNAME52980(G52980,G57895,G52658);
  nand GNAME52981(G52981,G52980,G52979);
  or GNAME52982(G52982,G57905,G52646);
  or GNAME52983(G52983,G57899,G52677);
  nand GNAME52984(G52984,G52983,G52982);
  or GNAME52985(G52985,G52659,G57884);
  or GNAME52986(G52986,G57896,G52660);
  nand GNAME52987(G52987,G52986,G52985);
  or GNAME52988(G52988,G57939,G52636);
  or GNAME52989(G52989,G57948,G52661);
  nand GNAME52990(G52990,G52989,G52988);
  or GNAME52991(G52991,G52652,G57882);
  or GNAME52992(G52992,G57894,G52686);
  nand GNAME52993(G52993,G52992,G52991);
  or GNAME52994(G52994,G57940,G52647);
  or GNAME52995(G52995,G57949,G52662);
  nand GNAME52996(G52996,G52995,G52994);
  or GNAME52997(G52997,G52658,G57883);
  or GNAME52998(G52998,G57895,G52687);
  nand GNAME52999(G52999,G52998,G52997);
  or GNAME53000(G53000,G57941,G52648);
  or GNAME53001(G53001,G57950,G52663);
  nand GNAME53002(G53002,G53001,G53000);
  or GNAME53003(G53003,G52660,G57884);
  or GNAME53004(G53004,G57896,G52688);
  nand GNAME53005(G53005,G53004,G53003);
  or GNAME53006(G53006,G57901,G52670);
  or GNAME53007(G53007,G57897,G52679);
  nand GNAME53008(G53008,G53007,G53006);
  or GNAME53009(G53009,G52686,G57882);
  or GNAME53010(G53010,G57894,G52685);
  nand GNAME53011(G53011,G53010,G53009);
  or GNAME53012(G53012,G57903,G52674);
  or GNAME53013(G53013,G57898,G52681);
  nand GNAME53014(G53014,G53013,G53012);
  or GNAME53015(G53015,G52687,G57883);
  or GNAME53016(G53016,G57895,G52689);
  nand GNAME53017(G53017,G53016,G53015);
  or GNAME53018(G53018,G57905,G52678);
  or GNAME53019(G53019,G57899,G52683);
  nand GNAME53020(G53020,G53019,G53018);
  or GNAME53021(G53021,G52688,G57884);
  or GNAME53022(G53022,G57896,G52690);
  nand GNAME53023(G53023,G53022,G53021);
  or GNAME53024(G53024,G57900,G52680);
  or GNAME53025(G53025,G57945,G52664);
  nand GNAME53026(G53026,G53025,G53024);
  or GNAME53027(G53027,G57951,G51042);
  or GNAME53028(G53028,G57933,G54659);
  nand GNAME53029(G53029,G53028,G53027);
  or GNAME53030(G53030,G57902,G52682);
  or GNAME53031(G53031,G57946,G52665);
  nand GNAME53032(G53032,G53031,G53030);
  or GNAME53033(G53033,G57952,G51045);
  or GNAME53034(G53034,G57934,G54656);
  nand GNAME53035(G53035,G53034,G53033);
  or GNAME53036(G53036,G57904,G52684);
  or GNAME53037(G53037,G57947,G52666);
  nand GNAME53038(G53038,G53037,G53036);
  or GNAME53039(G53039,G57953,G51048);
  or GNAME53040(G53040,G57935,G54657);
  nand GNAME53041(G53041,G53040,G53039);
  or GNAME53042(G53042,G57901,G52691);
  or GNAME53043(G53043,G57897,G52692);
  nand GNAME53044(G53044,G53043,G53042);
  or GNAME53045(G53045,G52697,G57882);
  or GNAME53046(G53046,G57894,G52698);
  nand GNAME53047(G53047,G53046,G53045);
  or GNAME53048(G53048,G57903,G52693);
  or GNAME53049(G53049,G57898,G52694);
  nand GNAME53050(G53050,G53049,G53048);
  or GNAME53051(G53051,G52699,G57883);
  or GNAME53052(G53052,G57895,G52700);
  nand GNAME53053(G53053,G53052,G53051);
  or GNAME53054(G53054,G57905,G52695);
  or GNAME53055(G53055,G57899,G52696);
  nand GNAME53056(G53056,G53055,G53054);
  or GNAME53057(G53057,G52701,G57884);
  or GNAME53058(G53058,G57896,G52702);
  nand GNAME53059(G53059,G53058,G53057);
  or GNAME53060(G53060,G52703,G57882);
  or GNAME53061(G53061,G57894,G52704);
  nand GNAME53062(G53062,G53061,G53060);
  or GNAME53063(G53063,G52705,G57883);
  or GNAME53064(G53064,G57895,G52706);
  nand GNAME53065(G53065,G53064,G53063);
  or GNAME53066(G53066,G52707,G57884);
  or GNAME53067(G53067,G57896,G52708);
  nand GNAME53068(G53068,G53067,G53066);
  or GNAME53069(G53069,G52704,G57882);
  or GNAME53070(G53070,G57894,G52709);
  nand GNAME53071(G53071,G53070,G53069);
  or GNAME53072(G53072,G52706,G57883);
  or GNAME53073(G53073,G57895,G52710);
  nand GNAME53074(G53074,G53073,G53072);
  or GNAME53075(G53075,G52708,G57884);
  or GNAME53076(G53076,G57896,G52711);
  nand GNAME53077(G53077,G53076,G53075);
  or GNAME53078(G53078,G51051,G57891);
  or GNAME53079(G53079,G57885,G54662);
  nand GNAME53080(G53080,G53079,G53078);
  or GNAME53081(G53081,G51054,G57892);
  or GNAME53082(G53082,G57886,G54663);
  nand GNAME53083(G53083,G53082,G53081);
  or GNAME53084(G53084,G51057,G57893);
  or GNAME53085(G53085,G57887,G54664);
  nand GNAME53086(G53086,G53085,G53084);
  or GNAME53087(G53087,G57901,G52692);
  or GNAME53088(G53088,G57897,G52712);
  nand GNAME53089(G53089,G53088,G53087);
  or GNAME53090(G53090,G57903,G52694);
  or GNAME53091(G53091,G57898,G52713);
  nand GNAME53092(G53092,G53091,G53090);
  or GNAME53093(G53093,G57905,G52696);
  or GNAME53094(G53094,G57899,G52714);
  nand GNAME53095(G53095,G53094,G53093);
  or GNAME53096(G53096,G57921,G54640);
  or GNAME53097(G53097,G57853,G52139);
  nand GNAME53098(G53098,G53097,G53096);
  or GNAME53099(G53099,G57922,G54639);
  or GNAME53100(G53100,G57854,G52141);
  nand GNAME53101(G53101,G53100,G53099);
  or GNAME53102(G53102,G57923,G54641);
  or GNAME53103(G53103,G57855,G52143);
  nand GNAME53104(G53104,G53103,G53102);
  or GNAME53105(G53105,G57927,G54642);
  or GNAME53106(G53106,G57861,G52146);
  nand GNAME53107(G53107,G53106,G53105);
  or GNAME53108(G53108,G57921,G52140);
  or GNAME53109(G53109,G57853,G52145);
  nand GNAME53110(G53110,G53109,G53108);
  or GNAME53111(G53111,G57928,G54643);
  or GNAME53112(G53112,G57862,G52150);
  nand GNAME53113(G53113,G53112,G53111);
  or GNAME53114(G53114,G57922,G52142);
  or GNAME53115(G53115,G57854,G52149);
  nand GNAME53116(G53116,G53115,G53114);
  or GNAME53117(G53117,G57929,G54644);
  or GNAME53118(G53118,G57863,G52154);
  nand GNAME53119(G53119,G53118,G53117);
  or GNAME53120(G53120,G57923,G52144);
  or GNAME53121(G53121,G57855,G52153);
  nand GNAME53122(G53122,G53121,G53120);
  or GNAME53123(G53123,G57921,G52145);
  or GNAME53124(G53124,G57853,G52148);
  nand GNAME53125(G53125,G53124,G53123);
  or GNAME53126(G53126,G57922,G52149);
  or GNAME53127(G53127,G57854,G52152);
  nand GNAME53128(G53128,G53127,G53126);
  or GNAME53129(G53129,G57923,G52153);
  or GNAME53130(G53130,G57855,G52156);
  nand GNAME53131(G53131,G53130,G53129);
  or GNAME53132(G53132,G57921,G52148);
  or GNAME53133(G53133,G57853,G52165);
  nand GNAME53134(G53134,G53133,G53132);
  or GNAME53135(G53135,G57922,G52152);
  or GNAME53136(G53136,G57854,G52170);
  nand GNAME53137(G53137,G53136,G53135);
  or GNAME53138(G53138,G57923,G52156);
  or GNAME53139(G53139,G57855,G52171);
  nand GNAME53140(G53140,G53139,G53138);
  or GNAME53141(G53141,G57876,G54647);
  or GNAME53142(G53142,G57867,G52164);
  nand GNAME53143(G53143,G53142,G53141);
  or GNAME53144(G53144,G57927,G52147);
  or GNAME53145(G53145,G57861,G52163);
  nand GNAME53146(G53146,G53145,G53144);
  or GNAME53147(G53147,G57878,G54649);
  or GNAME53148(G53148,G57869,G52167);
  nand GNAME53149(G53149,G53148,G53147);
  or GNAME53150(G53150,G57928,G52151);
  or GNAME53151(G53151,G57862,G52166);
  nand GNAME53152(G53152,G53151,G53150);
  or GNAME53153(G53153,G57879,G54650);
  or GNAME53154(G53154,G57870,G52169);
  nand GNAME53155(G53155,G53154,G53153);
  or GNAME53156(G53156,G57929,G52155);
  or GNAME53157(G53157,G57863,G52168);
  nand GNAME53158(G53158,G53157,G53156);
  or GNAME53159(G53159,G57921,G52165);
  or GNAME53160(G53160,G57853,G52157);
  nand GNAME53161(G53161,G53160,G53159);
  or GNAME53162(G53162,G57927,G52163);
  or GNAME53163(G53163,G57861,G52158);
  nand GNAME53164(G53164,G53163,G53162);
  or GNAME53165(G53165,G57922,G52170);
  or GNAME53166(G53166,G57854,G52159);
  nand GNAME53167(G53167,G53166,G53165);
  or GNAME53168(G53168,G57928,G52166);
  or GNAME53169(G53169,G57862,G52160);
  nand GNAME53170(G53170,G53169,G53168);
  or GNAME53171(G53171,G57923,G52171);
  or GNAME53172(G53172,G57855,G52161);
  nand GNAME53173(G53173,G53172,G53171);
  or GNAME53174(G53174,G57929,G52168);
  or GNAME53175(G53175,G57863,G52162);
  nand GNAME53176(G53176,G53175,G53174);
  or GNAME53177(G53177,G57877,G54648);
  or GNAME53178(G53178,G57868,G52174);
  nand GNAME53179(G53179,G53178,G53177);
  or GNAME53180(G53180,G57876,G52172);
  or GNAME53181(G53181,G57867,G52173);
  nand GNAME53182(G53182,G53181,G53180);
  or GNAME53183(G53183,G57880,G54651);
  or GNAME53184(G53184,G57871,G52179);
  nand GNAME53185(G53185,G53184,G53183);
  or GNAME53186(G53186,G57878,G52177);
  or GNAME53187(G53187,G57869,G52178);
  nand GNAME53188(G53188,G53187,G53186);
  or GNAME53189(G53189,G57881,G54652);
  or GNAME53190(G53190,G57872,G52182);
  nand GNAME53191(G53191,G53190,G53189);
  or GNAME53192(G53192,G57879,G52180);
  or GNAME53193(G53193,G57870,G52181);
  nand GNAME53194(G53194,G53193,G53192);
  or GNAME53195(G53195,G57927,G52158);
  or GNAME53196(G53196,G57861,G52176);
  nand GNAME53197(G53197,G53196,G53195);
  or GNAME53198(G53198,G57921,G52157);
  or GNAME53199(G53199,G57853,G52175);
  nand GNAME53200(G53200,G53199,G53198);
  or GNAME53201(G53201,G57928,G52160);
  or GNAME53202(G53202,G57862,G52184);
  nand GNAME53203(G53203,G53202,G53201);
  or GNAME53204(G53204,G57922,G52159);
  or GNAME53205(G53205,G57854,G52183);
  nand GNAME53206(G53206,G53205,G53204);
  or GNAME53207(G53207,G57929,G52162);
  or GNAME53208(G53208,G57863,G52186);
  nand GNAME53209(G53209,G53208,G53207);
  or GNAME53210(G53210,G57923,G52161);
  or GNAME53211(G53211,G57855,G52185);
  nand GNAME53212(G53212,G53211,G53210);
  or GNAME53213(G53213,G57954,G54653);
  or GNAME53214(G53214,G57930,G52191);
  nand GNAME53215(G53215,G53214,G53213);
  or GNAME53216(G53216,G57877,G52204);
  or GNAME53217(G53217,G57868,G52205);
  nand GNAME53218(G53218,G53217,G53216);
  or GNAME53219(G53219,G57955,G54654);
  or GNAME53220(G53220,G57931,G52199);
  nand GNAME53221(G53221,G53220,G53219);
  or GNAME53222(G53222,G57880,G52208);
  or GNAME53223(G53223,G57871,G52209);
  nand GNAME53224(G53224,G53223,G53222);
  or GNAME53225(G53225,G57956,G54655);
  or GNAME53226(G53226,G57932,G52201);
  nand GNAME53227(G53227,G53226,G53225);
  or GNAME53228(G53228,G57881,G52212);
  or GNAME53229(G53229,G57872,G52213);
  nand GNAME53230(G53230,G53229,G53228);
  or GNAME53231(G53231,G57877,G52174);
  or GNAME53232(G53232,G57868,G52204);
  nand GNAME53233(G53233,G53232,G53231);
  or GNAME53234(G53234,G57880,G52179);
  or GNAME53235(G53235,G57871,G52208);
  nand GNAME53236(G53236,G53235,G53234);
  or GNAME53237(G53237,G57881,G52182);
  or GNAME53238(G53238,G57872,G52212);
  nand GNAME53239(G53239,G53238,G53237);
  or GNAME53240(G53240,G57921,G52188);
  or GNAME53241(G53241,G57853,G52203);
  nand GNAME53242(G53242,G53241,G53240);
  or GNAME53243(G53243,G57927,G52189);
  or GNAME53244(G53244,G57861,G52190);
  nand GNAME53245(G53245,G53244,G53243);
  or GNAME53246(G53246,G57876,G52187);
  or GNAME53247(G53247,G57867,G52202);
  nand GNAME53248(G53248,G53247,G53246);
  or GNAME53249(G53249,G57922,G52193);
  or GNAME53250(G53250,G57854,G52207);
  nand GNAME53251(G53251,G53250,G53249);
  or GNAME53252(G53252,G57928,G52194);
  or GNAME53253(G53253,G57862,G52198);
  nand GNAME53254(G53254,G53253,G53252);
  or GNAME53255(G53255,G57878,G52192);
  or GNAME53256(G53256,G57869,G52206);
  nand GNAME53257(G53257,G53256,G53255);
  or GNAME53258(G53258,G57923,G52196);
  or GNAME53259(G53259,G57855,G52211);
  nand GNAME53260(G53260,G53259,G53258);
  or GNAME53261(G53261,G57929,G52197);
  or GNAME53262(G53262,G57863,G52200);
  nand GNAME53263(G53263,G53262,G53261);
  or GNAME53264(G53264,G57879,G52195);
  or GNAME53265(G53265,G57870,G52210);
  nand GNAME53266(G53266,G53265,G53264);
  or GNAME53267(G53267,G57927,G52176);
  or GNAME53268(G53268,G57861,G52189);
  nand GNAME53269(G53269,G53268,G53267);
  or GNAME53270(G53270,G57921,G52175);
  or GNAME53271(G53271,G57853,G52188);
  nand GNAME53272(G53272,G53271,G53270);
  or GNAME53273(G53273,G57928,G52184);
  or GNAME53274(G53274,G57862,G52194);
  nand GNAME53275(G53275,G53274,G53273);
  or GNAME53276(G53276,G57922,G52183);
  or GNAME53277(G53277,G57854,G52193);
  nand GNAME53278(G53278,G53277,G53276);
  or GNAME53279(G53279,G57929,G52186);
  or GNAME53280(G53280,G57863,G52197);
  nand GNAME53281(G53281,G53280,G53279);
  or GNAME53282(G53282,G57923,G52185);
  or GNAME53283(G53283,G57855,G52196);
  nand GNAME53284(G53284,G53283,G53282);
  or GNAME53285(G53285,G57876,G52202);
  or GNAME53286(G53286,G57867,G52219);
  nand GNAME53287(G53287,G53286,G53285);
  or GNAME53288(G53288,G57921,G52203);
  or GNAME53289(G53289,G57853,G52218);
  nand GNAME53290(G53290,G53289,G53288);
  or GNAME53291(G53291,G57878,G52206);
  or GNAME53292(G53292,G57869,G52229);
  nand GNAME53293(G53293,G53292,G53291);
  or GNAME53294(G53294,G57922,G52207);
  or GNAME53295(G53295,G57854,G52228);
  nand GNAME53296(G53296,G53295,G53294);
  or GNAME53297(G53297,G57879,G52210);
  or GNAME53298(G53298,G57870,G52232);
  nand GNAME53299(G53299,G53298,G53297);
  or GNAME53300(G53300,G57923,G52211);
  or GNAME53301(G53301,G57855,G52231);
  nand GNAME53302(G53302,G53301,G53300);
  or GNAME53303(G53303,G57954,G52191);
  or GNAME53304(G53304,G57930,G52220);
  nand GNAME53305(G53305,G53304,G53303);
  or GNAME53306(G53306,G57927,G52190);
  or GNAME53307(G53307,G57861,G52214);
  nand GNAME53308(G53308,G53307,G53306);
  or GNAME53309(G53309,G57955,G52199);
  or GNAME53310(G53310,G57931,G52233);
  nand GNAME53311(G53311,G53310,G53309);
  or GNAME53312(G53312,G57928,G52198);
  or GNAME53313(G53313,G57862,G52215);
  nand GNAME53314(G53314,G53313,G53312);
  or GNAME53315(G53315,G57956,G52201);
  or GNAME53316(G53316,G57932,G52240);
  nand GNAME53317(G53317,G53316,G53315);
  or GNAME53318(G53318,G57929,G52200);
  or GNAME53319(G53319,G57863,G52216);
  nand GNAME53320(G53320,G53319,G53318);
  or GNAME53321(G53321,G57951,G54659);
  or GNAME53322(G53322,G57933,G52222);
  nand GNAME53323(G53323,G53322,G53321);
  or GNAME53324(G53324,G57954,G52220);
  or GNAME53325(G53325,G57930,G52221);
  nand GNAME53326(G53326,G53325,G53324);
  or GNAME53327(G53327,G57952,G54656);
  or GNAME53328(G53328,G57934,G52235);
  nand GNAME53329(G53329,G53328,G53327);
  or GNAME53330(G53330,G57955,G52233);
  or GNAME53331(G53331,G57931,G52234);
  nand GNAME53332(G53332,G53331,G53330);
  or GNAME53333(G53333,G57953,G54657);
  or GNAME53334(G53334,G57935,G52242);
  nand GNAME53335(G53335,G53334,G53333);
  or GNAME53336(G53336,G57956,G52240);
  or GNAME53337(G53337,G57932,G52241);
  nand GNAME53338(G53338,G53337,G53336);
  or GNAME53339(G53339,G57877,G52217);
  or GNAME53340(G53340,G57868,G52225);
  nand GNAME53341(G53341,G53340,G53339);
  or GNAME53342(G53342,G57921,G52218);
  or GNAME53343(G53343,G57853,G52224);
  nand GNAME53344(G53344,G53343,G53342);
  or GNAME53345(G53345,G57876,G52219);
  or GNAME53346(G53346,G57867,G52223);
  nand GNAME53347(G53347,G53346,G53345);
  or GNAME53348(G53348,G57880,G52227);
  or GNAME53349(G53349,G57871,G52238);
  nand GNAME53350(G53350,G53349,G53348);
  or GNAME53351(G53351,G57922,G52228);
  or GNAME53352(G53352,G57854,G52237);
  nand GNAME53353(G53353,G53352,G53351);
  or GNAME53354(G53354,G57878,G52229);
  or GNAME53355(G53355,G57869,G52236);
  nand GNAME53356(G53356,G53355,G53354);
  or GNAME53357(G53357,G57881,G52230);
  or GNAME53358(G53358,G57872,G52245);
  nand GNAME53359(G53359,G53358,G53357);
  or GNAME53360(G53360,G57923,G52231);
  or GNAME53361(G53361,G57855,G52244);
  nand GNAME53362(G53362,G53361,G53360);
  or GNAME53363(G53363,G57879,G52232);
  or GNAME53364(G53364,G57870,G52243);
  nand GNAME53365(G53365,G53364,G53363);
  or GNAME53366(G53366,G57876,G52223);
  or GNAME53367(G53367,G57867,G52252);
  nand GNAME53368(G53368,G53367,G53366);
  or GNAME53369(G53369,G57927,G52226);
  or GNAME53370(G53370,G57861,G52251);
  nand GNAME53371(G53371,G53370,G53369);
  or GNAME53372(G53372,G57878,G52236);
  or GNAME53373(G53373,G57869,G52265);
  nand GNAME53374(G53374,G53373,G53372);
  or GNAME53375(G53375,G57928,G52239);
  or GNAME53376(G53376,G57862,G52264);
  nand GNAME53377(G53377,G53376,G53375);
  or GNAME53378(G53378,G57879,G52243);
  or GNAME53379(G53379,G57870,G52271);
  nand GNAME53380(G53380,G53379,G53378);
  or GNAME53381(G53381,G57929,G52246);
  or GNAME53382(G53382,G57863,G52270);
  nand GNAME53383(G53383,G53382,G53381);
  or GNAME53384(G53384,G57927,G52214);
  or GNAME53385(G53385,G57861,G52226);
  nand GNAME53386(G53386,G53385,G53384);
  or GNAME53387(G53387,G57928,G52215);
  or GNAME53388(G53388,G57862,G52239);
  nand GNAME53389(G53389,G53388,G53387);
  or GNAME53390(G53390,G57929,G52216);
  or GNAME53391(G53391,G57863,G52246);
  nand GNAME53392(G53392,G53391,G53390);
  or GNAME53393(G53393,G57951,G52222);
  or GNAME53394(G53394,G57933,G52249);
  nand GNAME53395(G53395,G53394,G53393);
  or GNAME53396(G53396,G57921,G52224);
  or GNAME53397(G53397,G57915,G52248);
  nand GNAME53398(G53398,G53397,G53396);
  or GNAME53399(G53399,G57954,G52221);
  or GNAME53400(G53400,G57930,G52247);
  nand GNAME53401(G53401,G53400,G53399);
  or GNAME53402(G53402,G57954,G52247);
  or GNAME53403(G53403,G57930,G52255);
  nand GNAME53404(G53404,G53403,G53402);
  or GNAME53405(G53405,G57876,G52252);
  or GNAME53406(G53406,G57867,G52254);
  nand GNAME53407(G53407,G53406,G53405);
  or GNAME53408(G53408,G57877,G52250);
  or GNAME53409(G53409,G57868,G52253);
  nand GNAME53410(G53410,G53409,G53408);
  or GNAME53411(G53411,G57952,G52235);
  or GNAME53412(G53412,G57934,G52262);
  nand GNAME53413(G53413,G53412,G53411);
  or GNAME53414(G53414,G57922,G52237);
  or GNAME53415(G53415,G57917,G52261);
  nand GNAME53416(G53416,G53415,G53414);
  or GNAME53417(G53417,G57955,G52234);
  or GNAME53418(G53418,G57931,G52260);
  nand GNAME53419(G53419,G53418,G53417);
  or GNAME53420(G53420,G57953,G52242);
  or GNAME53421(G53421,G57935,G52268);
  nand GNAME53422(G53422,G53421,G53420);
  or GNAME53423(G53423,G57923,G52244);
  or GNAME53424(G53424,G57918,G52267);
  nand GNAME53425(G53425,G53424,G53423);
  or GNAME53426(G53426,G57956,G52241);
  or GNAME53427(G53427,G57932,G52266);
  nand GNAME53428(G53428,G53427,G53426);
  or GNAME53429(G53429,G57955,G52260);
  or GNAME53430(G53430,G57931,G52274);
  nand GNAME53431(G53431,G53430,G53429);
  or GNAME53432(G53432,G57878,G52265);
  or GNAME53433(G53433,G57869,G52273);
  nand GNAME53434(G53434,G53433,G53432);
  or GNAME53435(G53435,G57880,G52263);
  or GNAME53436(G53436,G57871,G52272);
  nand GNAME53437(G53437,G53436,G53435);
  or GNAME53438(G53438,G57956,G52266);
  or GNAME53439(G53439,G57932,G52281);
  nand GNAME53440(G53440,G53439,G53438);
  or GNAME53441(G53441,G57879,G52271);
  or GNAME53442(G53442,G57870,G52280);
  nand GNAME53443(G53443,G53442,G53441);
  or GNAME53444(G53444,G57881,G52269);
  or GNAME53445(G53445,G57872,G52279);
  nand GNAME53446(G53446,G53445,G53444);
  or GNAME53447(G53447,G57951,G52249);
  or GNAME53448(G53448,G57933,G52258);
  nand GNAME53449(G53449,G53448,G53447);
  or GNAME53450(G53450,G57858,G52248);
  or GNAME53451(G53451,G57915,G52257);
  nand GNAME53452(G53452,G53451,G53450);
  or GNAME53453(G53453,G57927,G52251);
  or GNAME53454(G53454,G57861,G52256);
  nand GNAME53455(G53455,G53454,G53453);
  or GNAME53456(G53456,G57952,G52262);
  or GNAME53457(G53457,G57934,G52277);
  nand GNAME53458(G53458,G53457,G53456);
  or GNAME53459(G53459,G57859,G52261);
  or GNAME53460(G53460,G57917,G52276);
  nand GNAME53461(G53461,G53460,G53459);
  or GNAME53462(G53462,G57928,G52264);
  or GNAME53463(G53463,G57862,G52275);
  nand GNAME53464(G53464,G53463,G53462);
  or GNAME53465(G53465,G57953,G52268);
  or GNAME53466(G53466,G57935,G52284);
  nand GNAME53467(G53467,G53466,G53465);
  or GNAME53468(G53468,G57860,G52267);
  or GNAME53469(G53469,G57918,G52283);
  nand GNAME53470(G53470,G53469,G53468);
  or GNAME53471(G53471,G57929,G52270);
  or GNAME53472(G53472,G57863,G52282);
  nand GNAME53473(G53473,G53472,G53471);
  or GNAME53474(G53474,G57877,G52253);
  or GNAME53475(G53475,G57868,G52287);
  nand GNAME53476(G53476,G53475,G53474);
  or GNAME53477(G53477,G57858,G52257);
  or GNAME53478(G53478,G57915,G52286);
  nand GNAME53479(G53479,G53478,G53477);
  or GNAME53480(G53480,G57880,G52272);
  or GNAME53481(G53481,G57871,G52301);
  nand GNAME53482(G53482,G53481,G53480);
  or GNAME53483(G53483,G57859,G52276);
  or GNAME53484(G53484,G57917,G52300);
  nand GNAME53485(G53485,G53484,G53483);
  or GNAME53486(G53486,G57881,G52279);
  or GNAME53487(G53487,G57872,G52308);
  nand GNAME53488(G53488,G53487,G53486);
  or GNAME53489(G53489,G57860,G52283);
  or GNAME53490(G53490,G57918,G52307);
  nand GNAME53491(G53491,G53490,G53489);
  or GNAME53492(G53492,G57954,G52291);
  or GNAME53493(G53493,G57930,G52295);
  nand GNAME53494(G53494,G53493,G53492);
  or GNAME53495(G53495,G57876,G52289);
  or GNAME53496(G53496,G57867,G52294);
  nand GNAME53497(G53497,G53496,G53495);
  or GNAME53498(G53498,G57877,G52287);
  or GNAME53499(G53499,G57868,G52293);
  nand GNAME53500(G53500,G53499,G53498);
  or GNAME53501(G53501,G57955,G52305);
  or GNAME53502(G53502,G57931,G52316);
  nand GNAME53503(G53503,G53502,G53501);
  or GNAME53504(G53504,G57878,G52303);
  or GNAME53505(G53505,G57869,G52315);
  nand GNAME53506(G53506,G53505,G53504);
  or GNAME53507(G53507,G57880,G52301);
  or GNAME53508(G53508,G57871,G52314);
  nand GNAME53509(G53509,G53508,G53507);
  or GNAME53510(G53510,G57956,G52312);
  or GNAME53511(G53511,G57932,G52323);
  nand GNAME53512(G53512,G53511,G53510);
  or GNAME53513(G53513,G57879,G52310);
  or GNAME53514(G53514,G57870,G52322);
  nand GNAME53515(G53515,G53514,G53513);
  or GNAME53516(G53516,G57881,G52308);
  or GNAME53517(G53517,G57872,G52321);
  nand GNAME53518(G53518,G53517,G53516);
  or GNAME53519(G53519,G57906,G52290);
  or GNAME53520(G53520,G57888,G52299);
  nand GNAME53521(G53521,G53520,G53519);
  or GNAME53522(G53522,G54662,G57891);
  or GNAME53523(G53523,G57885,G52328);
  nand GNAME53524(G53524,G53523,G53522);
  or GNAME53525(G53525,G57907,G52304);
  or GNAME53526(G53526,G57889,G52320);
  nand GNAME53527(G53527,G53526,G53525);
  or GNAME53528(G53528,G54663,G57892);
  or GNAME53529(G53529,G57886,G52329);
  nand GNAME53530(G53530,G53529,G53528);
  or GNAME53531(G53531,G57908,G52311);
  or GNAME53532(G53532,G57890,G52327);
  nand GNAME53533(G53533,G53532,G53531);
  or GNAME53534(G53534,G54664,G57893);
  or GNAME53535(G53535,G57887,G52330);
  nand GNAME53536(G53536,G53535,G53534);
  or GNAME53537(G53537,G57927,G52256);
  or GNAME53538(G53538,G57916,G52292);
  nand GNAME53539(G53539,G53538,G53537);
  or GNAME53540(G53540,G57954,G52255);
  or GNAME53541(G53541,G57930,G52291);
  nand GNAME53542(G53542,G53541,G53540);
  or GNAME53543(G53543,G57928,G52275);
  or GNAME53544(G53544,G57919,G52306);
  nand GNAME53545(G53545,G53544,G53543);
  or GNAME53546(G53546,G57955,G52274);
  or GNAME53547(G53547,G57931,G52305);
  nand GNAME53548(G53548,G53547,G53546);
  or GNAME53549(G53549,G57929,G52282);
  or GNAME53550(G53550,G57920,G52313);
  nand GNAME53551(G53551,G53550,G53549);
  or GNAME53552(G53552,G57956,G52281);
  or GNAME53553(G53553,G57932,G52312);
  nand GNAME53554(G53554,G53553,G53552);
  or GNAME53555(G53555,G57906,G52259);
  or GNAME53556(G53556,G57888,G52290);
  nand GNAME53557(G53557,G53556,G53555);
  or GNAME53558(G53558,G57876,G52254);
  or GNAME53559(G53559,G57867,G52289);
  nand GNAME53560(G53560,G53559,G53558);
  or GNAME53561(G53561,G57951,G52258);
  or GNAME53562(G53562,G57933,G52288);
  nand GNAME53563(G53563,G53562,G53561);
  or GNAME53564(G53564,G57951,G52288);
  or GNAME53565(G53565,G57933,G52298);
  nand GNAME53566(G53566,G53565,G53564);
  or GNAME53567(G53567,G57858,G52286);
  or GNAME53568(G53568,G57915,G52297);
  nand GNAME53569(G53569,G53568,G53567);
  or GNAME53570(G53570,G57864,G52292);
  or GNAME53571(G53571,G57916,G52296);
  nand GNAME53572(G53572,G53571,G53570);
  or GNAME53573(G53573,G57907,G52278);
  or GNAME53574(G53574,G57889,G52304);
  nand GNAME53575(G53575,G53574,G53573);
  or GNAME53576(G53576,G57878,G52273);
  or GNAME53577(G53577,G57869,G52303);
  nand GNAME53578(G53578,G53577,G53576);
  or GNAME53579(G53579,G57952,G52277);
  or GNAME53580(G53580,G57934,G52302);
  nand GNAME53581(G53581,G53580,G53579);
  or GNAME53582(G53582,G57908,G52285);
  or GNAME53583(G53583,G57890,G52311);
  nand GNAME53584(G53584,G53583,G53582);
  or GNAME53585(G53585,G57879,G52280);
  or GNAME53586(G53586,G57870,G52310);
  nand GNAME53587(G53587,G53586,G53585);
  or GNAME53588(G53588,G57953,G52284);
  or GNAME53589(G53589,G57935,G52309);
  nand GNAME53590(G53590,G53589,G53588);
  or GNAME53591(G53591,G57952,G52302);
  or GNAME53592(G53592,G57934,G52319);
  nand GNAME53593(G53593,G53592,G53591);
  or GNAME53594(G53594,G57859,G52300);
  or GNAME53595(G53595,G57917,G52318);
  nand GNAME53596(G53596,G53595,G53594);
  or GNAME53597(G53597,G57865,G52306);
  or GNAME53598(G53598,G57919,G52317);
  nand GNAME53599(G53599,G53598,G53597);
  or GNAME53600(G53600,G57953,G52309);
  or GNAME53601(G53601,G57935,G52326);
  nand GNAME53602(G53602,G53601,G53600);
  or GNAME53603(G53603,G57860,G52307);
  or GNAME53604(G53604,G57918,G52325);
  nand GNAME53605(G53605,G53604,G53603);
  or GNAME53606(G53606,G57866,G52313);
  or GNAME53607(G53607,G57920,G52324);
  nand GNAME53608(G53608,G53607,G53606);
  or GNAME53609(G53609,G57954,G52295);
  or GNAME53610(G53610,G57930,G52333);
  nand GNAME53611(G53611,G53610,G53609);
  or GNAME53612(G53612,G57876,G52294);
  or GNAME53613(G53613,G57924,G52332);
  nand GNAME53614(G53614,G53613,G53612);
  or GNAME53615(G53615,G57877,G52293);
  or GNAME53616(G53616,G57868,G52331);
  nand GNAME53617(G53617,G53616,G53615);
  or GNAME53618(G53618,G57954,G52333);
  or GNAME53619(G53619,G57930,G52340);
  nand GNAME53620(G53620,G53619,G53618);
  or GNAME53621(G53621,G57873,G52332);
  or GNAME53622(G53622,G57924,G52339);
  nand GNAME53623(G53623,G53622,G53621);
  or GNAME53624(G53624,G57877,G52331);
  or GNAME53625(G53625,G57868,G52338);
  nand GNAME53626(G53626,G53625,G53624);
  or GNAME53627(G53627,G57955,G52316);
  or GNAME53628(G53628,G57931,G52347);
  nand GNAME53629(G53629,G53628,G53627);
  or GNAME53630(G53630,G57878,G52315);
  or GNAME53631(G53631,G57925,G52346);
  nand GNAME53632(G53632,G53631,G53630);
  or GNAME53633(G53633,G57880,G52314);
  or GNAME53634(G53634,G57871,G52345);
  nand GNAME53635(G53635,G53634,G53633);
  or GNAME53636(G53636,G57956,G52323);
  or GNAME53637(G53637,G57932,G52354);
  nand GNAME53638(G53638,G53637,G53636);
  or GNAME53639(G53639,G57879,G52322);
  or GNAME53640(G53640,G57926,G52353);
  nand GNAME53641(G53641,G53640,G53639);
  or GNAME53642(G53642,G57881,G52321);
  or GNAME53643(G53643,G57872,G52352);
  nand GNAME53644(G53644,G53643,G53642);
  or GNAME53645(G53645,G57955,G52347);
  or GNAME53646(G53646,G57931,G52361);
  nand GNAME53647(G53647,G53646,G53645);
  or GNAME53648(G53648,G57874,G52346);
  or GNAME53649(G53649,G57925,G52360);
  nand GNAME53650(G53650,G53649,G53648);
  or GNAME53651(G53651,G57880,G52345);
  or GNAME53652(G53652,G57871,G52359);
  nand GNAME53653(G53653,G53652,G53651);
  or GNAME53654(G53654,G57956,G52354);
  or GNAME53655(G53655,G57932,G52368);
  nand GNAME53656(G53656,G53655,G53654);
  or GNAME53657(G53657,G57875,G52353);
  or GNAME53658(G53658,G57926,G52367);
  nand GNAME53659(G53659,G53658,G53657);
  or GNAME53660(G53660,G57881,G52352);
  or GNAME53661(G53661,G57872,G52366);
  nand GNAME53662(G53662,G53661,G53660);
  or GNAME53663(G53663,G57906,G52299);
  or GNAME53664(G53664,G57888,G52337);
  nand GNAME53665(G53665,G53664,G53663);
  or GNAME53666(G53666,G52328,G57891);
  or GNAME53667(G53667,G57885,G52373);
  nand GNAME53668(G53668,G53667,G53666);
  or GNAME53669(G53669,G57906,G52337);
  or GNAME53670(G53670,G57888,G52344);
  nand GNAME53671(G53671,G53670,G53669);
  or GNAME53672(G53672,G52373,G57891);
  or GNAME53673(G53673,G57885,G52374);
  nand GNAME53674(G53674,G53673,G53672);
  or GNAME53675(G53675,G57907,G52320);
  or GNAME53676(G53676,G57889,G52351);
  nand GNAME53677(G53677,G53676,G53675);
  or GNAME53678(G53678,G52329,G57892);
  or GNAME53679(G53679,G57886,G52375);
  nand GNAME53680(G53680,G53679,G53678);
  or GNAME53681(G53681,G57908,G52327);
  or GNAME53682(G53682,G57890,G52358);
  nand GNAME53683(G53683,G53682,G53681);
  or GNAME53684(G53684,G52330,G57893);
  or GNAME53685(G53685,G57887,G52376);
  nand GNAME53686(G53686,G53685,G53684);
  or GNAME53687(G53687,G57907,G52351);
  or GNAME53688(G53688,G57889,G52365);
  nand GNAME53689(G53689,G53688,G53687);
  or GNAME53690(G53690,G52375,G57892);
  or GNAME53691(G53691,G57886,G52377);
  nand GNAME53692(G53692,G53691,G53690);
  or GNAME53693(G53693,G57908,G52358);
  or GNAME53694(G53694,G57890,G52372);
  nand GNAME53695(G53695,G53694,G53693);
  or GNAME53696(G53696,G52376,G57893);
  or GNAME53697(G53697,G57887,G52378);
  nand GNAME53698(G53698,G53697,G53696);
  or GNAME53699(G53699,G57951,G52298);
  or GNAME53700(G53700,G57933,G52336);
  nand GNAME53701(G53701,G53700,G53699);
  or GNAME53702(G53702,G57858,G52297);
  or GNAME53703(G53703,G57915,G52335);
  nand GNAME53704(G53704,G53703,G53702);
  or GNAME53705(G53705,G57864,G52296);
  or GNAME53706(G53706,G57916,G52334);
  nand GNAME53707(G53707,G53706,G53705);
  or GNAME53708(G53708,G57951,G52336);
  or GNAME53709(G53709,G57933,G52343);
  nand GNAME53710(G53710,G53709,G53708);
  or GNAME53711(G53711,G57858,G52335);
  or GNAME53712(G53712,G57915,G52342);
  nand GNAME53713(G53713,G53712,G53711);
  or GNAME53714(G53714,G57864,G52334);
  or GNAME53715(G53715,G57916,G52341);
  nand GNAME53716(G53716,G53715,G53714);
  or GNAME53717(G53717,G57952,G52319);
  or GNAME53718(G53718,G57934,G52350);
  nand GNAME53719(G53719,G53718,G53717);
  or GNAME53720(G53720,G57859,G52318);
  or GNAME53721(G53721,G57917,G52349);
  nand GNAME53722(G53722,G53721,G53720);
  or GNAME53723(G53723,G57865,G52317);
  or GNAME53724(G53724,G57919,G52348);
  nand GNAME53725(G53725,G53724,G53723);
  or GNAME53726(G53726,G57953,G52326);
  or GNAME53727(G53727,G57935,G52357);
  nand GNAME53728(G53728,G53727,G53726);
  or GNAME53729(G53729,G57860,G52325);
  or GNAME53730(G53730,G57918,G52356);
  nand GNAME53731(G53731,G53730,G53729);
  or GNAME53732(G53732,G57866,G52324);
  or GNAME53733(G53733,G57920,G52355);
  nand GNAME53734(G53734,G53733,G53732);
  or GNAME53735(G53735,G57952,G52350);
  or GNAME53736(G53736,G57934,G52364);
  nand GNAME53737(G53737,G53736,G53735);
  or GNAME53738(G53738,G57859,G52349);
  or GNAME53739(G53739,G57917,G52363);
  nand GNAME53740(G53740,G53739,G53738);
  or GNAME53741(G53741,G57865,G52348);
  or GNAME53742(G53742,G57919,G52362);
  nand GNAME53743(G53743,G53742,G53741);
  or GNAME53744(G53744,G57953,G52357);
  or GNAME53745(G53745,G57935,G52371);
  nand GNAME53746(G53746,G53745,G53744);
  or GNAME53747(G53747,G57860,G52356);
  or GNAME53748(G53748,G57918,G52370);
  nand GNAME53749(G53749,G53748,G53747);
  or GNAME53750(G53750,G57866,G52355);
  or GNAME53751(G53751,G57920,G52369);
  nand GNAME53752(G53752,G53751,G53750);
  or GNAME53753(G53753,G57954,G52340);
  or GNAME53754(G53754,G57930,G52381);
  nand GNAME53755(G53755,G53754,G53753);
  or GNAME53756(G53756,G57873,G52339);
  or GNAME53757(G53757,G57924,G52380);
  nand GNAME53758(G53758,G53757,G53756);
  or GNAME53759(G53759,G57877,G52338);
  or GNAME53760(G53760,G57942,G52379);
  nand GNAME53761(G53761,G53760,G53759);
  or GNAME53762(G53762,G57954,G52381);
  or GNAME53763(G53763,G57930,G52388);
  nand GNAME53764(G53764,G53763,G53762);
  or GNAME53765(G53765,G57873,G52380);
  or GNAME53766(G53766,G57924,G52387);
  nand GNAME53767(G53767,G53766,G53765);
  or GNAME53768(G53768,G57936,G52379);
  or GNAME53769(G53769,G57942,G52386);
  nand GNAME53770(G53770,G53769,G53768);
  or GNAME53771(G53771,G57955,G52361);
  or GNAME53772(G53772,G57931,G52395);
  nand GNAME53773(G53773,G53772,G53771);
  or GNAME53774(G53774,G57874,G52360);
  or GNAME53775(G53775,G57925,G52394);
  nand GNAME53776(G53776,G53775,G53774);
  or GNAME53777(G53777,G57880,G52359);
  or GNAME53778(G53778,G57943,G52393);
  nand GNAME53779(G53779,G53778,G53777);
  or GNAME53780(G53780,G57956,G52368);
  or GNAME53781(G53781,G57932,G52402);
  nand GNAME53782(G53782,G53781,G53780);
  or GNAME53783(G53783,G57875,G52367);
  or GNAME53784(G53784,G57926,G52401);
  nand GNAME53785(G53785,G53784,G53783);
  or GNAME53786(G53786,G57881,G52366);
  or GNAME53787(G53787,G57944,G52400);
  nand GNAME53788(G53788,G53787,G53786);
  or GNAME53789(G53789,G57955,G52395);
  or GNAME53790(G53790,G57931,G52409);
  nand GNAME53791(G53791,G53790,G53789);
  or GNAME53792(G53792,G57874,G52394);
  or GNAME53793(G53793,G57925,G52408);
  nand GNAME53794(G53794,G53793,G53792);
  or GNAME53795(G53795,G57937,G52393);
  or GNAME53796(G53796,G57943,G52407);
  nand GNAME53797(G53797,G53796,G53795);
  or GNAME53798(G53798,G57956,G52402);
  or GNAME53799(G53799,G57932,G52416);
  nand GNAME53800(G53800,G53799,G53798);
  or GNAME53801(G53801,G57875,G52401);
  or GNAME53802(G53802,G57926,G52415);
  nand GNAME53803(G53803,G53802,G53801);
  or GNAME53804(G53804,G57938,G52400);
  or GNAME53805(G53805,G57944,G52414);
  nand GNAME53806(G53806,G53805,G53804);
  or GNAME53807(G53807,G57906,G52344);
  or GNAME53808(G53808,G57888,G52385);
  nand GNAME53809(G53809,G53808,G53807);
  or GNAME53810(G53810,G52374,G57891);
  or GNAME53811(G53811,G57885,G52421);
  nand GNAME53812(G53812,G53811,G53810);
  or GNAME53813(G53813,G57906,G52385);
  or GNAME53814(G53814,G57888,G52392);
  nand GNAME53815(G53815,G53814,G53813);
  or GNAME53816(G53816,G52421,G57891);
  or GNAME53817(G53817,G57885,G52422);
  nand GNAME53818(G53818,G53817,G53816);
  or GNAME53819(G53819,G57907,G52365);
  or GNAME53820(G53820,G57889,G52399);
  nand GNAME53821(G53821,G53820,G53819);
  or GNAME53822(G53822,G52377,G57892);
  or GNAME53823(G53823,G57886,G52423);
  nand GNAME53824(G53824,G53823,G53822);
  or GNAME53825(G53825,G57908,G52372);
  or GNAME53826(G53826,G57890,G52406);
  nand GNAME53827(G53827,G53826,G53825);
  or GNAME53828(G53828,G52378,G57893);
  or GNAME53829(G53829,G57887,G52424);
  nand GNAME53830(G53830,G53829,G53828);
  or GNAME53831(G53831,G57907,G52399);
  or GNAME53832(G53832,G57889,G52413);
  nand GNAME53833(G53833,G53832,G53831);
  or GNAME53834(G53834,G52423,G57892);
  or GNAME53835(G53835,G57886,G52425);
  nand GNAME53836(G53836,G53835,G53834);
  or GNAME53837(G53837,G57908,G52406);
  or GNAME53838(G53838,G57890,G52420);
  nand GNAME53839(G53839,G53838,G53837);
  or GNAME53840(G53840,G52424,G57893);
  or GNAME53841(G53841,G57887,G52426);
  nand GNAME53842(G53842,G53841,G53840);
  or GNAME53843(G53843,G57951,G52343);
  or GNAME53844(G53844,G57933,G52384);
  nand GNAME53845(G53845,G53844,G53843);
  or GNAME53846(G53846,G57858,G52342);
  or GNAME53847(G53847,G57915,G52383);
  nand GNAME53848(G53848,G53847,G53846);
  or GNAME53849(G53849,G57864,G52341);
  or GNAME53850(G53850,G57916,G52382);
  nand GNAME53851(G53851,G53850,G53849);
  or GNAME53852(G53852,G57951,G52384);
  or GNAME53853(G53853,G57933,G52391);
  nand GNAME53854(G53854,G53853,G53852);
  or GNAME53855(G53855,G57858,G52383);
  or GNAME53856(G53856,G57915,G52390);
  nand GNAME53857(G53857,G53856,G53855);
  or GNAME53858(G53858,G57864,G52382);
  or GNAME53859(G53859,G57916,G52389);
  nand GNAME53860(G53860,G53859,G53858);
  or GNAME53861(G53861,G57952,G52364);
  or GNAME53862(G53862,G57934,G52398);
  nand GNAME53863(G53863,G53862,G53861);
  or GNAME53864(G53864,G57859,G52363);
  or GNAME53865(G53865,G57917,G52397);
  nand GNAME53866(G53866,G53865,G53864);
  or GNAME53867(G53867,G57865,G52362);
  or GNAME53868(G53868,G57919,G52396);
  nand GNAME53869(G53869,G53868,G53867);
  or GNAME53870(G53870,G57953,G52371);
  or GNAME53871(G53871,G57935,G52405);
  nand GNAME53872(G53872,G53871,G53870);
  or GNAME53873(G53873,G57860,G52370);
  or GNAME53874(G53874,G57918,G52404);
  nand GNAME53875(G53875,G53874,G53873);
  or GNAME53876(G53876,G57866,G52369);
  or GNAME53877(G53877,G57920,G52403);
  nand GNAME53878(G53878,G53877,G53876);
  or GNAME53879(G53879,G57952,G52398);
  or GNAME53880(G53880,G57934,G52412);
  nand GNAME53881(G53881,G53880,G53879);
  or GNAME53882(G53882,G57859,G52397);
  or GNAME53883(G53883,G57917,G52411);
  nand GNAME53884(G53884,G53883,G53882);
  or GNAME53885(G53885,G57865,G52396);
  or GNAME53886(G53886,G57919,G52410);
  nand GNAME53887(G53887,G53886,G53885);
  or GNAME53888(G53888,G57953,G52405);
  or GNAME53889(G53889,G57935,G52419);
  nand GNAME53890(G53890,G53889,G53888);
  or GNAME53891(G53891,G57860,G52404);
  or GNAME53892(G53892,G57918,G52418);
  nand GNAME53893(G53893,G53892,G53891);
  or GNAME53894(G53894,G57866,G52403);
  or GNAME53895(G53895,G57920,G52417);
  nand GNAME53896(G53896,G53895,G53894);
  or GNAME53897(G53897,G57954,G52388);
  or GNAME53898(G53898,G57948,G52429);
  nand GNAME53899(G53899,G53898,G53897);
  or GNAME53900(G53900,G57873,G52387);
  or GNAME53901(G53901,G57924,G52428);
  nand GNAME53902(G53902,G53901,G53900);
  or GNAME53903(G53903,G57936,G52386);
  or GNAME53904(G53904,G57942,G52427);
  nand GNAME53905(G53905,G53904,G53903);
  or GNAME53906(G53906,G57939,G52429);
  or GNAME53907(G53907,G57948,G52436);
  nand GNAME53908(G53908,G53907,G53906);
  or GNAME53909(G53909,G57873,G52428);
  or GNAME53910(G53910,G57924,G52435);
  nand GNAME53911(G53911,G53910,G53909);
  or GNAME53912(G53912,G57936,G52427);
  or GNAME53913(G53913,G57942,G52434);
  nand GNAME53914(G53914,G53913,G53912);
  or GNAME53915(G53915,G57955,G52409);
  or GNAME53916(G53916,G57949,G52443);
  nand GNAME53917(G53917,G53916,G53915);
  or GNAME53918(G53918,G57874,G52408);
  or GNAME53919(G53919,G57925,G52442);
  nand GNAME53920(G53920,G53919,G53918);
  or GNAME53921(G53921,G57937,G52407);
  or GNAME53922(G53922,G57943,G52441);
  nand GNAME53923(G53923,G53922,G53921);
  or GNAME53924(G53924,G57956,G52416);
  or GNAME53925(G53925,G57950,G52450);
  nand GNAME53926(G53926,G53925,G53924);
  or GNAME53927(G53927,G57875,G52415);
  or GNAME53928(G53928,G57926,G52449);
  nand GNAME53929(G53929,G53928,G53927);
  or GNAME53930(G53930,G57938,G52414);
  or GNAME53931(G53931,G57944,G52448);
  nand GNAME53932(G53932,G53931,G53930);
  or GNAME53933(G53933,G57940,G52443);
  or GNAME53934(G53934,G57949,G52457);
  nand GNAME53935(G53935,G53934,G53933);
  or GNAME53936(G53936,G57874,G52442);
  or GNAME53937(G53937,G57925,G52456);
  nand GNAME53938(G53938,G53937,G53936);
  or GNAME53939(G53939,G57937,G52441);
  or GNAME53940(G53940,G57943,G52455);
  nand GNAME53941(G53941,G53940,G53939);
  or GNAME53942(G53942,G57941,G52450);
  or GNAME53943(G53943,G57950,G52464);
  nand GNAME53944(G53944,G53943,G53942);
  or GNAME53945(G53945,G57875,G52449);
  or GNAME53946(G53946,G57926,G52463);
  nand GNAME53947(G53947,G53946,G53945);
  or GNAME53948(G53948,G57938,G52448);
  or GNAME53949(G53949,G57944,G52462);
  nand GNAME53950(G53950,G53949,G53948);
  or GNAME53951(G53951,G57906,G52392);
  or GNAME53952(G53952,G57888,G52433);
  nand GNAME53953(G53953,G53952,G53951);
  or GNAME53954(G53954,G52422,G57891);
  or GNAME53955(G53955,G57885,G52469);
  nand GNAME53956(G53956,G53955,G53954);
  or GNAME53957(G53957,G57906,G52433);
  or GNAME53958(G53958,G57888,G52440);
  nand GNAME53959(G53959,G53958,G53957);
  or GNAME53960(G53960,G52469,G57891);
  or GNAME53961(G53961,G57885,G52470);
  nand GNAME53962(G53962,G53961,G53960);
  or GNAME53963(G53963,G57907,G52413);
  or GNAME53964(G53964,G57889,G52447);
  nand GNAME53965(G53965,G53964,G53963);
  or GNAME53966(G53966,G52425,G57892);
  or GNAME53967(G53967,G57886,G52471);
  nand GNAME53968(G53968,G53967,G53966);
  or GNAME53969(G53969,G57908,G52420);
  or GNAME53970(G53970,G57890,G52454);
  nand GNAME53971(G53971,G53970,G53969);
  or GNAME53972(G53972,G52426,G57893);
  or GNAME53973(G53973,G57887,G52472);
  nand GNAME53974(G53974,G53973,G53972);
  or GNAME53975(G53975,G57907,G52447);
  or GNAME53976(G53976,G57889,G52461);
  nand GNAME53977(G53977,G53976,G53975);
  or GNAME53978(G53978,G52471,G57892);
  or GNAME53979(G53979,G57886,G52473);
  nand GNAME53980(G53980,G53979,G53978);
  or GNAME53981(G53981,G57908,G52454);
  or GNAME53982(G53982,G57890,G52468);
  nand GNAME53983(G53983,G53982,G53981);
  or GNAME53984(G53984,G52472,G57893);
  or GNAME53985(G53985,G57887,G52474);
  nand GNAME53986(G53986,G53985,G53984);
  or GNAME53987(G53987,G57951,G52391);
  or GNAME53988(G53988,G57933,G52432);
  nand GNAME53989(G53989,G53988,G53987);
  or GNAME53990(G53990,G57858,G52390);
  or GNAME53991(G53991,G57915,G52431);
  nand GNAME53992(G53992,G53991,G53990);
  or GNAME53993(G53993,G57864,G52389);
  or GNAME53994(G53994,G57916,G52430);
  nand GNAME53995(G53995,G53994,G53993);
  or GNAME53996(G53996,G57951,G52432);
  or GNAME53997(G53997,G57933,G52439);
  nand GNAME53998(G53998,G53997,G53996);
  or GNAME53999(G53999,G57858,G52431);
  or GNAME54000(G54000,G57915,G52438);
  nand GNAME54001(G54001,G54000,G53999);
  or GNAME54002(G54002,G57864,G52430);
  or GNAME54003(G54003,G57916,G52437);
  nand GNAME54004(G54004,G54003,G54002);
  or GNAME54005(G54005,G57952,G52412);
  or GNAME54006(G54006,G57934,G52446);
  nand GNAME54007(G54007,G54006,G54005);
  or GNAME54008(G54008,G57859,G52411);
  or GNAME54009(G54009,G57917,G52445);
  nand GNAME54010(G54010,G54009,G54008);
  or GNAME54011(G54011,G57865,G52410);
  or GNAME54012(G54012,G57919,G52444);
  nand GNAME54013(G54013,G54012,G54011);
  or GNAME54014(G54014,G57953,G52419);
  or GNAME54015(G54015,G57935,G52453);
  nand GNAME54016(G54016,G54015,G54014);
  or GNAME54017(G54017,G57860,G52418);
  or GNAME54018(G54018,G57918,G52452);
  nand GNAME54019(G54019,G54018,G54017);
  or GNAME54020(G54020,G57866,G52417);
  or GNAME54021(G54021,G57920,G52451);
  nand GNAME54022(G54022,G54021,G54020);
  or GNAME54023(G54023,G57952,G52446);
  or GNAME54024(G54024,G57934,G52460);
  nand GNAME54025(G54025,G54024,G54023);
  or GNAME54026(G54026,G57859,G52445);
  or GNAME54027(G54027,G57917,G52459);
  nand GNAME54028(G54028,G54027,G54026);
  or GNAME54029(G54029,G57865,G52444);
  or GNAME54030(G54030,G57919,G52458);
  nand GNAME54031(G54031,G54030,G54029);
  or GNAME54032(G54032,G57953,G52453);
  or GNAME54033(G54033,G57935,G52467);
  nand GNAME54034(G54034,G54033,G54032);
  or GNAME54035(G54035,G57860,G52452);
  or GNAME54036(G54036,G57918,G52466);
  nand GNAME54037(G54037,G54036,G54035);
  or GNAME54038(G54038,G57866,G52451);
  or GNAME54039(G54039,G57920,G52465);
  nand GNAME54040(G54040,G54039,G54038);
  or GNAME54041(G54041,G57939,G52436);
  or GNAME54042(G54042,G57948,G52480);
  nand GNAME54043(G54043,G54042,G54041);
  or GNAME54044(G54044,G57873,G52435);
  or GNAME54045(G54045,G57924,G52479);
  nand GNAME54046(G54046,G54045,G54044);
  or GNAME54047(G54047,G57936,G52434);
  or GNAME54048(G54048,G57942,G52478);
  nand GNAME54049(G54049,G54048,G54047);
  or GNAME54050(G54050,G57939,G52480);
  or GNAME54051(G54051,G57948,G52487);
  nand GNAME54052(G54052,G54051,G54050);
  or GNAME54053(G54053,G57873,G52479);
  or GNAME54054(G54054,G57924,G52486);
  nand GNAME54055(G54055,G54054,G54053);
  or GNAME54056(G54056,G57936,G52478);
  or GNAME54057(G54057,G57942,G52485);
  nand GNAME54058(G54058,G54057,G54056);
  or GNAME54059(G54059,G57940,G52457);
  or GNAME54060(G54060,G57949,G52492);
  nand GNAME54061(G54061,G54060,G54059);
  or GNAME54062(G54062,G57874,G52456);
  or GNAME54063(G54063,G57925,G52491);
  nand GNAME54064(G54064,G54063,G54062);
  or GNAME54065(G54065,G57937,G52455);
  or GNAME54066(G54066,G57943,G52490);
  nand GNAME54067(G54067,G54066,G54065);
  or GNAME54068(G54068,G57941,G52464);
  or GNAME54069(G54069,G57950,G52499);
  nand GNAME54070(G54070,G54069,G54068);
  or GNAME54071(G54071,G57875,G52463);
  or GNAME54072(G54072,G57926,G52498);
  nand GNAME54073(G54073,G54072,G54071);
  or GNAME54074(G54074,G57938,G52462);
  or GNAME54075(G54075,G57944,G52497);
  nand GNAME54076(G54076,G54075,G54074);
  or GNAME54077(G54077,G57940,G52492);
  or GNAME54078(G54078,G57949,G52506);
  nand GNAME54079(G54079,G54078,G54077);
  or GNAME54080(G54080,G57874,G52491);
  or GNAME54081(G54081,G57925,G52505);
  nand GNAME54082(G54082,G54081,G54080);
  or GNAME54083(G54083,G57937,G52490);
  or GNAME54084(G54084,G57943,G52504);
  nand GNAME54085(G54085,G54084,G54083);
  or GNAME54086(G54086,G57941,G52499);
  or GNAME54087(G54087,G57950,G52511);
  nand GNAME54088(G54088,G54087,G54086);
  or GNAME54089(G54089,G57875,G52498);
  or GNAME54090(G54090,G57926,G52510);
  nand GNAME54091(G54091,G54090,G54089);
  or GNAME54092(G54092,G57938,G52497);
  or GNAME54093(G54093,G57944,G52509);
  nand GNAME54094(G54094,G54093,G54092);
  or GNAME54095(G54095,G57906,G52440);
  or GNAME54096(G54096,G57888,G52484);
  nand GNAME54097(G54097,G54096,G54095);
  or GNAME54098(G54098,G52470,G57891);
  or GNAME54099(G54099,G57885,G52514);
  nand GNAME54100(G54100,G54099,G54098);
  or GNAME54101(G54101,G57907,G52461);
  or GNAME54102(G54102,G57889,G52496);
  nand GNAME54103(G54103,G54102,G54101);
  or GNAME54104(G54104,G52473,G57892);
  or GNAME54105(G54105,G57886,G52515);
  nand GNAME54106(G54106,G54105,G54104);
  or GNAME54107(G54107,G57908,G52468);
  or GNAME54108(G54108,G57890,G52503);
  nand GNAME54109(G54109,G54108,G54107);
  or GNAME54110(G54110,G52474,G57893);
  or GNAME54111(G54111,G57887,G52516);
  nand GNAME54112(G54112,G54111,G54110);
  or GNAME54113(G54113,G57951,G52439);
  or GNAME54114(G54114,G57945,G52483);
  nand GNAME54115(G54115,G54114,G54113);
  or GNAME54116(G54116,G57858,G52438);
  or GNAME54117(G54117,G57915,G52482);
  nand GNAME54118(G54118,G54117,G54116);
  or GNAME54119(G54119,G57864,G52437);
  or GNAME54120(G54120,G57916,G52481);
  nand GNAME54121(G54121,G54120,G54119);
  or GNAME54122(G54122,G57900,G52483);
  or GNAME54123(G54123,G57945,G52475);
  nand GNAME54124(G54124,G54123,G54122);
  or GNAME54125(G54125,G57858,G52482);
  or GNAME54126(G54126,G57915,G52526);
  nand GNAME54127(G54127,G54126,G54125);
  or GNAME54128(G54128,G57864,G52481);
  or GNAME54129(G54129,G57916,G52488);
  nand GNAME54130(G54130,G54129,G54128);
  or GNAME54131(G54131,G57952,G52460);
  or GNAME54132(G54132,G57946,G52495);
  nand GNAME54133(G54133,G54132,G54131);
  or GNAME54134(G54134,G57859,G52459);
  or GNAME54135(G54135,G57917,G52494);
  nand GNAME54136(G54136,G54135,G54134);
  or GNAME54137(G54137,G57865,G52458);
  or GNAME54138(G54138,G57919,G52493);
  nand GNAME54139(G54139,G54138,G54137);
  or GNAME54140(G54140,G57953,G52467);
  or GNAME54141(G54141,G57947,G52502);
  nand GNAME54142(G54142,G54141,G54140);
  or GNAME54143(G54143,G57860,G52466);
  or GNAME54144(G54144,G57918,G52501);
  nand GNAME54145(G54145,G54144,G54143);
  or GNAME54146(G54146,G57866,G52465);
  or GNAME54147(G54147,G57920,G52500);
  nand GNAME54148(G54148,G54147,G54146);
  or GNAME54149(G54149,G57902,G52495);
  or GNAME54150(G54150,G57946,G52476);
  nand GNAME54151(G54151,G54150,G54149);
  or GNAME54152(G54152,G57859,G52494);
  or GNAME54153(G54153,G57917,G52539);
  nand GNAME54154(G54154,G54153,G54152);
  or GNAME54155(G54155,G57865,G52493);
  or GNAME54156(G54156,G57919,G52507);
  nand GNAME54157(G54157,G54156,G54155);
  or GNAME54158(G54158,G57904,G52502);
  or GNAME54159(G54159,G57947,G52477);
  nand GNAME54160(G54160,G54159,G54158);
  or GNAME54161(G54161,G57860,G52501);
  or GNAME54162(G54162,G57918,G52545);
  nand GNAME54163(G54163,G54162,G54161);
  or GNAME54164(G54164,G57866,G52500);
  or GNAME54165(G54165,G57920,G52512);
  nand GNAME54166(G54166,G54165,G54164);
  or GNAME54167(G54167,G57873,G52486);
  or GNAME54168(G54168,G57924,G52529);
  nand GNAME54169(G54169,G54168,G54167);
  or GNAME54170(G54170,G57906,G52489);
  or GNAME54171(G54171,G57897,G52528);
  nand GNAME54172(G54172,G54171,G54170);
  or GNAME54173(G54173,G57939,G52487);
  or GNAME54174(G54174,G57948,G52527);
  nand GNAME54175(G54175,G54174,G54173);
  or GNAME54176(G54176,G57874,G52505);
  or GNAME54177(G54177,G57925,G52542);
  nand GNAME54178(G54178,G54177,G54176);
  or GNAME54179(G54179,G57907,G52508);
  or GNAME54180(G54180,G57898,G52541);
  nand GNAME54181(G54181,G54180,G54179);
  or GNAME54182(G54182,G57940,G52506);
  or GNAME54183(G54183,G57949,G52540);
  nand GNAME54184(G54184,G54183,G54182);
  or GNAME54185(G54185,G57875,G52510);
  or GNAME54186(G54186,G57926,G52548);
  nand GNAME54187(G54187,G54186,G54185);
  or GNAME54188(G54188,G57908,G52513);
  or GNAME54189(G54189,G57899,G52547);
  nand GNAME54190(G54190,G54189,G54188);
  or GNAME54191(G54191,G57941,G52511);
  or GNAME54192(G54192,G57950,G52546);
  nand GNAME54193(G54193,G54192,G54191);
  or GNAME54194(G54194,G57939,G52527);
  or GNAME54195(G54195,G57948,G52538);
  nand GNAME54196(G54196,G54195,G54194);
  or GNAME54197(G54197,G57936,G52531);
  or GNAME54198(G54198,G57942,G52537);
  nand GNAME54199(G54199,G54198,G54197);
  or GNAME54200(G54200,G57940,G52540);
  or GNAME54201(G54201,G57949,G52557);
  nand GNAME54202(G54202,G54201,G54200);
  or GNAME54203(G54203,G57937,G52544);
  or GNAME54204(G54204,G57943,G52556);
  nand GNAME54205(G54205,G54204,G54203);
  or GNAME54206(G54206,G57941,G52546);
  or GNAME54207(G54207,G57950,G52564);
  nand GNAME54208(G54208,G54207,G54206);
  or GNAME54209(G54209,G57938,G52550);
  or GNAME54210(G54210,G57944,G52563);
  nand GNAME54211(G54211,G54210,G54209);
  or GNAME54212(G54212,G57900,G52475);
  or GNAME54213(G54213,G57945,G52535);
  nand GNAME54214(G54214,G54213,G54212);
  or GNAME54215(G54215,G57902,G52476);
  or GNAME54216(G54216,G57946,G52554);
  nand GNAME54217(G54217,G54216,G54215);
  or GNAME54218(G54218,G57904,G52477);
  or GNAME54219(G54219,G57947,G52561);
  nand GNAME54220(G54220,G54219,G54218);
  or GNAME54221(G54221,G57936,G52485);
  or GNAME54222(G54222,G57942,G52531);
  nand GNAME54223(G54223,G54222,G54221);
  or GNAME54224(G54224,G57864,G52488);
  or GNAME54225(G54225,G57916,G52530);
  nand GNAME54226(G54226,G54225,G54224);
  or GNAME54227(G54227,G57921,G50988);
  or GNAME54228(G54228,G57853,G54640);
  nand GNAME54229(G54229,G54228,G54227);
  or GNAME54230(G54230,G57900,G52535);
  or GNAME54231(G54231,G57945,G52536);
  nand GNAME54232(G54232,G54231,G54230);
  or GNAME54233(G54233,G57864,G52530);
  or GNAME54234(G54234,G57916,G52534);
  nand GNAME54235(G54235,G54234,G54233);
  or GNAME54236(G54236,G57873,G52529);
  or GNAME54237(G54237,G57924,G52533);
  nand GNAME54238(G54238,G54237,G54236);
  or GNAME54239(G54239,G57937,G52504);
  or GNAME54240(G54240,G57943,G52544);
  nand GNAME54241(G54241,G54240,G54239);
  or GNAME54242(G54242,G57865,G52507);
  or GNAME54243(G54243,G57919,G52543);
  nand GNAME54244(G54244,G54243,G54242);
  or GNAME54245(G54245,G57922,G50991);
  or GNAME54246(G54246,G57854,G54639);
  nand GNAME54247(G54247,G54246,G54245);
  or GNAME54248(G54248,G57938,G52509);
  or GNAME54249(G54249,G57944,G52550);
  nand GNAME54250(G54250,G54249,G54248);
  or GNAME54251(G54251,G57866,G52512);
  or GNAME54252(G54252,G57920,G52549);
  nand GNAME54253(G54253,G54252,G54251);
  or GNAME54254(G54254,G57923,G50994);
  or GNAME54255(G54255,G57855,G54641);
  nand GNAME54256(G54256,G54255,G54254);
  or GNAME54257(G54257,G57902,G52554);
  or GNAME54258(G54258,G57946,G52555);
  nand GNAME54259(G54259,G54258,G54257);
  or GNAME54260(G54260,G57865,G52543);
  or GNAME54261(G54261,G57919,G52553);
  nand GNAME54262(G54262,G54261,G54260);
  or GNAME54263(G54263,G57874,G52542);
  or GNAME54264(G54264,G57925,G52552);
  nand GNAME54265(G54265,G54264,G54263);
  or GNAME54266(G54266,G57904,G52561);
  or GNAME54267(G54267,G57947,G52562);
  nand GNAME54268(G54268,G54267,G54266);
  or GNAME54269(G54269,G57866,G52549);
  or GNAME54270(G54270,G57920,G52560);
  nand GNAME54271(G54271,G54270,G54269);
  or GNAME54272(G54272,G57875,G52548);
  or GNAME54273(G54273,G57926,G52559);
  nand GNAME54274(G54274,G54273,G54272);
  or GNAME54275(G54275,G57936,G52537);
  or GNAME54276(G54276,G57942,G52592);
  nand GNAME54277(G54277,G54276,G54275);
  or GNAME54278(G54278,G57901,G52532);
  or GNAME54279(G54279,G57897,G52591);
  nand GNAME54280(G54280,G54279,G54278);
  or GNAME54281(G54281,G57900,G52536);
  or GNAME54282(G54282,G57945,G52590);
  nand GNAME54283(G54283,G54282,G54281);
  or GNAME54284(G54284,G57900,G52590);
  or GNAME54285(G54285,G57945,G52576);
  nand GNAME54286(G54286,G54285,G54284);
  or GNAME54287(G54287,G57873,G52589);
  or GNAME54288(G54288,G57924,G52593);
  nand GNAME54289(G54289,G54288,G54287);
  or GNAME54290(G54290,G57936,G52592);
  or GNAME54291(G54291,G57942,G52574);
  nand GNAME54292(G54292,G54291,G54290);
  or GNAME54293(G54293,G57937,G52556);
  or GNAME54294(G54294,G57943,G52599);
  nand GNAME54295(G54295,G54294,G54293);
  or GNAME54296(G54296,G57903,G52551);
  or GNAME54297(G54297,G57898,G52598);
  nand GNAME54298(G54298,G54297,G54296);
  or GNAME54299(G54299,G57902,G52555);
  or GNAME54300(G54300,G57946,G52597);
  nand GNAME54301(G54301,G54300,G54299);
  or GNAME54302(G54302,G57938,G52563);
  or GNAME54303(G54303,G57944,G52603);
  nand GNAME54304(G54304,G54303,G54302);
  or GNAME54305(G54305,G57905,G52558);
  or GNAME54306(G54306,G57899,G52602);
  nand GNAME54307(G54307,G54306,G54305);
  or GNAME54308(G54308,G57904,G52562);
  or GNAME54309(G54309,G57947,G52601);
  nand GNAME54310(G54310,G54309,G54308);
  or GNAME54311(G54311,G57902,G52597);
  or GNAME54312(G54312,G57946,G52581);
  nand GNAME54313(G54313,G54312,G54311);
  or GNAME54314(G54314,G57874,G52596);
  or GNAME54315(G54315,G57925,G52604);
  nand GNAME54316(G54316,G54315,G54314);
  or GNAME54317(G54317,G57937,G52599);
  or GNAME54318(G54318,G57943,G52579);
  nand GNAME54319(G54319,G54318,G54317);
  or GNAME54320(G54320,G57904,G52601);
  or GNAME54321(G54321,G57947,G52586);
  nand GNAME54322(G54322,G54321,G54320);
  or GNAME54323(G54323,G57875,G52600);
  or GNAME54324(G54324,G57926,G52607);
  nand GNAME54325(G54325,G54324,G54323);
  or GNAME54326(G54326,G57938,G52603);
  or GNAME54327(G54327,G57944,G52584);
  nand GNAME54328(G54328,G54327,G54326);
  or GNAME54329(G54329,G57939,G52523);
  or GNAME54330(G54330,G57948,G52595);
  nand GNAME54331(G54331,G54330,G54329);
  or GNAME54332(G54332,G57900,G52576);
  or GNAME54333(G54333,G57945,G52577);
  nand GNAME54334(G54334,G54333,G54332);
  or GNAME54335(G54335,G57936,G52574);
  or GNAME54336(G54336,G57942,G52575);
  nand GNAME54337(G54337,G54336,G54335);
  or GNAME54338(G54338,G57940,G52524);
  or GNAME54339(G54339,G57949,G52606);
  nand GNAME54340(G54340,G54339,G54338);
  or GNAME54341(G54341,G57941,G52525);
  or GNAME54342(G54342,G57950,G52609);
  nand GNAME54343(G54343,G54342,G54341);
  or GNAME54344(G54344,G57902,G52581);
  or GNAME54345(G54345,G57946,G52582);
  nand GNAME54346(G54346,G54345,G54344);
  or GNAME54347(G54347,G57937,G52579);
  or GNAME54348(G54348,G57943,G52580);
  nand GNAME54349(G54349,G54348,G54347);
  or GNAME54350(G54350,G57904,G52586);
  or GNAME54351(G54351,G57947,G52587);
  nand GNAME54352(G54352,G54351,G54350);
  or GNAME54353(G54353,G57938,G52584);
  or GNAME54354(G54354,G57944,G52585);
  nand GNAME54355(G54355,G54354,G54353);
  or GNAME54356(G54356,G57939,G52538);
  or GNAME54357(G54357,G57948,G52523);
  nand GNAME54358(G54358,G54357,G54356);
  or GNAME54359(G54359,G57873,G52533);
  or GNAME54360(G54360,G57924,G52589);
  nand GNAME54361(G54361,G54360,G54359);
  or GNAME54362(G54362,G57927,G50997);
  or GNAME54363(G54363,G57861,G54642);
  nand GNAME54364(G54364,G54363,G54362);
  or GNAME54365(G54365,G57940,G52557);
  or GNAME54366(G54366,G57949,G52524);
  nand GNAME54367(G54367,G54366,G54365);
  or GNAME54368(G54368,G57874,G52552);
  or GNAME54369(G54369,G57925,G52596);
  nand GNAME54370(G54370,G54369,G54368);
  or GNAME54371(G54371,G57928,G51000);
  or GNAME54372(G54372,G57862,G54643);
  nand GNAME54373(G54373,G54372,G54371);
  or GNAME54374(G54374,G57941,G52564);
  or GNAME54375(G54375,G57950,G52525);
  nand GNAME54376(G54376,G54375,G54374);
  or GNAME54377(G54377,G57875,G52559);
  or GNAME54378(G54378,G57926,G52600);
  nand GNAME54379(G54379,G54378,G54377);
  or GNAME54380(G54380,G57929,G51003);
  or GNAME54381(G54381,G57863,G54644);
  nand GNAME54382(G54382,G54381,G54380);
  or GNAME54383(G54383,G57939,G52595);
  or GNAME54384(G54384,G57948,G52578);
  nand GNAME54385(G54385,G54384,G54383);
  or GNAME54386(G54386,G57901,G52594);
  or GNAME54387(G54387,G57897,G52634);
  nand GNAME54388(G54388,G54387,G54386);
  or GNAME54389(G54389,G57876,G51006);
  or GNAME54390(G54390,G57867,G54647);
  nand GNAME54391(G54391,G54390,G54389);
  or GNAME54392(G54392,G57940,G52606);
  or GNAME54393(G54393,G57949,G52583);
  nand GNAME54394(G54394,G54393,G54392);
  or GNAME54395(G54395,G57903,G52605);
  or GNAME54396(G54396,G57898,G52640);
  nand GNAME54397(G54397,G54396,G54395);
  or GNAME54398(G54398,G57878,G51009);
  or GNAME54399(G54399,G57869,G54649);
  nand GNAME54400(G54400,G54399,G54398);
  or GNAME54401(G54401,G57941,G52609);
  or GNAME54402(G54402,G57950,G52588);
  nand GNAME54403(G54403,G54402,G54401);
  or GNAME54404(G54404,G57905,G52608);
  or GNAME54405(G54405,G57899,G52644);
  nand GNAME54406(G54406,G54405,G54404);
  or GNAME54407(G54407,G57879,G51012);
  or GNAME54408(G54408,G57870,G54650);
  nand GNAME54409(G54409,G54408,G54407);
  or GNAME54410(G54410,G57939,G52631);
  or GNAME54411(G54411,G57948,G52623);
  nand GNAME54412(G54412,G54411,G54410);
  or GNAME54413(G54413,G57900,G52633);
  or GNAME54414(G54414,G57945,G52624);
  nand GNAME54415(G54415,G54414,G54413);
  or GNAME54416(G54416,G57877,G51015);
  or GNAME54417(G54417,G57868,G54648);
  nand GNAME54418(G54418,G54417,G54416);
  or GNAME54419(G54419,G57940,G52637);
  or GNAME54420(G54420,G57949,G52627);
  nand GNAME54421(G54421,G54420,G54419);
  or GNAME54422(G54422,G57902,G52639);
  or GNAME54423(G54423,G57946,G52628);
  nand GNAME54424(G54424,G54423,G54422);
  or GNAME54425(G54425,G57880,G51018);
  or GNAME54426(G54426,G57871,G54651);
  nand GNAME54427(G54427,G54426,G54425);
  or GNAME54428(G54428,G57941,G52641);
  or GNAME54429(G54429,G57950,G52629);
  nand GNAME54430(G54430,G54429,G54428);
  or GNAME54431(G54431,G57904,G52643);
  or GNAME54432(G54432,G57947,G52630);
  nand GNAME54433(G54433,G54432,G54431);
  or GNAME54434(G54434,G57881,G51021);
  or GNAME54435(G54435,G57872,G54652);
  nand GNAME54436(G54436,G54435,G54434);
  or GNAME54437(G54437,G57900,G52577);
  or GNAME54438(G54438,G57945,G52633);
  nand GNAME54439(G54439,G54438,G54437);
  or GNAME54440(G54440,G57936,G52575);
  or GNAME54441(G54441,G57942,G52632);
  nand GNAME54442(G54442,G54441,G54440);
  or GNAME54443(G54443,G57939,G52578);
  or GNAME54444(G54444,G57948,G52631);
  nand GNAME54445(G54445,G54444,G54443);
  or GNAME54446(G54446,G57902,G52582);
  or GNAME54447(G54447,G57946,G52639);
  nand GNAME54448(G54448,G54447,G54446);
  or GNAME54449(G54449,G57937,G52580);
  or GNAME54450(G54450,G57943,G52638);
  nand GNAME54451(G54451,G54450,G54449);
  or GNAME54452(G54452,G57940,G52583);
  or GNAME54453(G54453,G57949,G52637);
  nand GNAME54454(G54454,G54453,G54452);
  or GNAME54455(G54455,G57904,G52587);
  or GNAME54456(G54456,G57947,G52643);
  nand GNAME54457(G54457,G54456,G54455);
  or GNAME54458(G54458,G57938,G52585);
  or GNAME54459(G54459,G57944,G52642);
  nand GNAME54460(G54460,G54459,G54458);
  or GNAME54461(G54461,G57941,G52588);
  or GNAME54462(G54462,G57950,G52641);
  nand GNAME54463(G54463,G54462,G54461);
  or GNAME54464(G54464,G57901,G52669);
  or GNAME54465(G54465,G57897,G52670);
  nand GNAME54466(G54466,G54465,G54464);
  or GNAME54467(G54467,G57900,G52668);
  or GNAME54468(G54468,G57945,G52667);
  nand GNAME54469(G54469,G54468,G54467);
  or GNAME54470(G54470,G57954,G51024);
  or GNAME54471(G54471,G57930,G54653);
  nand GNAME54472(G54472,G54471,G54470);
  or GNAME54473(G54473,G57903,G52673);
  or GNAME54474(G54474,G57898,G52674);
  nand GNAME54475(G54475,G54474,G54473);
  or GNAME54476(G54476,G57902,G52671);
  or GNAME54477(G54477,G57946,G52672);
  nand GNAME54478(G54478,G54477,G54476);
  or GNAME54479(G54479,G57955,G51027);
  or GNAME54480(G54480,G57931,G54654);
  nand GNAME54481(G54481,G54480,G54479);
  or GNAME54482(G54482,G57905,G52677);
  or GNAME54483(G54483,G57899,G52678);
  nand GNAME54484(G54484,G54483,G54482);
  or GNAME54485(G54485,G57904,G52675);
  or GNAME54486(G54486,G57947,G52676);
  nand GNAME54487(G54487,G54486,G54485);
  or GNAME54488(G54488,G57956,G51030);
  or GNAME54489(G54489,G57932,G54655);
  nand GNAME54490(G54490,G54489,G54488);
  or GNAME54491(G54491,G57900,G52624);
  or GNAME54492(G54492,G57945,G52668);
  nand GNAME54493(G54493,G54492,G54491);
  or GNAME54494(G54494,G57939,G52623);
  or GNAME54495(G54495,G57948,G52636);
  nand GNAME54496(G54496,G54495,G54494);
  or GNAME54497(G54497,G57902,G52628);
  or GNAME54498(G54498,G57946,G52671);
  nand GNAME54499(G54499,G54498,G54497);
  or GNAME54500(G54500,G57940,G52627);
  or GNAME54501(G54501,G57949,G52647);
  nand GNAME54502(G54502,G54501,G54500);
  or GNAME54503(G54503,G57904,G52630);
  or GNAME54504(G54504,G57947,G52675);
  nand GNAME54505(G54505,G54504,G54503);
  or GNAME54506(G54506,G57941,G52629);
  or GNAME54507(G54507,G57950,G52648);
  nand GNAME54508(G54508,G54507,G54506);
  or GNAME54509(G54509,G57901,G52622);
  or GNAME54510(G54510,G57897,G52635);
  nand GNAME54511(G54511,G54510,G54509);
  or GNAME54512(G54512,G57903,G52625);
  or GNAME54513(G54513,G57898,G52645);
  nand GNAME54514(G54514,G54513,G54512);
  or GNAME54515(G54515,G57905,G52626);
  or GNAME54516(G54516,G57899,G52646);
  nand GNAME54517(G54517,G54516,G54515);
  or GNAME54518(G54518,G57900,G52667);
  or GNAME54519(G54519,G57945,G52680);
  nand GNAME54520(G54520,G54519,G54518);
  or GNAME54521(G54521,G57902,G52672);
  or GNAME54522(G54522,G57946,G52682);
  nand GNAME54523(G54523,G54522,G54521);
  or GNAME54524(G54524,G57904,G52676);
  or GNAME54525(G54525,G57947,G52684);
  nand GNAME54526(G54526,G54525,G54524);
  or GNAME54527(G54527,G57906,G51033);
  or GNAME54528(G54528,G57888,G54658);
  nand GNAME54529(G54529,G54528,G54527);
  or GNAME54530(G54530,G57907,G51036);
  or GNAME54531(G54531,G57889,G54660);
  nand GNAME54532(G54532,G54531,G54530);
  or GNAME54533(G54533,G57908,G51039);
  or GNAME54534(G54534,G57890,G54661);
  nand GNAME54535(G54535,G54534,G54533);
  or GNAME54536(G54536,G57901,G52679);
  or GNAME54537(G54537,G57897,G52691);
  nand GNAME54538(G54538,G54537,G54536);
  or GNAME54539(G54539,G52685,G57882);
  or GNAME54540(G54540,G57894,G52697);
  nand GNAME54541(G54541,G54540,G54539);
  or GNAME54542(G54542,G57903,G52681);
  or GNAME54543(G54543,G57898,G52693);
  nand GNAME54544(G54544,G54543,G54542);
  or GNAME54545(G54545,G52689,G57883);
  or GNAME54546(G54546,G57895,G52699);
  nand GNAME54547(G54547,G54546,G54545);
  or GNAME54548(G54548,G57905,G52683);
  or GNAME54549(G54549,G57899,G52695);
  nand GNAME54550(G54550,G54549,G54548);
  or GNAME54551(G54551,G52690,G57884);
  or GNAME54552(G54552,G57896,G52701);
  nand GNAME54553(G54553,G54552,G54551);
  or GNAME54554(G54554,G52698,G57882);
  or GNAME54555(G54555,G57894,G52703);
  nand GNAME54556(G54556,G54555,G54554);
  or GNAME54557(G54557,G52700,G57883);
  or GNAME54558(G54558,G57895,G52705);
  nand GNAME54559(G54559,G54558,G54557);
  or GNAME54560(G54560,G52702,G57884);
  or GNAME54561(G54561,G57896,G52707);
  nand GNAME54562(G54562,G54561,G54560);
  not GNAME54563(G54563,G55990);
  not GNAME54564(G54564,G54755);
  not GNAME54565(G54565,G54768);
  not GNAME54566(G54566,G2344);
  not GNAME54567(G54567,G1928);
  not GNAME54568(G54568,G1512);
  not GNAME54569(G54569,G57724);
  not GNAME54570(G54570,G57729);
  not GNAME54571(G54571,G57728);
  not GNAME54572(G54572,G57730);
  not GNAME54573(G54573,G57738);
  not GNAME54574(G54574,G57737);
  not GNAME54575(G54575,G57739);
  not GNAME54576(G54576,G57734);
  not GNAME54577(G54577,G57735);
  not GNAME54578(G54578,G57736);
  not GNAME54579(G54579,G57746);
  not GNAME54580(G54580,G57747);
  not GNAME54581(G54581,G57748);
  not GNAME54582(G54582,G57743);
  not GNAME54583(G54583,G57744);
  not GNAME54584(G54584,G57745);
  not GNAME54585(G54585,G57755);
  not GNAME54586(G54586,G57756);
  not GNAME54587(G54587,G57757);
  not GNAME54588(G54588,G57752);
  not GNAME54589(G54589,G57753);
  not GNAME54590(G54590,G57754);
  not GNAME54591(G54591,G57764);
  not GNAME54592(G54592,G57765);
  not GNAME54593(G54593,G57766);
  not GNAME54594(G54594,G57761);
  not GNAME54595(G54595,G57762);
  not GNAME54596(G54596,G57763);
  not GNAME54597(G54597,G57771);
  not GNAME54598(G54598,G57773);
  not GNAME54599(G54599,G57775);
  not GNAME54600(G54600,G57770);
  not GNAME54601(G54601,G57772);
  not GNAME54602(G54602,G57774);
  not GNAME54603(G54603,G57789);
  not GNAME54604(G54604,G57792);
  not GNAME54605(G54605,G57794);
  not GNAME54606(G54606,G57808);
  not GNAME54607(G54607,G57810);
  not GNAME54608(G54608,G57812);
  not GNAME54609(G54609,G57790);
  not GNAME54610(G54610,G57793);
  not GNAME54611(G54611,G57795);
  not GNAME54612(G54612,G57791);
  not GNAME54613(G54613,G57796);
  not GNAME54614(G54614,G57797);
  not GNAME54615(G54615,G57813);
  not GNAME54616(G54616,G57814);
  not GNAME54617(G54617,G57815);
  not GNAME54618(G54618,G57807);
  not GNAME54619(G54619,G57822);
  not GNAME54620(G54620,G57809);
  not GNAME54621(G54621,G57811);
  not GNAME54622(G54622,G57823);
  not GNAME54623(G54623,G57824);
  not GNAME54624(G54624,G57819);
  not GNAME54625(G54625,G57820);
  not GNAME54626(G54626,G57827);
  not GNAME54627(G54627,G57830);
  not GNAME54628(G54628,G57826);
  not GNAME54629(G54629,G57829);
  not GNAME54630(G54630,G57821);
  not GNAME54631(G54631,G57840);
  not GNAME54632(G54632,G57825);
  not GNAME54633(G54633,G57828);
  not GNAME54634(G54634,G57842);
  not GNAME54635(G54635,G57844);
  not GNAME54636(G54636,G57841);
  not GNAME54637(G54637,G57843);
  not GNAME54638(G54638,G57845);
  not GNAME54639(G54639,G57782);
  not GNAME54640(G54640,G57781);
  not GNAME54641(G54641,G57783);
  not GNAME54642(G54642,G57784);
  not GNAME54643(G54643,G57785);
  not GNAME54644(G54644,G57786);
  not GNAME54645(G54645,G57787);
  not GNAME54646(G54646,G57788);
  not GNAME54647(G54647,G57801);
  not GNAME54648(G54648,G57816);
  not GNAME54649(G54649,G57802);
  not GNAME54650(G54650,G57803);
  not GNAME54651(G54651,G57817);
  not GNAME54652(G54652,G57818);
  not GNAME54653(G54653,G57831);
  not GNAME54654(G54654,G57832);
  not GNAME54655(G54655,G57833);
  not GNAME54656(G54656,G57835);
  not GNAME54657(G54657,G57836);
  not GNAME54658(G54658,G57846);
  not GNAME54659(G54659,G57834);
  not GNAME54660(G54660,G57847);
  not GNAME54661(G54661,G57848);
  not GNAME54662(G54662,G57849);
  not GNAME54663(G54663,G57850);
  not GNAME54664(G54664,G57851);
  not GNAME54665(G54665,G52049);
  not GNAME54666(G54666,G52048);
  not GNAME54667(G54667,G52050);
  not GNAME54668(G54668,G52054);
  not GNAME54669(G54669,G52055);
  not GNAME54670(G54670,G52056);
  not GNAME54671(G54671,G52060);
  not GNAME54672(G54672,G52061);
  not GNAME54673(G54673,G52062);
  not GNAME54674(G54674,G52066);
  not GNAME54675(G54675,G52067);
  not GNAME54676(G54676,G52068);
  not GNAME54677(G54677,G52072);
  not GNAME54678(G54678,G52073);
  not GNAME54679(G54679,G52074);
  not GNAME54680(G54680,G52078);
  not GNAME54681(G54681,G52079);
  not GNAME54682(G54682,G52080);
  not GNAME54683(G54683,G52087);
  not GNAME54684(G54684,G52088);
  not GNAME54685(G54685,G52089);
  nand GNAME54686(G54686,G52118,G54715);
  nand GNAME54687(G54687,G52119,G54716);
  nand GNAME54688(G54688,G52120,G54717);
  nand GNAME54689(G54689,G52121,G54718);
  nand GNAME54690(G54690,G52122,G54719);
  nand GNAME54691(G54691,G52123,G54720);
  nand GNAME54692(G54692,G52124,G54721);
  nand GNAME54693(G54693,G52125,G54722);
  nand GNAME54694(G54694,G52126,G54723);
  nand GNAME54695(G54695,G52127,G54724);
  nand GNAME54696(G54696,G52128,G54725);
  nand GNAME54697(G54697,G52129,G54726);
  nand GNAME54698(G54698,G52133,G54727);
  nand GNAME54699(G54699,G52130,G54728);
  nand GNAME54700(G54700,G52131,G54729);
  nand GNAME54701(G54701,G52132,G54730);
  nand GNAME54702(G54702,G52134,G54731);
  nand GNAME54703(G54703,G52135,G54732);
  nand GNAME54704(G54704,G54733,G54566);
  nand GNAME54705(G54705,G54734,G54567);
  nand GNAME54706(G54706,G54735,G54568);
  nand GNAME54707(G54707,G52136,G54736);
  nand GNAME54708(G54708,G52137,G54737);
  nand GNAME54709(G54709,G52138,G54738);
  xor GNAME54710(G54710,G54833,G54807);
  xor GNAME54711(G54711,G51728,G57576);
  xor GNAME54712(G54712,G51710,G57563);
  xor GNAME54713(G54713,G51716,G57589);
  xor GNAME54714(G54714,G57719,G49328);
  xor GNAME54715(G54715,G2678,G2699);
  xor GNAME54716(G54716,G2262,G2283);
  xor GNAME54717(G54717,G1846,G1867);
  xor GNAME54718(G54718,G2636,G2657);
  xor GNAME54719(G54719,G2220,G2241);
  xor GNAME54720(G54720,G1804,G1825);
  xor GNAME54721(G54721,G2552,G2573);
  xor GNAME54722(G54722,G2136,G2157);
  xor GNAME54723(G54723,G1720,G1741);
  xor GNAME54724(G54724,G2594,G2615);
  xor GNAME54725(G54725,G2178,G2199);
  xor GNAME54726(G54726,G1762,G1783);
  xor GNAME54727(G54727,G2428,G2449);
  xor GNAME54728(G54728,G2470,G2491);
  xor GNAME54729(G54729,G2054,G2075);
  xor GNAME54730(G54730,G1638,G1659);
  xor GNAME54731(G54731,G2012,G2033);
  xor GNAME54732(G54732,G1596,G1617);
  xor GNAME54733(G54733,G2344,G2365);
  xor GNAME54734(G54734,G1928,G1949);
  xor GNAME54735(G54735,G1512,G1533);
  xor GNAME54736(G54736,G2386,G2407);
  xor GNAME54737(G54737,G1970,G1991);
  xor GNAME54738(G54738,G1554,G1575);
  xor GNAME54739(G54739,G50984,G50987);
  xor GNAME54740(G54740,G41048,G51060);
  xor GNAME54741(G54741,G47303,G54740);
  xor GNAME54742(G54742,G41033,G51062);
  xor GNAME54743(G54743,G47288,G54742);
  xor GNAME54744(G54744,G41063,G51064);
  xor GNAME54745(G54745,G47318,G54744);
  dff DFF_54754(CK,G54753,G47268);
  and GNAME54755(G54755,G54753,G54756);
  nand GNAME54756(G54756,G80,G54758);
  buf GNAME54757(G54757,G54753);
  buf GNAME54758(G54758,G54748);
  dff DFF_54767(CK,G54766,G47253);
  and GNAME54768(G54768,G54766,G54769);
  nand GNAME54769(G54769,G80,G54771);
  buf GNAME54770(G54770,G54766);
  buf GNAME54771(G54771,G54761);
  dff DFF_54780(CK,G54779,G44973);
  and GNAME54781(G54781,G54779,G54782);
  nand GNAME54782(G54782,G80,G54784);
  buf GNAME54783(G54783,G54779);
  buf GNAME54784(G54784,G54774);
  dff DFF_54793(CK,G54792,G44943);
  and GNAME54794(G54794,G54792,G54795);
  nand GNAME54795(G54795,G80,G54797);
  buf GNAME54796(G54796,G54792);
  buf GNAME54797(G54797,G54787);
  dff DFF_54806(CK,G54805,G50714);
  and GNAME54807(G54807,G54805,G54808);
  nand GNAME54808(G54808,G80,G54810);
  buf GNAME54809(G54809,G54805);
  buf GNAME54810(G54810,G54800);
  dff DFF_54819(CK,G54818,G54710);
  and GNAME54820(G54820,G54818,G54821);
  nand GNAME54821(G54821,G80,G54823);
  buf GNAME54822(G54822,G54818);
  buf GNAME54823(G54823,G54813);
  dff DFF_54832(CK,G54831,G54739);
  and GNAME54833(G54833,G54831,G54834);
  nand GNAME54834(G54834,G80,G54836);
  buf GNAME54835(G54835,G54831);
  buf GNAME54836(G54836,G54826);
  dff DFF_54845(CK,G54844,G47238);
  and GNAME54846(G54846,G54844,G54847);
  nand GNAME54847(G54847,G80,G54849);
  buf GNAME54848(G54848,G54844);
  buf GNAME54849(G54849,G54839);
  dff DFF_54858(CK,G54857,G48933);
  and GNAME54859(G54859,G54857,G54860);
  nand GNAME54860(G54860,G80,G54862);
  buf GNAME54861(G54861,G54857);
  buf GNAME54862(G54862,G54852);
  dff DFF_54871(CK,G54870,G47223);
  and GNAME54872(G54872,G54870,G54873);
  nand GNAME54873(G54873,G80,G54875);
  buf GNAME54874(G54874,G54870);
  buf GNAME54875(G54875,G54865);
  dff DFF_54884(CK,G54883,G48918);
  and GNAME54885(G54885,G54883,G54886);
  nand GNAME54886(G54886,G80,G54888);
  buf GNAME54887(G54887,G54883);
  buf GNAME54888(G54888,G54878);
  dff DFF_54897(CK,G54896,G49353);
  and GNAME54898(G54898,G54896,G54899);
  nand GNAME54899(G54899,G80,G54901);
  buf GNAME54900(G54900,G54896);
  buf GNAME54901(G54901,G54891);
  dff DFF_54910(CK,G54909,G49818);
  and GNAME54911(G54911,G54909,G54912);
  nand GNAME54912(G54912,G80,G54914);
  buf GNAME54913(G54913,G54909);
  buf GNAME54914(G54914,G54904);
  dff DFF_54923(CK,G54922,G49368);
  and GNAME54924(G54924,G54922,G54925);
  nand GNAME54925(G54925,G80,G54927);
  buf GNAME54926(G54926,G54922);
  buf GNAME54927(G54927,G54917);
  dff DFF_54936(CK,G54935,G50711);
  and GNAME54937(G54937,G54935,G54938);
  nand GNAME54938(G54938,G80,G54940);
  buf GNAME54939(G54939,G54935);
  buf GNAME54940(G54940,G54930);
  dff DFF_54949(CK,G54948,G48903);
  and GNAME54950(G54950,G54948,G54951);
  nand GNAME54951(G54951,G80,G54953);
  buf GNAME54952(G54952,G54948);
  buf GNAME54953(G54953,G54943);
  dff DFF_54962(CK,G54961,G48888);
  and GNAME54963(G54963,G54961,G54964);
  nand GNAME54964(G54964,G80,G54966);
  buf GNAME54965(G54965,G54961);
  buf GNAME54966(G54966,G54956);
  dff DFF_54975(CK,G54974,G48873);
  and GNAME54976(G54976,G54974,G54977);
  nand GNAME54977(G54977,G80,G54979);
  buf GNAME54978(G54978,G54974);
  buf GNAME54979(G54979,G54969);
  dff DFF_54988(CK,G54987,G48858);
  and GNAME54989(G54989,G54987,G54990);
  nand GNAME54990(G54990,G80,G54992);
  buf GNAME54991(G54991,G54987);
  buf GNAME54992(G54992,G54982);
  dff DFF_55001(CK,G55000,G49833);
  and GNAME55002(G55002,G55000,G55003);
  nand GNAME55003(G55003,G80,G55005);
  buf GNAME55004(G55004,G55000);
  buf GNAME55005(G55005,G54995);
  dff DFF_55014(CK,G55013,G49848);
  and GNAME55015(G55015,G55013,G55016);
  nand GNAME55016(G55016,G80,G55018);
  buf GNAME55017(G55017,G55013);
  buf GNAME55018(G55018,G55008);
  dff DFF_55027(CK,G55026,G49863);
  and GNAME55028(G55028,G55026,G55029);
  nand GNAME55029(G55029,G80,G55031);
  buf GNAME55030(G55030,G55026);
  buf GNAME55031(G55031,G55021);
  dff DFF_55040(CK,G55039,G49908);
  and GNAME55041(G55041,G55039,G55042);
  nand GNAME55042(G55042,G80,G55044);
  buf GNAME55043(G55043,G55039);
  buf GNAME55044(G55044,G55034);
  dff DFF_55053(CK,G55052,G50708);
  and GNAME55054(G55054,G55052,G55055);
  nand GNAME55055(G55055,G80,G55057);
  buf GNAME55056(G55056,G55052);
  buf GNAME55057(G55057,G55047);
  dff DFF_55066(CK,G55065,G50705);
  and GNAME55067(G55067,G55065,G55068);
  nand GNAME55068(G55068,G80,G55070);
  buf GNAME55069(G55069,G55065);
  buf GNAME55070(G55070,G55060);
  dff DFF_55079(CK,G55078,G48843);
  and GNAME55080(G55080,G55078,G55081);
  nand GNAME55081(G55081,G80,G55083);
  buf GNAME55082(G55082,G55078);
  buf GNAME55083(G55083,G55073);
  dff DFF_55092(CK,G55091,G48828);
  and GNAME55093(G55093,G55091,G55094);
  nand GNAME55094(G55094,G80,G55096);
  buf GNAME55095(G55095,G55091);
  buf GNAME55096(G55096,G55086);
  dff DFF_55105(CK,G55104,G48813);
  and GNAME55106(G55106,G55104,G55107);
  nand GNAME55107(G55107,G80,G55109);
  buf GNAME55108(G55108,G55104);
  buf GNAME55109(G55109,G55099);
  dff DFF_55118(CK,G55117,G48798);
  and GNAME55119(G55119,G55117,G55120);
  nand GNAME55120(G55120,G80,G55122);
  buf GNAME55121(G55121,G55117);
  buf GNAME55122(G55122,G55112);
  dff DFF_55131(CK,G55130,G49878);
  and GNAME55132(G55132,G55130,G55133);
  nand GNAME55133(G55133,G80,G55135);
  buf GNAME55134(G55134,G55130);
  buf GNAME55135(G55135,G55125);
  dff DFF_55144(CK,G55143,G49893);
  and GNAME55145(G55145,G55143,G55146);
  nand GNAME55146(G55146,G80,G55148);
  buf GNAME55147(G55147,G55143);
  buf GNAME55148(G55148,G55138);
  dff DFF_55157(CK,G55156,G49923);
  and GNAME55158(G55158,G55156,G55159);
  nand GNAME55159(G55159,G80,G55161);
  buf GNAME55160(G55160,G55156);
  buf GNAME55161(G55161,G55151);
  dff DFF_55170(CK,G55169,G49968);
  and GNAME55171(G55171,G55169,G55172);
  nand GNAME55172(G55172,G80,G55174);
  buf GNAME55173(G55173,G55169);
  buf GNAME55174(G55174,G55164);
  dff DFF_55183(CK,G55182,G50702);
  and GNAME55184(G55184,G55182,G55185);
  nand GNAME55185(G55185,G80,G55187);
  buf GNAME55186(G55186,G55182);
  buf GNAME55187(G55187,G55177);
  dff DFF_55196(CK,G55195,G50723);
  and GNAME55197(G55197,G55195,G55198);
  nand GNAME55198(G55198,G80,G55200);
  buf GNAME55199(G55199,G55195);
  buf GNAME55200(G55200,G55190);
  dff DFF_55209(CK,G55208,G48783);
  and GNAME55210(G55210,G55208,G55211);
  nand GNAME55211(G55211,G80,G55213);
  buf GNAME55212(G55212,G55208);
  buf GNAME55213(G55213,G55203);
  dff DFF_55222(CK,G55221,G48768);
  and GNAME55223(G55223,G55221,G55224);
  nand GNAME55224(G55224,G80,G55226);
  buf GNAME55225(G55225,G55221);
  buf GNAME55226(G55226,G55216);
  dff DFF_55235(CK,G55234,G48753);
  and GNAME55236(G55236,G55234,G55237);
  nand GNAME55237(G55237,G80,G55239);
  buf GNAME55238(G55238,G55234);
  buf GNAME55239(G55239,G55229);
  dff DFF_55248(CK,G55247,G48738);
  and GNAME55249(G55249,G55247,G55250);
  nand GNAME55250(G55250,G80,G55252);
  buf GNAME55251(G55251,G55247);
  buf GNAME55252(G55252,G55242);
  dff DFF_55261(CK,G55260,G49938);
  and GNAME55262(G55262,G55260,G55263);
  nand GNAME55263(G55263,G80,G55265);
  buf GNAME55264(G55264,G55260);
  buf GNAME55265(G55265,G55255);
  dff DFF_55274(CK,G55273,G49953);
  and GNAME55275(G55275,G55273,G55276);
  nand GNAME55276(G55276,G80,G55278);
  buf GNAME55277(G55277,G55273);
  buf GNAME55278(G55278,G55268);
  dff DFF_55287(CK,G55286,G49983);
  and GNAME55288(G55288,G55286,G55289);
  nand GNAME55289(G55289,G80,G55291);
  buf GNAME55290(G55290,G55286);
  buf GNAME55291(G55291,G55281);
  dff DFF_55300(CK,G55299,G50028);
  and GNAME55301(G55301,G55299,G55302);
  nand GNAME55302(G55302,G80,G55304);
  buf GNAME55303(G55303,G55299);
  buf GNAME55304(G55304,G55294);
  dff DFF_55313(CK,G55312,G50720);
  and GNAME55314(G55314,G55312,G55315);
  nand GNAME55315(G55315,G80,G55317);
  buf GNAME55316(G55316,G55312);
  buf GNAME55317(G55317,G55307);
  dff DFF_55326(CK,G55325,G50717);
  and GNAME55327(G55327,G55325,G55328);
  nand GNAME55328(G55328,G80,G55330);
  buf GNAME55329(G55329,G55325);
  buf GNAME55330(G55330,G55320);
  dff DFF_55339(CK,G55338,G48723);
  and GNAME55340(G55340,G55338,G55341);
  nand GNAME55341(G55341,G80,G55343);
  buf GNAME55342(G55342,G55338);
  buf GNAME55343(G55343,G55333);
  dff DFF_55352(CK,G55351,G49293);
  and GNAME55353(G55353,G55351,G55354);
  nand GNAME55354(G55354,G80,G55356);
  buf GNAME55355(G55355,G55351);
  buf GNAME55356(G55356,G55346);
  dff DFF_55365(CK,G55364,G48708);
  and GNAME55366(G55366,G55364,G55367);
  nand GNAME55367(G55367,G80,G55369);
  buf GNAME55368(G55368,G55364);
  buf GNAME55369(G55369,G55359);
  dff DFF_55378(CK,G55377,G49278);
  and GNAME55379(G55379,G55377,G55380);
  nand GNAME55380(G55380,G80,G55382);
  buf GNAME55381(G55381,G55377);
  buf GNAME55382(G55382,G55372);
  dff DFF_55391(CK,G55390,G49998);
  and GNAME55392(G55392,G55390,G55393);
  nand GNAME55393(G55393,G80,G55395);
  buf GNAME55394(G55394,G55390);
  buf GNAME55395(G55395,G55385);
  dff DFF_55404(CK,G55403,G50013);
  and GNAME55405(G55405,G55403,G55406);
  nand GNAME55406(G55406,G80,G55408);
  buf GNAME55407(G55407,G55403);
  buf GNAME55408(G55408,G55398);
  dff DFF_55417(CK,G55416,G50043);
  and GNAME55418(G55418,G55416,G55419);
  nand GNAME55419(G55419,G80,G55421);
  buf GNAME55420(G55420,G55416);
  buf GNAME55421(G55421,G55411);
  dff DFF_55430(CK,G55429,G50058);
  and GNAME55431(G55431,G55429,G55432);
  nand GNAME55432(G55432,G80,G55434);
  buf GNAME55433(G55433,G55429);
  buf GNAME55434(G55434,G55424);
  dff DFF_55443(CK,G55442,G50726);
  and GNAME55444(G55444,G55442,G55445);
  nand GNAME55445(G55445,G80,G55447);
  buf GNAME55446(G55446,G55442);
  buf GNAME55447(G55447,G55437);
  dff DFF_55456(CK,G55455,G50729);
  and GNAME55457(G55457,G55455,G55458);
  nand GNAME55458(G55458,G80,G55460);
  buf GNAME55459(G55459,G55455);
  buf GNAME55460(G55460,G55450);
  dff DFF_55469(CK,G55468,G49263);
  and GNAME55470(G55470,G55468,G55471);
  nand GNAME55471(G55471,G80,G55473);
  buf GNAME55472(G55472,G55468);
  buf GNAME55473(G55473,G55463);
  dff DFF_55482(CK,G55481,G49248);
  and GNAME55483(G55483,G55481,G55484);
  nand GNAME55484(G55484,G80,G55486);
  buf GNAME55485(G55485,G55481);
  buf GNAME55486(G55486,G55476);
  dff DFF_55495(CK,G55494,G49233);
  and GNAME55496(G55496,G55494,G55497);
  nand GNAME55497(G55497,G80,G55499);
  buf GNAME55498(G55498,G55494);
  buf GNAME55499(G55499,G55489);
  dff DFF_55508(CK,G55507,G49218);
  and GNAME55509(G55509,G55507,G55510);
  nand GNAME55510(G55510,G80,G55512);
  buf GNAME55511(G55511,G55507);
  buf GNAME55512(G55512,G55502);
  dff DFF_55521(CK,G55520,G50073);
  and GNAME55522(G55522,G55520,G55523);
  nand GNAME55523(G55523,G80,G55525);
  buf GNAME55524(G55524,G55520);
  buf GNAME55525(G55525,G55515);
  dff DFF_55534(CK,G55533,G50088);
  and GNAME55535(G55535,G55533,G55536);
  nand GNAME55536(G55536,G80,G55538);
  buf GNAME55537(G55537,G55533);
  buf GNAME55538(G55538,G55528);
  dff DFF_55547(CK,G55546,G50103);
  and GNAME55548(G55548,G55546,G55549);
  nand GNAME55549(G55549,G80,G55551);
  buf GNAME55550(G55550,G55546);
  buf GNAME55551(G55551,G55541);
  dff DFF_55560(CK,G55559,G50118);
  and GNAME55561(G55561,G55559,G55562);
  nand GNAME55562(G55562,G80,G55564);
  buf GNAME55563(G55563,G55559);
  buf GNAME55564(G55564,G55554);
  dff DFF_55573(CK,G55572,G50741);
  and GNAME55574(G55574,G55572,G55575);
  nand GNAME55575(G55575,G80,G55577);
  buf GNAME55576(G55576,G55572);
  buf GNAME55577(G55577,G55567);
  dff DFF_55586(CK,G55585,G50738);
  and GNAME55587(G55587,G55585,G55588);
  nand GNAME55588(G55588,G80,G55590);
  buf GNAME55589(G55589,G55585);
  buf GNAME55590(G55590,G55580);
  dff DFF_55599(CK,G55598,G49203);
  and GNAME55600(G55600,G55598,G55601);
  nand GNAME55601(G55601,G80,G55603);
  buf GNAME55602(G55602,G55598);
  buf GNAME55603(G55603,G55593);
  dff DFF_55612(CK,G55611,G49188);
  and GNAME55613(G55613,G55611,G55614);
  nand GNAME55614(G55614,G80,G55616);
  buf GNAME55615(G55615,G55611);
  buf GNAME55616(G55616,G55606);
  dff DFF_55625(CK,G55624,G49173);
  and GNAME55626(G55626,G55624,G55627);
  nand GNAME55627(G55627,G80,G55629);
  buf GNAME55628(G55628,G55624);
  buf GNAME55629(G55629,G55619);
  dff DFF_55638(CK,G55637,G49158);
  and GNAME55639(G55639,G55637,G55640);
  nand GNAME55640(G55640,G80,G55642);
  buf GNAME55641(G55641,G55637);
  buf GNAME55642(G55642,G55632);
  dff DFF_55651(CK,G55650,G50133);
  and GNAME55652(G55652,G55650,G55653);
  nand GNAME55653(G55653,G80,G55655);
  buf GNAME55654(G55654,G55650);
  buf GNAME55655(G55655,G55645);
  dff DFF_55664(CK,G55663,G50148);
  and GNAME55665(G55665,G55663,G55666);
  nand GNAME55666(G55666,G80,G55668);
  buf GNAME55667(G55667,G55663);
  buf GNAME55668(G55668,G55658);
  dff DFF_55677(CK,G55676,G50163);
  and GNAME55678(G55678,G55676,G55679);
  nand GNAME55679(G55679,G80,G55681);
  buf GNAME55680(G55680,G55676);
  buf GNAME55681(G55681,G55671);
  dff DFF_55690(CK,G55689,G50178);
  and GNAME55691(G55691,G55689,G55692);
  nand GNAME55692(G55692,G80,G55694);
  buf GNAME55693(G55693,G55689);
  buf GNAME55694(G55694,G55684);
  dff DFF_55703(CK,G55702,G50735);
  and GNAME55704(G55704,G55702,G55705);
  nand GNAME55705(G55705,G80,G55707);
  buf GNAME55706(G55706,G55702);
  buf GNAME55707(G55707,G55697);
  dff DFF_55716(CK,G55715,G50732);
  and GNAME55717(G55717,G55715,G55718);
  nand GNAME55718(G55718,G80,G55720);
  buf GNAME55719(G55719,G55715);
  buf GNAME55720(G55720,G55710);
  dff DFF_55729(CK,G55728,G49143);
  and GNAME55730(G55730,G55728,G55731);
  nand GNAME55731(G55731,G80,G55733);
  buf GNAME55732(G55732,G55728);
  buf GNAME55733(G55733,G55723);
  dff DFF_55742(CK,G55741,G49128);
  and GNAME55743(G55743,G55741,G55744);
  nand GNAME55744(G55744,G80,G55746);
  buf GNAME55745(G55745,G55741);
  buf GNAME55746(G55746,G55736);
  dff DFF_55755(CK,G55754,G49113);
  and GNAME55756(G55756,G55754,G55757);
  nand GNAME55757(G55757,G80,G55759);
  buf GNAME55758(G55758,G55754);
  buf GNAME55759(G55759,G55749);
  dff DFF_55768(CK,G55767,G49098);
  and GNAME55769(G55769,G55767,G55770);
  nand GNAME55770(G55770,G80,G55772);
  buf GNAME55771(G55771,G55767);
  buf GNAME55772(G55772,G55762);
  dff DFF_55781(CK,G55780,G50193);
  and GNAME55782(G55782,G55780,G55783);
  nand GNAME55783(G55783,G80,G55785);
  buf GNAME55784(G55784,G55780);
  buf GNAME55785(G55785,G55775);
  dff DFF_55794(CK,G55793,G50208);
  and GNAME55795(G55795,G55793,G55796);
  nand GNAME55796(G55796,G80,G55798);
  buf GNAME55797(G55797,G55793);
  buf GNAME55798(G55798,G55788);
  dff DFF_55807(CK,G55806,G50223);
  and GNAME55808(G55808,G55806,G55809);
  nand GNAME55809(G55809,G80,G55811);
  buf GNAME55810(G55810,G55806);
  buf GNAME55811(G55811,G55801);
  dff DFF_55820(CK,G55819,G50238);
  and GNAME55821(G55821,G55819,G55822);
  nand GNAME55822(G55822,G80,G55824);
  buf GNAME55823(G55823,G55819);
  buf GNAME55824(G55824,G55814);
  dff DFF_55833(CK,G55832,G50756);
  and GNAME55834(G55834,G55832,G55835);
  nand GNAME55835(G55835,G80,G55837);
  buf GNAME55836(G55836,G55832);
  buf GNAME55837(G55837,G55827);
  dff DFF_55846(CK,G55845,G50753);
  and GNAME55847(G55847,G55845,G55848);
  nand GNAME55848(G55848,G80,G55850);
  buf GNAME55849(G55849,G55845);
  buf GNAME55850(G55850,G55840);
  dff DFF_55859(CK,G55858,G49083);
  and GNAME55860(G55860,G55858,G55861);
  nand GNAME55861(G55861,G80,G55863);
  buf GNAME55862(G55862,G55858);
  buf GNAME55863(G55863,G55853);
  dff DFF_55872(CK,G55871,G48693);
  and GNAME55873(G55873,G55871,G55874);
  nand GNAME55874(G55874,G80,G55876);
  buf GNAME55875(G55875,G55871);
  buf GNAME55876(G55876,G55866);
  dff DFF_55885(CK,G55884,G49068);
  and GNAME55886(G55886,G55884,G55887);
  nand GNAME55887(G55887,G80,G55889);
  buf GNAME55888(G55888,G55884);
  buf GNAME55889(G55889,G55879);
  dff DFF_55898(CK,G55897,G48678);
  and GNAME55899(G55899,G55897,G55900);
  nand GNAME55900(G55900,G80,G55902);
  buf GNAME55901(G55901,G55897);
  buf GNAME55902(G55902,G55892);
  dff DFF_55911(CK,G55910,G50253);
  and GNAME55912(G55912,G55910,G55913);
  nand GNAME55913(G55913,G80,G55915);
  buf GNAME55914(G55914,G55910);
  buf GNAME55915(G55915,G55905);
  dff DFF_55924(CK,G55923,G50268);
  and GNAME55925(G55925,G55923,G55926);
  nand GNAME55926(G55926,G80,G55928);
  buf GNAME55927(G55927,G55923);
  buf GNAME55928(G55928,G55918);
  dff DFF_55937(CK,G55936,G50283);
  and GNAME55938(G55938,G55936,G55939);
  nand GNAME55939(G55939,G80,G55941);
  buf GNAME55940(G55940,G55936);
  buf GNAME55941(G55941,G55931);
  dff DFF_55950(CK,G55949,G50298);
  and GNAME55951(G55951,G55949,G55952);
  nand GNAME55952(G55952,G80,G55954);
  buf GNAME55953(G55953,G55949);
  buf GNAME55954(G55954,G55944);
  dff DFF_55963(CK,G55962,G50750);
  and GNAME55964(G55964,G55962,G55965);
  nand GNAME55965(G55965,G80,G55967);
  buf GNAME55966(G55966,G55962);
  buf GNAME55967(G55967,G55957);
  dff DFF_55976(CK,G55975,G50747);
  and GNAME55977(G55977,G55975,G55978);
  nand GNAME55978(G55978,G80,G55980);
  buf GNAME55979(G55979,G55975);
  buf GNAME55980(G55980,G55970);
  dff DFF_55989(CK,G55988,G47208);
  and GNAME55990(G55990,G55988,G55991);
  nand GNAME55991(G55991,G80,G55993);
  buf GNAME55992(G55992,G55988);
  buf GNAME55993(G55993,G55983);
  dff DFF_56002(CK,G56001,G48663);
  and GNAME56003(G56003,G56001,G56004);
  nand GNAME56004(G56004,G80,G56006);
  buf GNAME56005(G56005,G56001);
  buf GNAME56006(G56006,G55996);
  dff DFF_56015(CK,G56014,G48648);
  and GNAME56016(G56016,G56014,G56017);
  nand GNAME56017(G56017,G80,G56019);
  buf GNAME56018(G56018,G56014);
  buf GNAME56019(G56019,G56009);
  dff DFF_56028(CK,G56027,G47193);
  and GNAME56029(G56029,G56027,G56030);
  nand GNAME56030(G56030,G80,G56032);
  buf GNAME56031(G56031,G56027);
  buf GNAME56032(G56032,G56022);
  dff DFF_56041(CK,G56040,G48633);
  and GNAME56042(G56042,G56040,G56043);
  nand GNAME56043(G56043,G80,G56045);
  buf GNAME56044(G56044,G56040);
  buf GNAME56045(G56045,G56035);
  dff DFF_56054(CK,G56053,G48618);
  and GNAME56055(G56055,G56053,G56056);
  nand GNAME56056(G56056,G80,G56058);
  buf GNAME56057(G56057,G56053);
  buf GNAME56058(G56058,G56048);
  dff DFF_56067(CK,G56066,G48603);
  and GNAME56068(G56068,G56066,G56069);
  nand GNAME56069(G56069,G80,G56071);
  buf GNAME56070(G56070,G56066);
  buf GNAME56071(G56071,G56061);
  dff DFF_56080(CK,G56079,G48588);
  and GNAME56081(G56081,G56079,G56082);
  nand GNAME56082(G56082,G80,G56084);
  buf GNAME56083(G56083,G56079);
  buf GNAME56084(G56084,G56074);
  dff DFF_56093(CK,G56092,G48573);
  and GNAME56094(G56094,G56092,G56095);
  nand GNAME56095(G56095,G80,G56097);
  buf GNAME56096(G56096,G56092);
  buf GNAME56097(G56097,G56087);
  dff DFF_56106(CK,G56105,G50313);
  and GNAME56107(G56107,G56105,G56108);
  nand GNAME56108(G56108,G80,G56110);
  buf GNAME56109(G56109,G56105);
  buf GNAME56110(G56110,G56100);
  dff DFF_56119(CK,G56118,G50328);
  and GNAME56120(G56120,G56118,G56121);
  nand GNAME56121(G56121,G80,G56123);
  buf GNAME56122(G56122,G56118);
  buf GNAME56123(G56123,G56113);
  dff DFF_56132(CK,G56131,G50358);
  and GNAME56133(G56133,G56131,G56134);
  nand GNAME56134(G56134,G80,G56136);
  buf GNAME56135(G56135,G56131);
  buf GNAME56136(G56136,G56126);
  dff DFF_56145(CK,G56144,G50373);
  and GNAME56146(G56146,G56144,G56147);
  nand GNAME56147(G56147,G80,G56149);
  buf GNAME56148(G56148,G56144);
  buf GNAME56149(G56149,G56139);
  dff DFF_56158(CK,G56157,G50744);
  and GNAME56159(G56159,G56157,G56160);
  nand GNAME56160(G56160,G80,G56162);
  buf GNAME56161(G56161,G56157);
  buf GNAME56162(G56162,G56152);
  dff DFF_56171(CK,G56170,G50768);
  and GNAME56172(G56172,G56170,G56173);
  nand GNAME56173(G56173,G80,G56175);
  buf GNAME56174(G56174,G56170);
  buf GNAME56175(G56175,G56165);
  dff DFF_56184(CK,G56183,G48558);
  and GNAME56185(G56185,G56183,G56186);
  nand GNAME56186(G56186,G80,G56188);
  buf GNAME56187(G56187,G56183);
  buf GNAME56188(G56188,G56178);
  dff DFF_56197(CK,G56196,G48543);
  and GNAME56198(G56198,G56196,G56199);
  nand GNAME56199(G56199,G80,G56201);
  buf GNAME56200(G56200,G56196);
  buf GNAME56201(G56201,G56191);
  dff DFF_56210(CK,G56209,G48528);
  and GNAME56211(G56211,G56209,G56212);
  nand GNAME56212(G56212,G80,G56214);
  buf GNAME56213(G56213,G56209);
  buf GNAME56214(G56214,G56204);
  dff DFF_56223(CK,G56222,G48513);
  and GNAME56224(G56224,G56222,G56225);
  nand GNAME56225(G56225,G80,G56227);
  buf GNAME56226(G56226,G56222);
  buf GNAME56227(G56227,G56217);
  dff DFF_56236(CK,G56235,G48498);
  and GNAME56237(G56237,G56235,G56238);
  nand GNAME56238(G56238,G80,G56240);
  buf GNAME56239(G56239,G56235);
  buf GNAME56240(G56240,G56230);
  dff DFF_56249(CK,G56248,G48483);
  and GNAME56250(G56250,G56248,G56251);
  nand GNAME56251(G56251,G80,G56253);
  buf GNAME56252(G56252,G56248);
  buf GNAME56253(G56253,G56243);
  dff DFF_56262(CK,G56261,G48468);
  and GNAME56263(G56263,G56261,G56264);
  nand GNAME56264(G56264,G80,G56266);
  buf GNAME56265(G56265,G56261);
  buf GNAME56266(G56266,G56256);
  dff DFF_56275(CK,G56274,G48453);
  and GNAME56276(G56276,G56274,G56277);
  nand GNAME56277(G56277,G80,G56279);
  buf GNAME56278(G56278,G56274);
  buf GNAME56279(G56279,G56269);
  dff DFF_56288(CK,G56287,G50343);
  and GNAME56289(G56289,G56287,G56290);
  nand GNAME56290(G56290,G80,G56292);
  buf GNAME56291(G56291,G56287);
  buf GNAME56292(G56292,G56282);
  dff DFF_56301(CK,G56300,G50388);
  and GNAME56302(G56302,G56300,G56303);
  nand GNAME56303(G56303,G80,G56305);
  buf GNAME56304(G56304,G56300);
  buf GNAME56305(G56305,G56295);
  dff DFF_56314(CK,G56313,G50403);
  and GNAME56315(G56315,G56313,G56316);
  nand GNAME56316(G56316,G80,G56318);
  buf GNAME56317(G56317,G56313);
  buf GNAME56318(G56318,G56308);
  dff DFF_56327(CK,G56326,G50418);
  and GNAME56328(G56328,G56326,G56329);
  nand GNAME56329(G56329,G80,G56331);
  buf GNAME56330(G56330,G56326);
  buf GNAME56331(G56331,G56321);
  dff DFF_56340(CK,G56339,G50433);
  and GNAME56341(G56341,G56339,G56342);
  nand GNAME56342(G56342,G80,G56344);
  buf GNAME56343(G56343,G56339);
  buf GNAME56344(G56344,G56334);
  dff DFF_56353(CK,G56352,G50765);
  and GNAME56354(G56354,G56352,G56355);
  nand GNAME56355(G56355,G80,G56357);
  buf GNAME56356(G56356,G56352);
  buf GNAME56357(G56357,G56347);
  dff DFF_56366(CK,G56365,G50762);
  and GNAME56367(G56367,G56365,G56368);
  nand GNAME56368(G56368,G80,G56370);
  buf GNAME56369(G56369,G56365);
  buf GNAME56370(G56370,G56360);
  dff DFF_56379(CK,G56378,G48438);
  and GNAME56380(G56380,G56378,G56381);
  nand GNAME56381(G56381,G80,G56383);
  buf GNAME56382(G56382,G56378);
  buf GNAME56383(G56383,G56373);
  dff DFF_56392(CK,G56391,G48423);
  and GNAME56393(G56393,G56391,G56394);
  nand GNAME56394(G56394,G80,G56396);
  buf GNAME56395(G56395,G56391);
  buf GNAME56396(G56396,G56386);
  dff DFF_56405(CK,G56404,G48408);
  and GNAME56406(G56406,G56404,G56407);
  nand GNAME56407(G56407,G80,G56409);
  buf GNAME56408(G56408,G56404);
  buf GNAME56409(G56409,G56399);
  dff DFF_56418(CK,G56417,G49053);
  and GNAME56419(G56419,G56417,G56420);
  nand GNAME56420(G56420,G80,G56422);
  buf GNAME56421(G56421,G56417);
  buf GNAME56422(G56422,G56412);
  dff DFF_56431(CK,G56430,G49038);
  and GNAME56432(G56432,G56430,G56433);
  nand GNAME56433(G56433,G80,G56435);
  buf GNAME56434(G56434,G56430);
  buf GNAME56435(G56435,G56425);
  dff DFF_56444(CK,G56443,G49023);
  and GNAME56445(G56445,G56443,G56446);
  nand GNAME56446(G56446,G80,G56448);
  buf GNAME56447(G56447,G56443);
  buf GNAME56448(G56448,G56438);
  dff DFF_56457(CK,G56456,G49008);
  and GNAME56458(G56458,G56456,G56459);
  nand GNAME56459(G56459,G80,G56461);
  buf GNAME56460(G56460,G56456);
  buf GNAME56461(G56461,G56451);
  dff DFF_56470(CK,G56469,G48393);
  and GNAME56471(G56471,G56469,G56472);
  nand GNAME56472(G56472,G80,G56474);
  buf GNAME56473(G56473,G56469);
  buf GNAME56474(G56474,G56464);
  dff DFF_56483(CK,G56482,G48378);
  and GNAME56484(G56484,G56482,G56485);
  nand GNAME56485(G56485,G80,G56487);
  buf GNAME56486(G56486,G56482);
  buf GNAME56487(G56487,G56477);
  dff DFF_56496(CK,G56495,G50448);
  and GNAME56497(G56497,G56495,G56498);
  nand GNAME56498(G56498,G80,G56500);
  buf GNAME56499(G56499,G56495);
  buf GNAME56500(G56500,G56490);
  dff DFF_56509(CK,G56508,G50463);
  and GNAME56510(G56510,G56508,G56511);
  nand GNAME56511(G56511,G80,G56513);
  buf GNAME56512(G56512,G56508);
  buf GNAME56513(G56513,G56503);
  dff DFF_56522(CK,G56521,G50478);
  and GNAME56523(G56523,G56521,G56524);
  nand GNAME56524(G56524,G80,G56526);
  buf GNAME56525(G56525,G56521);
  buf GNAME56526(G56526,G56516);
  dff DFF_56535(CK,G56534,G50493);
  and GNAME56536(G56536,G56534,G56537);
  nand GNAME56537(G56537,G80,G56539);
  buf GNAME56538(G56538,G56534);
  buf GNAME56539(G56539,G56529);
  dff DFF_56548(CK,G56547,G50759);
  and GNAME56549(G56549,G56547,G56550);
  nand GNAME56550(G56550,G80,G56552);
  buf GNAME56551(G56551,G56547);
  buf GNAME56552(G56552,G56542);
  dff DFF_56561(CK,G56560,G50783);
  and GNAME56562(G56562,G56560,G56563);
  nand GNAME56563(G56563,G80,G56565);
  buf GNAME56564(G56564,G56560);
  buf GNAME56565(G56565,G56555);
  dff DFF_56574(CK,G56573,G48363);
  and GNAME56575(G56575,G56573,G56576);
  nand GNAME56576(G56576,G80,G56578);
  buf GNAME56577(G56577,G56573);
  buf GNAME56578(G56578,G56568);
  dff DFF_56587(CK,G56586,G48348);
  and GNAME56588(G56588,G56586,G56589);
  nand GNAME56589(G56589,G80,G56591);
  buf GNAME56590(G56590,G56586);
  buf GNAME56591(G56591,G56581);
  dff DFF_56600(CK,G56599,G48993);
  and GNAME56601(G56601,G56599,G56602);
  nand GNAME56602(G56602,G80,G56604);
  buf GNAME56603(G56603,G56599);
  buf GNAME56604(G56604,G56594);
  dff DFF_56613(CK,G56612,G48978);
  and GNAME56614(G56614,G56612,G56615);
  nand GNAME56615(G56615,G80,G56617);
  buf GNAME56616(G56616,G56612);
  buf GNAME56617(G56617,G56607);
  dff DFF_56626(CK,G56625,G48963);
  and GNAME56627(G56627,G56625,G56628);
  nand GNAME56628(G56628,G80,G56630);
  buf GNAME56629(G56629,G56625);
  buf GNAME56630(G56630,G56620);
  dff DFF_56639(CK,G56638,G48948);
  and GNAME56640(G56640,G56638,G56641);
  nand GNAME56641(G56641,G80,G56643);
  buf GNAME56642(G56642,G56638);
  buf GNAME56643(G56643,G56633);
  dff DFF_56652(CK,G56651,G48333);
  and GNAME56653(G56653,G56651,G56654);
  nand GNAME56654(G56654,G80,G56656);
  buf GNAME56655(G56655,G56651);
  buf GNAME56656(G56656,G56646);
  dff DFF_56665(CK,G56664,G48318);
  and GNAME56666(G56666,G56664,G56667);
  nand GNAME56667(G56667,G80,G56669);
  buf GNAME56668(G56668,G56664);
  buf GNAME56669(G56669,G56659);
  dff DFF_56678(CK,G56677,G50508);
  and GNAME56679(G56679,G56677,G56680);
  nand GNAME56680(G56680,G80,G56682);
  buf GNAME56681(G56681,G56677);
  buf GNAME56682(G56682,G56672);
  dff DFF_56691(CK,G56690,G50523);
  and GNAME56692(G56692,G56690,G56693);
  nand GNAME56693(G56693,G80,G56695);
  buf GNAME56694(G56694,G56690);
  buf GNAME56695(G56695,G56685);
  dff DFF_56704(CK,G56703,G50538);
  and GNAME56705(G56705,G56703,G56706);
  nand GNAME56706(G56706,G80,G56708);
  buf GNAME56707(G56707,G56703);
  buf GNAME56708(G56708,G56698);
  dff DFF_56717(CK,G56716,G50553);
  and GNAME56718(G56718,G56716,G56719);
  nand GNAME56719(G56719,G80,G56721);
  buf GNAME56720(G56720,G56716);
  buf GNAME56721(G56721,G56711);
  dff DFF_56730(CK,G56729,G50780);
  and GNAME56731(G56731,G56729,G56732);
  nand GNAME56732(G56732,G80,G56734);
  buf GNAME56733(G56733,G56729);
  buf GNAME56734(G56734,G56724);
  dff DFF_56743(CK,G56742,G50777);
  and GNAME56744(G56744,G56742,G56745);
  nand GNAME56745(G56745,G80,G56747);
  buf GNAME56746(G56746,G56742);
  buf GNAME56747(G56747,G56737);
  dff DFF_56756(CK,G56755,G47178);
  and GNAME56757(G56757,G56755,G56758);
  nand GNAME56758(G56758,G80,G56760);
  buf GNAME56759(G56759,G56755);
  buf GNAME56760(G56760,G56750);
  dff DFF_56769(CK,G56768,G47163);
  and GNAME56770(G56770,G56768,G56771);
  nand GNAME56771(G56771,G80,G56773);
  buf GNAME56772(G56772,G56768);
  buf GNAME56773(G56773,G56763);
  dff DFF_56782(CK,G56781,G48303);
  and GNAME56783(G56783,G56781,G56784);
  nand GNAME56784(G56784,G80,G56786);
  buf GNAME56785(G56785,G56781);
  buf GNAME56786(G56786,G56776);
  dff DFF_56795(CK,G56794,G48288);
  and GNAME56796(G56796,G56794,G56797);
  nand GNAME56797(G56797,G80,G56799);
  buf GNAME56798(G56798,G56794);
  buf GNAME56799(G56799,G56789);
  dff DFF_56808(CK,G56807,G48273);
  and GNAME56809(G56809,G56807,G56810);
  nand GNAME56810(G56810,G80,G56812);
  buf GNAME56811(G56811,G56807);
  buf GNAME56812(G56812,G56802);
  dff DFF_56821(CK,G56820,G48258);
  and GNAME56822(G56822,G56820,G56823);
  nand GNAME56823(G56823,G80,G56825);
  buf GNAME56824(G56824,G56820);
  buf GNAME56825(G56825,G56815);
  dff DFF_56834(CK,G56833,G48243);
  and GNAME56835(G56835,G56833,G56836);
  nand GNAME56836(G56836,G80,G56838);
  buf GNAME56837(G56837,G56833);
  buf GNAME56838(G56838,G56828);
  dff DFF_56847(CK,G56846,G47148);
  and GNAME56848(G56848,G56846,G56849);
  nand GNAME56849(G56849,G80,G56851);
  buf GNAME56850(G56850,G56846);
  buf GNAME56851(G56851,G56841);
  dff DFF_56860(CK,G56859,G47133);
  and GNAME56861(G56861,G56859,G56862);
  nand GNAME56862(G56862,G80,G56864);
  buf GNAME56863(G56863,G56859);
  buf GNAME56864(G56864,G56854);
  dff DFF_56873(CK,G56872,G50568);
  and GNAME56874(G56874,G56872,G56875);
  nand GNAME56875(G56875,G80,G56877);
  buf GNAME56876(G56876,G56872);
  buf GNAME56877(G56877,G56867);
  dff DFF_56886(CK,G56885,G50583);
  and GNAME56887(G56887,G56885,G56888);
  nand GNAME56888(G56888,G80,G56890);
  buf GNAME56889(G56889,G56885);
  buf GNAME56890(G56890,G56880);
  dff DFF_56899(CK,G56898,G50598);
  and GNAME56900(G56900,G56898,G56901);
  nand GNAME56901(G56901,G80,G56903);
  buf GNAME56902(G56902,G56898);
  buf GNAME56903(G56903,G56893);
  dff DFF_56912(CK,G56911,G50613);
  and GNAME56913(G56913,G56911,G56914);
  nand GNAME56914(G56914,G80,G56916);
  buf GNAME56915(G56915,G56911);
  buf GNAME56916(G56916,G56906);
  dff DFF_56925(CK,G56924,G50774);
  and GNAME56926(G56926,G56924,G56927);
  nand GNAME56927(G56927,G80,G56929);
  buf GNAME56928(G56928,G56924);
  buf GNAME56929(G56929,G56919);
  dff DFF_56938(CK,G56937,G50771);
  and GNAME56939(G56939,G56937,G56940);
  nand GNAME56940(G56940,G80,G56942);
  buf GNAME56941(G56941,G56937);
  buf GNAME56942(G56942,G56932);
  dff DFF_56951(CK,G56950,G47118);
  and GNAME56952(G56952,G56950,G56953);
  nand GNAME56953(G56953,G80,G56955);
  buf GNAME56954(G56954,G56950);
  buf GNAME56955(G56955,G56945);
  dff DFF_56964(CK,G56963,G47313);
  and GNAME56965(G56965,G56963,G56966);
  nand GNAME56966(G56966,G80,G56968);
  buf GNAME56967(G56967,G56963);
  buf GNAME56968(G56968,G56958);
  dff DFF_56977(CK,G56976,G48228);
  and GNAME56978(G56978,G56976,G56979);
  nand GNAME56979(G56979,G80,G56981);
  buf GNAME56980(G56980,G56976);
  buf GNAME56981(G56981,G56971);
  dff DFF_56990(CK,G56989,G48213);
  and GNAME56991(G56991,G56989,G56992);
  nand GNAME56992(G56992,G80,G56994);
  buf GNAME56993(G56993,G56989);
  buf GNAME56994(G56994,G56984);
  dff DFF_57003(CK,G57002,G48198);
  and GNAME57004(G57004,G57002,G57005);
  nand GNAME57005(G57005,G80,G57007);
  buf GNAME57006(G57006,G57002);
  buf GNAME57007(G57007,G56997);
  dff DFF_57016(CK,G57015,G48183);
  and GNAME57017(G57017,G57015,G57018);
  nand GNAME57018(G57018,G80,G57020);
  buf GNAME57019(G57019,G57015);
  buf GNAME57020(G57020,G57010);
  dff DFF_57029(CK,G57028,G47103);
  and GNAME57030(G57030,G57028,G57031);
  nand GNAME57031(G57031,G80,G57033);
  buf GNAME57032(G57032,G57028);
  buf GNAME57033(G57033,G57023);
  dff DFF_57042(CK,G57041,G47298);
  and GNAME57043(G57043,G57041,G57044);
  nand GNAME57044(G57044,G80,G57046);
  buf GNAME57045(G57045,G57041);
  buf GNAME57046(G57046,G57036);
  dff DFF_57055(CK,G57054,G50628);
  and GNAME57056(G57056,G57054,G57057);
  nand GNAME57057(G57057,G80,G57059);
  buf GNAME57058(G57058,G57054);
  buf GNAME57059(G57059,G57049);
  dff DFF_57068(CK,G57067,G49323);
  and GNAME57069(G57069,G57067,G57070);
  nand GNAME57070(G57070,G80,G57072);
  buf GNAME57071(G57071,G57067);
  buf GNAME57072(G57072,G57062);
  dff DFF_57081(CK,G57080,G50643);
  and GNAME57082(G57082,G57080,G57083);
  nand GNAME57083(G57083,G80,G57085);
  buf GNAME57084(G57084,G57080);
  buf GNAME57085(G57085,G57075);
  dff DFF_57094(CK,G57093,G50658);
  and GNAME57095(G57095,G57093,G57096);
  nand GNAME57096(G57096,G80,G57098);
  buf GNAME57097(G57097,G57093);
  buf GNAME57098(G57098,G57088);
  dff DFF_57107(CK,G57106,G50795);
  and GNAME57108(G57108,G57106,G57109);
  nand GNAME57109(G57109,G80,G57111);
  buf GNAME57110(G57110,G57106);
  buf GNAME57111(G57111,G57101);
  dff DFF_57120(CK,G57119,G50792);
  and GNAME57121(G57121,G57119,G57122);
  nand GNAME57122(G57122,G80,G57124);
  buf GNAME57123(G57123,G57119);
  buf GNAME57124(G57124,G57114);
  dff DFF_57133(CK,G57132,G44913);
  and GNAME57134(G57134,G57132,G57135);
  nand GNAME57135(G57135,G80,G57137);
  buf GNAME57136(G57136,G57132);
  buf GNAME57137(G57137,G57127);
  dff DFF_57146(CK,G57145,G52047);
  and GNAME57147(G57147,G57145,G57148);
  nand GNAME57148(G57148,G80,G57150);
  buf GNAME57149(G57149,G57145);
  buf GNAME57150(G57150,G57140);
  dff DFF_57159(CK,G57158,G51149);
  and GNAME57160(G57160,G57158,G57161);
  nand GNAME57161(G57161,G80,G57163);
  buf GNAME57162(G57162,G57158);
  buf GNAME57163(G57163,G57153);
  dff DFF_57172(CK,G57171,G51146);
  and GNAME57173(G57173,G57171,G57174);
  nand GNAME57174(G57174,G80,G57176);
  buf GNAME57175(G57175,G57171);
  buf GNAME57176(G57176,G57166);
  dff DFF_57185(CK,G57184,G51143);
  and GNAME57186(G57186,G57184,G57187);
  nand GNAME57187(G57187,G80,G57189);
  buf GNAME57188(G57188,G57184);
  buf GNAME57189(G57189,G57179);
  dff DFF_57198(CK,G57197,G51140);
  and GNAME57199(G57199,G57197,G57200);
  nand GNAME57200(G57200,G80,G57202);
  buf GNAME57201(G57201,G57197);
  buf GNAME57202(G57202,G57192);
  dff DFF_57211(CK,G57210,G51137);
  and GNAME57212(G57212,G57210,G57213);
  nand GNAME57213(G57213,G80,G57215);
  buf GNAME57214(G57214,G57210);
  buf GNAME57215(G57215,G57205);
  dff DFF_57224(CK,G57223,G51134);
  and GNAME57225(G57225,G57223,G57226);
  nand GNAME57226(G57226,G80,G57228);
  buf GNAME57227(G57227,G57223);
  buf GNAME57228(G57228,G57218);
  dff DFF_57237(CK,G57236,G51131);
  and GNAME57238(G57238,G57236,G57239);
  nand GNAME57239(G57239,G80,G57241);
  buf GNAME57240(G57240,G57236);
  buf GNAME57241(G57241,G57231);
  dff DFF_57250(CK,G57249,G51128);
  and GNAME57251(G57251,G57249,G57252);
  nand GNAME57252(G57252,G80,G57254);
  buf GNAME57253(G57253,G57249);
  buf GNAME57254(G57254,G57244);
  dff DFF_57263(CK,G57262,G51125);
  and GNAME57264(G57264,G57262,G57265);
  nand GNAME57265(G57265,G80,G57267);
  buf GNAME57266(G57266,G57262);
  buf GNAME57267(G57267,G57257);
  dff DFF_57276(CK,G57275,G51122);
  and GNAME57277(G57277,G57275,G57278);
  nand GNAME57278(G57278,G80,G57280);
  buf GNAME57279(G57279,G57275);
  buf GNAME57280(G57280,G57270);
  dff DFF_57289(CK,G57288,G51119);
  and GNAME57290(G57290,G57288,G57291);
  nand GNAME57291(G57291,G80,G57293);
  buf GNAME57292(G57292,G57288);
  buf GNAME57293(G57293,G57283);
  dff DFF_57302(CK,G57301,G51116);
  and GNAME57303(G57303,G57301,G57304);
  nand GNAME57304(G57304,G80,G57306);
  buf GNAME57305(G57305,G57301);
  buf GNAME57306(G57306,G57296);
  dff DFF_57315(CK,G57314,G51113);
  and GNAME57316(G57316,G57314,G57317);
  nand GNAME57317(G57317,G80,G57319);
  buf GNAME57318(G57318,G57314);
  buf GNAME57319(G57319,G57309);
  dff DFF_57328(CK,G57327,G51110);
  and GNAME57329(G57329,G57327,G57330);
  nand GNAME57330(G57330,G80,G57332);
  buf GNAME57331(G57331,G57327);
  buf GNAME57332(G57332,G57322);
  dff DFF_57341(CK,G57340,G57852);
  and GNAME57342(G57342,G57340,G57343);
  nand GNAME57343(G57343,G80,G57345);
  buf GNAME57344(G57344,G57340);
  buf GNAME57345(G57345,G57335);
  dff DFF_57354(CK,G57353,G51107);
  and GNAME57355(G57355,G57353,G57356);
  nand GNAME57356(G57356,G80,G57358);
  buf GNAME57357(G57357,G57353);
  buf GNAME57358(G57358,G57348);
  dff DFF_57367(CK,G57366,G51104);
  and GNAME57368(G57368,G57366,G57369);
  nand GNAME57369(G57369,G80,G57371);
  buf GNAME57370(G57370,G57366);
  buf GNAME57371(G57371,G57361);
  dff DFF_57380(CK,G57379,G51101);
  and GNAME57381(G57381,G57379,G57382);
  nand GNAME57382(G57382,G80,G57384);
  buf GNAME57383(G57383,G57379);
  buf GNAME57384(G57384,G57374);
  dff DFF_57393(CK,G57392,G51098);
  and GNAME57394(G57394,G57392,G57395);
  nand GNAME57395(G57395,G80,G57397);
  buf GNAME57396(G57396,G57392);
  buf GNAME57397(G57397,G57387);
  dff DFF_57406(CK,G57405,G51095);
  and GNAME57407(G57407,G57405,G57408);
  nand GNAME57408(G57408,G80,G57410);
  buf GNAME57409(G57409,G57405);
  buf GNAME57410(G57410,G57400);
  dff DFF_57419(CK,G57418,G51092);
  and GNAME57420(G57420,G57418,G57421);
  nand GNAME57421(G57421,G80,G57423);
  buf GNAME57422(G57422,G57418);
  buf GNAME57423(G57423,G57413);
  dff DFF_57432(CK,G57431,G51089);
  and GNAME57433(G57433,G57431,G57434);
  nand GNAME57434(G57434,G80,G57436);
  buf GNAME57435(G57435,G57431);
  buf GNAME57436(G57436,G57426);
  dff DFF_57445(CK,G57444,G51086);
  and GNAME57446(G57446,G57444,G57447);
  nand GNAME57447(G57447,G80,G57449);
  buf GNAME57448(G57448,G57444);
  buf GNAME57449(G57449,G57439);
  dff DFF_57458(CK,G57457,G51173);
  and GNAME57459(G57459,G57457,G57460);
  nand GNAME57460(G57460,G80,G57462);
  buf GNAME57461(G57461,G57457);
  buf GNAME57462(G57462,G57452);
  dff DFF_57471(CK,G57470,G51170);
  and GNAME57472(G57472,G57470,G57473);
  nand GNAME57473(G57473,G80,G57475);
  buf GNAME57474(G57474,G57470);
  buf GNAME57475(G57475,G57465);
  dff DFF_57484(CK,G57483,G51167);
  and GNAME57485(G57485,G57483,G57486);
  nand GNAME57486(G57486,G80,G57488);
  buf GNAME57487(G57487,G57483);
  buf GNAME57488(G57488,G57478);
  dff DFF_57497(CK,G57496,G51164);
  and GNAME57498(G57498,G57496,G57499);
  nand GNAME57499(G57499,G80,G57501);
  buf GNAME57500(G57500,G57496);
  buf GNAME57501(G57501,G57491);
  dff DFF_57510(CK,G57509,G51161);
  and GNAME57511(G57511,G57509,G57512);
  nand GNAME57512(G57512,G80,G57514);
  buf GNAME57513(G57513,G57509);
  buf GNAME57514(G57514,G57504);
  dff DFF_57523(CK,G57522,G51158);
  and GNAME57524(G57524,G57522,G57525);
  nand GNAME57525(G57525,G80,G57527);
  buf GNAME57526(G57526,G57522);
  buf GNAME57527(G57527,G57517);
  dff DFF_57536(CK,G57535,G51155);
  and GNAME57537(G57537,G57535,G57538);
  nand GNAME57538(G57538,G80,G57540);
  buf GNAME57539(G57539,G57535);
  buf GNAME57540(G57540,G57530);
  dff DFF_57549(CK,G57548,G51152);
  and GNAME57550(G57550,G57548,G57551);
  nand GNAME57551(G57551,G80,G57553);
  buf GNAME57552(G57552,G57548);
  buf GNAME57553(G57553,G57543);
  dff DFF_57562(CK,G57561,G54745);
  and GNAME57563(G57563,G57561,G57564);
  nand GNAME57564(G57564,G80,G57566);
  buf GNAME57565(G57565,G57561);
  buf GNAME57566(G57566,G57556);
  dff DFF_57575(CK,G57574,G54743);
  and GNAME57576(G57576,G57574,G57577);
  nand GNAME57577(G57577,G80,G57579);
  buf GNAME57578(G57578,G57574);
  buf GNAME57579(G57579,G57569);
  dff DFF_57588(CK,G57587,G54741);
  and GNAME57589(G57589,G57587,G57590);
  nand GNAME57590(G57590,G80,G57592);
  buf GNAME57591(G57591,G57587);
  buf GNAME57592(G57592,G57582);
  dff DFF_57601(CK,G57600,G47088);
  and GNAME57602(G57602,G57600,G57603);
  nand GNAME57603(G57603,G80,G57605);
  buf GNAME57604(G57604,G57600);
  buf GNAME57605(G57605,G57595);
  dff DFF_57614(CK,G57613,G47073);
  and GNAME57615(G57615,G57613,G57616);
  nand GNAME57616(G57616,G80,G57618);
  buf GNAME57617(G57617,G57613);
  buf GNAME57618(G57618,G57608);
  dff DFF_57627(CK,G57626,G47058);
  and GNAME57628(G57628,G57626,G57629);
  nand GNAME57629(G57629,G80,G57631);
  buf GNAME57630(G57630,G57626);
  buf GNAME57631(G57631,G57621);
  dff DFF_57640(CK,G57639,G47283);
  and GNAME57641(G57641,G57639,G57642);
  nand GNAME57642(G57642,G80,G57644);
  buf GNAME57643(G57643,G57639);
  buf GNAME57644(G57644,G57634);
  dff DFF_57653(CK,G57652,G50673);
  and GNAME57654(G57654,G57652,G57655);
  nand GNAME57655(G57655,G80,G57657);
  buf GNAME57656(G57656,G57652);
  buf GNAME57657(G57657,G57647);
  dff DFF_57666(CK,G57665,G50688);
  and GNAME57667(G57667,G57665,G57668);
  nand GNAME57668(G57668,G80,G57670);
  buf GNAME57669(G57669,G57665);
  buf GNAME57670(G57670,G57660);
  dff DFF_57679(CK,G57678,G50789);
  and GNAME57680(G57680,G57678,G57681);
  nand GNAME57681(G57681,G80,G57683);
  buf GNAME57682(G57682,G57678);
  buf GNAME57683(G57683,G57673);
  dff DFF_57692(CK,G57691,G50786);
  and GNAME57693(G57693,G57691,G57694);
  nand GNAME57694(G57694,G80,G57696);
  buf GNAME57695(G57695,G57691);
  buf GNAME57696(G57696,G57686);
  dff DFF_57705(CK,G57704,G54714);
  and GNAME57706(G57706,G57704,G57707);
  nand GNAME57707(G57707,G80,G57709);
  buf GNAME57708(G57708,G57704);
  buf GNAME57709(G57709,G57699);
  dff DFF_57718(CK,G57717,G50693);
  and GNAME57719(G57719,G57717,G57720);
  nand GNAME57720(G57720,G80,G57722);
  buf GNAME57721(G57721,G57717);
  buf GNAME57722(G57722,G57712);
  buf GNAME57723(G57723,G57134);
  buf GNAME57724(G57724,G57134);
  buf GNAME57725(G57725,G2699);
  buf GNAME57726(G57726,G2283);
  buf GNAME57727(G57727,G1867);
  buf GNAME57728(G57728,G10250);
  buf GNAME57729(G57729,G8378);
  buf GNAME57730(G57730,G6506);
  buf GNAME57731(G57731,G2657);
  buf GNAME57732(G57732,G2241);
  buf GNAME57733(G57733,G1825);
  buf GNAME57734(G57734,G10208);
  buf GNAME57735(G57735,G8336);
  buf GNAME57736(G57736,G6464);
  buf GNAME57737(G57737,G10229);
  buf GNAME57738(G57738,G8357);
  buf GNAME57739(G57739,G6485);
  buf GNAME57740(G57740,G2615);
  buf GNAME57741(G57741,G2199);
  buf GNAME57742(G57742,G1783);
  buf GNAME57743(G57743,G10166);
  buf GNAME57744(G57744,G8294);
  buf GNAME57745(G57745,G6422);
  buf GNAME57746(G57746,G10187);
  buf GNAME57747(G57747,G8315);
  buf GNAME57748(G57748,G6443);
  buf GNAME57749(G57749,G2573);
  buf GNAME57750(G57750,G2157);
  buf GNAME57751(G57751,G1741);
  buf GNAME57752(G57752,G10124);
  buf GNAME57753(G57753,G8252);
  buf GNAME57754(G57754,G6380);
  buf GNAME57755(G57755,G10145);
  buf GNAME57756(G57756,G8273);
  buf GNAME57757(G57757,G6401);
  buf GNAME57758(G57758,G2491);
  buf GNAME57759(G57759,G2075);
  buf GNAME57760(G57760,G1659);
  buf GNAME57761(G57761,G10042);
  buf GNAME57762(G57762,G8170);
  buf GNAME57763(G57763,G6298);
  buf GNAME57764(G57764,G10103);
  buf GNAME57765(G57765,G8231);
  buf GNAME57766(G57766,G6359);
  buf GNAME57767(G57767,G2449);
  buf GNAME57768(G57768,G2033);
  buf GNAME57769(G57769,G1617);
  buf GNAME57770(G57770,G10000);
  buf GNAME57771(G57771,G10021);
  buf GNAME57772(G57772,G8128);
  buf GNAME57773(G57773,G8149);
  buf GNAME57774(G57774,G6256);
  buf GNAME57775(G57775,G6277);
  buf GNAME57776(G57776,G2407);
  buf GNAME57777(G57777,G1991);
  buf GNAME57778(G57778,G1575);
  buf GNAME57779(G57779,G54794);
  buf GNAME57780(G57780,G54781);
  buf GNAME57781(G57781,G2699);
  buf GNAME57782(G57782,G2283);
  buf GNAME57783(G57783,G1867);
  buf GNAME57784(G57784,G2657);
  buf GNAME57785(G57785,G2241);
  buf GNAME57786(G57786,G1825);
  buf GNAME57787(G57787,G54794);
  buf GNAME57788(G57788,G54781);
  buf GNAME57789(G57789,G9979);
  buf GNAME57790(G57790,G9958);
  buf GNAME57791(G57791,G9937);
  buf GNAME57792(G57792,G8107);
  buf GNAME57793(G57793,G8086);
  buf GNAME57794(G57794,G6235);
  buf GNAME57795(G57795,G6214);
  buf GNAME57796(G57796,G8065);
  buf GNAME57797(G57797,G6193);
  buf GNAME57798(G57798,G2365);
  buf GNAME57799(G57799,G1949);
  buf GNAME57800(G57800,G1533);
  buf GNAME57801(G57801,G2615);
  buf GNAME57802(G57802,G2199);
  buf GNAME57803(G57803,G1783);
  buf GNAME57804(G57804,G9687);
  buf GNAME57805(G57805,G7815);
  buf GNAME57806(G57806,G5943);
  buf GNAME57807(G57807,G9834);
  buf GNAME57808(G57808,G9895);
  buf GNAME57809(G57809,G7962);
  buf GNAME57810(G57810,G8023);
  buf GNAME57811(G57811,G6090);
  buf GNAME57812(G57812,G6151);
  buf GNAME57813(G57813,G9916);
  buf GNAME57814(G57814,G8044);
  buf GNAME57815(G57815,G6172);
  buf GNAME57816(G57816,G2573);
  buf GNAME57817(G57817,G2157);
  buf GNAME57818(G57818,G1741);
  buf GNAME57819(G57819,G9792);
  buf GNAME57820(G57820,G9771);
  buf GNAME57821(G57821,G9750);
  buf GNAME57822(G57822,G9813);
  buf GNAME57823(G57823,G7941);
  buf GNAME57824(G57824,G6069);
  buf GNAME57825(G57825,G7878);
  buf GNAME57826(G57826,G7899);
  buf GNAME57827(G57827,G7920);
  buf GNAME57828(G57828,G6006);
  buf GNAME57829(G57829,G6027);
  buf GNAME57830(G57830,G6048);
  buf GNAME57831(G57831,G2491);
  buf GNAME57832(G57832,G2075);
  buf GNAME57833(G57833,G1659);
  buf GNAME57834(G57834,G2449);
  buf GNAME57835(G57835,G2033);
  buf GNAME57836(G57836,G1617);
  buf GNAME57837(G57837,G9687);
  buf GNAME57838(G57838,G7815);
  buf GNAME57839(G57839,G5943);
  buf GNAME57840(G57840,G9729);
  buf GNAME57841(G57841,G9708);
  buf GNAME57842(G57842,G7857);
  buf GNAME57843(G57843,G7836);
  buf GNAME57844(G57844,G5985);
  buf GNAME57845(G57845,G5964);
  buf GNAME57846(G57846,G2407);
  buf GNAME57847(G57847,G1991);
  buf GNAME57848(G57848,G1575);
  buf GNAME57849(G57849,G2365);
  buf GNAME57850(G57850,G1949);
  buf GNAME57851(G57851,G1533);
  buf GNAME57852(G57852,G51230);
  buf GNAME57853(G57853,G54686);
  buf GNAME57854(G57854,G54687);
  buf GNAME57855(G57855,G54688);
  buf GNAME57856(G57856,G51230);
  buf GNAME57857(G57857,G51230);
  buf GNAME57858(G57858,G52118);
  buf GNAME57859(G57859,G52119);
  buf GNAME57860(G57860,G52120);
  buf GNAME57861(G57861,G54689);
  buf GNAME57862(G57862,G54690);
  buf GNAME57863(G57863,G54691);
  buf GNAME57864(G57864,G52121);
  buf GNAME57865(G57865,G52122);
  buf GNAME57866(G57866,G52123);
  buf GNAME57867(G57867,G54695);
  buf GNAME57868(G57868,G54692);
  buf GNAME57869(G57869,G54696);
  buf GNAME57870(G57870,G54697);
  buf GNAME57871(G57871,G54693);
  buf GNAME57872(G57872,G54694);
  buf GNAME57873(G57873,G52127);
  buf GNAME57874(G57874,G52128);
  buf GNAME57875(G57875,G52129);
  buf GNAME57876(G57876,G52127);
  buf GNAME57877(G57877,G52124);
  buf GNAME57878(G57878,G52128);
  buf GNAME57879(G57879,G52129);
  buf GNAME57880(G57880,G52125);
  buf GNAME57881(G57881,G52126);
  buf GNAME57882(G57882,G54566);
  buf GNAME57883(G57883,G54567);
  buf GNAME57884(G57884,G54568);
  buf GNAME57885(G57885,G54704);
  buf GNAME57886(G57886,G54705);
  buf GNAME57887(G57887,G54706);
  buf GNAME57888(G57888,G54707);
  buf GNAME57889(G57889,G54708);
  buf GNAME57890(G57890,G54709);
  buf GNAME57891(G57891,G54566);
  buf GNAME57892(G57892,G54567);
  buf GNAME57893(G57893,G54568);
  buf GNAME57894(G57894,G54704);
  buf GNAME57895(G57895,G54705);
  buf GNAME57896(G57896,G54706);
  buf GNAME57897(G57897,G54707);
  buf GNAME57898(G57898,G54708);
  buf GNAME57899(G57899,G54709);
  buf GNAME57900(G57900,G52133);
  buf GNAME57901(G57901,G52136);
  buf GNAME57902(G57902,G52134);
  buf GNAME57903(G57903,G52137);
  buf GNAME57904(G57904,G52135);
  buf GNAME57905(G57905,G52138);
  buf GNAME57906(G57906,G52136);
  buf GNAME57907(G57907,G52137);
  buf GNAME57908(G57908,G52138);
  buf GNAME57909(G57909,G54639);
  buf GNAME57910(G57910,G54640);
  buf GNAME57911(G57911,G54641);
  buf GNAME57912(G57912,G54640);
  buf GNAME57913(G57913,G54639);
  buf GNAME57914(G57914,G54641);
  buf GNAME57915(G57915,G54686);
  buf GNAME57916(G57916,G54689);
  buf GNAME57917(G57917,G54687);
  buf GNAME57918(G57918,G54688);
  buf GNAME57919(G57919,G54690);
  buf GNAME57920(G57920,G54691);
  buf GNAME57921(G57921,G52118);
  buf GNAME57922(G57922,G52119);
  buf GNAME57923(G57923,G52120);
  buf GNAME57924(G57924,G54695);
  buf GNAME57925(G57925,G54696);
  buf GNAME57926(G57926,G54697);
  buf GNAME57927(G57927,G52121);
  buf GNAME57928(G57928,G52122);
  buf GNAME57929(G57929,G52123);
  buf GNAME57930(G57930,G54699);
  buf GNAME57931(G57931,G54700);
  buf GNAME57932(G57932,G54701);
  buf GNAME57933(G57933,G54698);
  buf GNAME57934(G57934,G54702);
  buf GNAME57935(G57935,G54703);
  buf GNAME57936(G57936,G52124);
  buf GNAME57937(G57937,G52125);
  buf GNAME57938(G57938,G52126);
  buf GNAME57939(G57939,G52130);
  buf GNAME57940(G57940,G52131);
  buf GNAME57941(G57941,G52132);
  buf GNAME57942(G57942,G54692);
  buf GNAME57943(G57943,G54693);
  buf GNAME57944(G57944,G54694);
  buf GNAME57945(G57945,G54698);
  buf GNAME57946(G57946,G54702);
  buf GNAME57947(G57947,G54703);
  buf GNAME57948(G57948,G54699);
  buf GNAME57949(G57949,G54700);
  buf GNAME57950(G57950,G54701);
  buf GNAME57951(G57951,G52133);
  buf GNAME57952(G57952,G52134);
  buf GNAME57953(G57953,G52135);
  buf GNAME57954(G57954,G52130);
  buf GNAME57955(G57955,G52131);
  buf GNAME57956(G57956,G52132);
  xor GNAME63480(G63480,G63481,G75892);
  xor GNAME63481(G63481,G75181,G75178);
  and GNAME63482(G63482,G75181,G75892);
  and GNAME63483(G63483,G75178,G75892);
  and GNAME63484(G63484,G75181,G75178);
  or GNAME63485(G63485,G63484,G63483,G63482);
  xor GNAME63495(G63495,G63496,G75895);
  xor GNAME63496(G63496,G75182,G75179);
  and GNAME63497(G63497,G75182,G75895);
  and GNAME63498(G63498,G75179,G75895);
  and GNAME63499(G63499,G75182,G75179);
  or GNAME63500(G63500,G63499,G63498,G63497);
  xor GNAME63510(G63510,G63511,G75898);
  xor GNAME63511(G63511,G75183,G75180);
  and GNAME63512(G63512,G75183,G75898);
  and GNAME63513(G63513,G75180,G75898);
  and GNAME63514(G63514,G75183,G75180);
  or GNAME63515(G63515,G63514,G63513,G63512);
  xor GNAME63525(G63525,G63526,G75901);
  xor GNAME63526(G63526,G75187,G75184);
  and GNAME63527(G63527,G75187,G75901);
  and GNAME63528(G63528,G75184,G75901);
  and GNAME63529(G63529,G75187,G75184);
  or GNAME63530(G63530,G63529,G63528,G63527);
  xor GNAME63540(G63540,G63541,G75904);
  xor GNAME63541(G63541,G75188,G75185);
  and GNAME63542(G63542,G75188,G75904);
  and GNAME63543(G63543,G75185,G75904);
  and GNAME63544(G63544,G75188,G75185);
  or GNAME63545(G63545,G63544,G63543,G63542);
  xor GNAME63555(G63555,G63556,G75907);
  xor GNAME63556(G63556,G75189,G75186);
  and GNAME63557(G63557,G75189,G75907);
  and GNAME63558(G63558,G75186,G75907);
  and GNAME63559(G63559,G75189,G75186);
  or GNAME63560(G63560,G63559,G63558,G63557);
  xor GNAME63570(G63570,G63571,G75910);
  xor GNAME63571(G63571,G75193,G75190);
  and GNAME63572(G63572,G75193,G75910);
  and GNAME63573(G63573,G75190,G75910);
  and GNAME63574(G63574,G75193,G75190);
  or GNAME63575(G63575,G63574,G63573,G63572);
  xor GNAME63585(G63585,G63586,G75913);
  xor GNAME63586(G63586,G75194,G75191);
  and GNAME63587(G63587,G75194,G75913);
  and GNAME63588(G63588,G75191,G75913);
  and GNAME63589(G63589,G75194,G75191);
  or GNAME63590(G63590,G63589,G63588,G63587);
  xor GNAME63600(G63600,G63601,G75916);
  xor GNAME63601(G63601,G75195,G75192);
  and GNAME63602(G63602,G75195,G75916);
  and GNAME63603(G63603,G75192,G75916);
  and GNAME63604(G63604,G75195,G75192);
  or GNAME63605(G63605,G63604,G63603,G63602);
  xor GNAME63615(G63615,G63616,G75919);
  xor GNAME63616(G63616,G75199,G75196);
  and GNAME63617(G63617,G75199,G75919);
  and GNAME63618(G63618,G75196,G75919);
  and GNAME63619(G63619,G75199,G75196);
  or GNAME63620(G63620,G63619,G63618,G63617);
  xor GNAME63630(G63630,G63631,G75922);
  xor GNAME63631(G63631,G75200,G75197);
  and GNAME63632(G63632,G75200,G75922);
  and GNAME63633(G63633,G75197,G75922);
  and GNAME63634(G63634,G75200,G75197);
  or GNAME63635(G63635,G63634,G63633,G63632);
  xor GNAME63645(G63645,G63646,G75925);
  xor GNAME63646(G63646,G75201,G75198);
  and GNAME63647(G63647,G75201,G75925);
  and GNAME63648(G63648,G75198,G75925);
  and GNAME63649(G63649,G75201,G75198);
  or GNAME63650(G63650,G63649,G63648,G63647);
  xor GNAME63660(G63660,G63661,G75928);
  xor GNAME63661(G63661,G75205,G75202);
  and GNAME63662(G63662,G75205,G75928);
  and GNAME63663(G63663,G75202,G75928);
  and GNAME63664(G63664,G75205,G75202);
  or GNAME63665(G63665,G63664,G63663,G63662);
  xor GNAME63675(G63675,G63676,G75931);
  xor GNAME63676(G63676,G75206,G75203);
  and GNAME63677(G63677,G75206,G75931);
  and GNAME63678(G63678,G75203,G75931);
  and GNAME63679(G63679,G75206,G75203);
  or GNAME63680(G63680,G63679,G63678,G63677);
  xor GNAME63690(G63690,G63691,G75934);
  xor GNAME63691(G63691,G75207,G75204);
  and GNAME63692(G63692,G75207,G75934);
  and GNAME63693(G63693,G75204,G75934);
  and GNAME63694(G63694,G75207,G75204);
  or GNAME63695(G63695,G63694,G63693,G63692);
  xor GNAME63705(G63705,G63706,G75937);
  xor GNAME63706(G63706,G75214,G75208);
  and GNAME63707(G63707,G75214,G75937);
  and GNAME63708(G63708,G75208,G75937);
  and GNAME63709(G63709,G75214,G75208);
  or GNAME63710(G63710,G63709,G63708,G63707);
  xor GNAME63720(G63720,G63721,G75940);
  xor GNAME63721(G63721,G75215,G75209);
  and GNAME63722(G63722,G75215,G75940);
  and GNAME63723(G63723,G75209,G75940);
  and GNAME63724(G63724,G75215,G75209);
  or GNAME63725(G63725,G63724,G63723,G63722);
  xor GNAME63735(G63735,G63736,G75943);
  xor GNAME63736(G63736,G75216,G75210);
  and GNAME63737(G63737,G75216,G75943);
  and GNAME63738(G63738,G75210,G75943);
  and GNAME63739(G63739,G75216,G75210);
  or GNAME63740(G63740,G63739,G63738,G63737);
  xor GNAME63750(G63750,G63751,G75946);
  xor GNAME63751(G63751,G75211,G77810);
  and GNAME63752(G63752,G75211,G75946);
  and GNAME63753(G63753,G77810,G75946);
  and GNAME63754(G63754,G75211,G77810);
  or GNAME63755(G63755,G63754,G63753,G63752);
  xor GNAME63765(G63765,G63766,G75949);
  xor GNAME63766(G63766,G75212,G77811);
  and GNAME63767(G63767,G75212,G75949);
  and GNAME63768(G63768,G77811,G75949);
  and GNAME63769(G63769,G75212,G77811);
  or GNAME63770(G63770,G63769,G63768,G63767);
  xor GNAME63780(G63780,G63781,G75952);
  xor GNAME63781(G63781,G75213,G77812);
  and GNAME63782(G63782,G75213,G75952);
  and GNAME63783(G63783,G77812,G75952);
  and GNAME63784(G63784,G75213,G77812);
  or GNAME63785(G63785,G63784,G63783,G63782);
  xor GNAME63795(G63795,G63796,G75955);
  xor GNAME63796(G63796,G74195,G75958);
  and GNAME63797(G63797,G74195,G75955);
  and GNAME63798(G63798,G75958,G75955);
  and GNAME63799(G63799,G74195,G75958);
  or GNAME63800(G63800,G63799,G63798,G63797);
  xor GNAME63810(G63810,G63811,G75961);
  xor GNAME63811(G63811,G74198,G75964);
  and GNAME63812(G63812,G74198,G75961);
  and GNAME63813(G63813,G75964,G75961);
  and GNAME63814(G63814,G74198,G75964);
  or GNAME63815(G63815,G63814,G63813,G63812);
  xor GNAME63825(G63825,G63826,G75967);
  xor GNAME63826(G63826,G74201,G75970);
  and GNAME63827(G63827,G74201,G75967);
  and GNAME63828(G63828,G75970,G75967);
  and GNAME63829(G63829,G74201,G75970);
  or GNAME63830(G63830,G63829,G63828,G63827);
  xor GNAME63840(G63840,G63841,G75973);
  xor GNAME63841(G63841,G74204,G75976);
  and GNAME63842(G63842,G74204,G75973);
  and GNAME63843(G63843,G75976,G75973);
  and GNAME63844(G63844,G74204,G75976);
  or GNAME63845(G63845,G63844,G63843,G63842);
  xor GNAME63855(G63855,G63856,G75979);
  xor GNAME63856(G63856,G74207,G75982);
  and GNAME63857(G63857,G74207,G75979);
  and GNAME63858(G63858,G75982,G75979);
  and GNAME63859(G63859,G74207,G75982);
  or GNAME63860(G63860,G63859,G63858,G63857);
  xor GNAME63870(G63870,G63871,G75985);
  xor GNAME63871(G63871,G74210,G75988);
  and GNAME63872(G63872,G74210,G75985);
  and GNAME63873(G63873,G75988,G75985);
  and GNAME63874(G63874,G74210,G75988);
  or GNAME63875(G63875,G63874,G63873,G63872);
  xor GNAME63885(G63885,G63886,G76027);
  xor GNAME63886(G63886,G74303,G76030);
  and GNAME63887(G63887,G74303,G76027);
  and GNAME63888(G63888,G76030,G76027);
  and GNAME63889(G63889,G74303,G76030);
  or GNAME63890(G63890,G63889,G63888,G63887);
  xor GNAME63900(G63900,G63901,G76033);
  xor GNAME63901(G63901,G74306,G76036);
  and GNAME63902(G63902,G74306,G76033);
  and GNAME63903(G63903,G76036,G76033);
  and GNAME63904(G63904,G74306,G76036);
  or GNAME63905(G63905,G63904,G63903,G63902);
  xor GNAME63915(G63915,G63916,G76039);
  xor GNAME63916(G63916,G74309,G76042);
  and GNAME63917(G63917,G74309,G76039);
  and GNAME63918(G63918,G76042,G76039);
  and GNAME63919(G63919,G74309,G76042);
  or GNAME63920(G63920,G63919,G63918,G63917);
  xor GNAME63930(G63930,G63931,G76063);
  xor GNAME63931(G63931,G74312,G76066);
  and GNAME63932(G63932,G74312,G76063);
  and GNAME63933(G63933,G76066,G76063);
  and GNAME63934(G63934,G74312,G76066);
  or GNAME63935(G63935,G63934,G63933,G63932);
  xor GNAME63945(G63945,G63946,G76069);
  xor GNAME63946(G63946,G74315,G76072);
  and GNAME63947(G63947,G74315,G76069);
  and GNAME63948(G63948,G76072,G76069);
  and GNAME63949(G63949,G74315,G76072);
  or GNAME63950(G63950,G63949,G63948,G63947);
  xor GNAME63960(G63960,G63961,G76075);
  xor GNAME63961(G63961,G74318,G76078);
  and GNAME63962(G63962,G74318,G76075);
  and GNAME63963(G63963,G76078,G76075);
  and GNAME63964(G63964,G74318,G76078);
  or GNAME63965(G63965,G63964,G63963,G63962);
  xor GNAME63975(G63975,G63976,G76099);
  xor GNAME63976(G63976,G74321,G76102);
  and GNAME63977(G63977,G74321,G76099);
  and GNAME63978(G63978,G76102,G76099);
  and GNAME63979(G63979,G74321,G76102);
  or GNAME63980(G63980,G63979,G63978,G63977);
  xor GNAME63990(G63990,G63991,G76105);
  xor GNAME63991(G63991,G74324,G76108);
  and GNAME63992(G63992,G74324,G76105);
  and GNAME63993(G63993,G76108,G76105);
  and GNAME63994(G63994,G74324,G76108);
  or GNAME63995(G63995,G63994,G63993,G63992);
  xor GNAME64005(G64005,G64006,G76111);
  xor GNAME64006(G64006,G74327,G76114);
  and GNAME64007(G64007,G74327,G76111);
  and GNAME64008(G64008,G76114,G76111);
  and GNAME64009(G64009,G74327,G76114);
  or GNAME64010(G64010,G64009,G64008,G64007);
  xor GNAME64020(G64020,G64021,G76135);
  xor GNAME64021(G64021,G74330,G76138);
  and GNAME64022(G64022,G74330,G76135);
  and GNAME64023(G64023,G76138,G76135);
  and GNAME64024(G64024,G74330,G76138);
  or GNAME64025(G64025,G64024,G64023,G64022);
  xor GNAME64035(G64035,G64036,G76141);
  xor GNAME64036(G64036,G74333,G76144);
  and GNAME64037(G64037,G74333,G76141);
  and GNAME64038(G64038,G76144,G76141);
  and GNAME64039(G64039,G74333,G76144);
  or GNAME64040(G64040,G64039,G64038,G64037);
  xor GNAME64050(G64050,G64051,G76147);
  xor GNAME64051(G64051,G74336,G76150);
  and GNAME64052(G64052,G74336,G76147);
  and GNAME64053(G64053,G76150,G76147);
  and GNAME64054(G64054,G74336,G76150);
  or GNAME64055(G64055,G64054,G64053,G64052);
  xor GNAME64065(G64065,G64066,G74470);
  xor GNAME64066(G64066,G76153,G76156);
  and GNAME64067(G64067,G76153,G74470);
  and GNAME64068(G64068,G76156,G74470);
  and GNAME64069(G64069,G76153,G76156);
  or GNAME64070(G64070,G64069,G64068,G64067);
  xor GNAME64080(G64080,G64081,G74476);
  xor GNAME64081(G64081,G76159,G76162);
  and GNAME64082(G64082,G76159,G74476);
  and GNAME64083(G64083,G76162,G74476);
  and GNAME64084(G64084,G76159,G76162);
  or GNAME64085(G64085,G64084,G64083,G64082);
  xor GNAME64095(G64095,G64096,G74482);
  xor GNAME64096(G64096,G76165,G76168);
  and GNAME64097(G64097,G76165,G74482);
  and GNAME64098(G64098,G76168,G74482);
  and GNAME64099(G64099,G76165,G76168);
  or GNAME64100(G64100,G64099,G64098,G64097);
  xor GNAME64110(G64110,G64111,G76171);
  xor GNAME64111(G64111,G74339,G76174);
  and GNAME64112(G64112,G74339,G76171);
  and GNAME64113(G64113,G76174,G76171);
  and GNAME64114(G64114,G74339,G76174);
  or GNAME64115(G64115,G64114,G64113,G64112);
  xor GNAME64125(G64125,G64126,G76177);
  xor GNAME64126(G64126,G74342,G76180);
  and GNAME64127(G64127,G74342,G76177);
  and GNAME64128(G64128,G76180,G76177);
  and GNAME64129(G64129,G74342,G76180);
  or GNAME64130(G64130,G64129,G64128,G64127);
  xor GNAME64140(G64140,G64141,G76183);
  xor GNAME64141(G64141,G74345,G76186);
  and GNAME64142(G64142,G74345,G76183);
  and GNAME64143(G64143,G76186,G76183);
  and GNAME64144(G64144,G74345,G76186);
  or GNAME64145(G64145,G64144,G64143,G64142);
  xor GNAME64155(G64155,G64156,G63485);
  xor GNAME64156(G64156,G77792,G76225);
  and GNAME64157(G64157,G77792,G63485);
  and GNAME64158(G64158,G76225,G63485);
  and GNAME64159(G64159,G77792,G76225);
  or GNAME64160(G64160,G64159,G64158,G64157);
  xor GNAME64170(G64170,G64171,G63500);
  xor GNAME64171(G64171,G77793,G76228);
  and GNAME64172(G64172,G77793,G63500);
  and GNAME64173(G64173,G76228,G63500);
  and GNAME64174(G64174,G77793,G76228);
  or GNAME64175(G64175,G64174,G64173,G64172);
  xor GNAME64185(G64185,G64186,G63515);
  xor GNAME64186(G64186,G77794,G76231);
  and GNAME64187(G64187,G77794,G63515);
  and GNAME64188(G64188,G76231,G63515);
  and GNAME64189(G64189,G77794,G76231);
  or GNAME64190(G64190,G64189,G64188,G64187);
  xor GNAME64200(G64200,G64201,G63480);
  xor GNAME64201(G64201,G75849,G64295);
  and GNAME64202(G64202,G75849,G63480);
  and GNAME64203(G64203,G64295,G63480);
  and GNAME64204(G64204,G75849,G64295);
  or GNAME64205(G64205,G64204,G64203,G64202);
  xor GNAME64215(G64215,G64216,G63495);
  xor GNAME64216(G64216,G75851,G64310);
  and GNAME64217(G64217,G75851,G63495);
  and GNAME64218(G64218,G64310,G63495);
  and GNAME64219(G64219,G75851,G64310);
  or GNAME64220(G64220,G64219,G64218,G64217);
  xor GNAME64230(G64230,G64231,G63510);
  xor GNAME64231(G64231,G75853,G64325);
  and GNAME64232(G64232,G75853,G63510);
  and GNAME64233(G64233,G64325,G63510);
  and GNAME64234(G64234,G75853,G64325);
  or GNAME64235(G64235,G64234,G64233,G64232);
  xor GNAME64245(G64245,G64246,G64340);
  xor GNAME64246(G64246,G63530,G64290);
  and GNAME64247(G64247,G63530,G64340);
  and GNAME64248(G64248,G64290,G64340);
  and GNAME64249(G64249,G63530,G64290);
  or GNAME64250(G64250,G64249,G64248,G64247);
  xor GNAME64260(G64260,G64261,G64355);
  xor GNAME64261(G64261,G63545,G64305);
  and GNAME64262(G64262,G63545,G64355);
  and GNAME64263(G64263,G64305,G64355);
  and GNAME64264(G64264,G63545,G64305);
  or GNAME64265(G64265,G64264,G64263,G64262);
  xor GNAME64275(G64275,G64276,G64370);
  xor GNAME64276(G64276,G63560,G64320);
  and GNAME64277(G64277,G63560,G64370);
  and GNAME64278(G64278,G64320,G64370);
  and GNAME64279(G64279,G63560,G64320);
  or GNAME64280(G64280,G64279,G64278,G64277);
  xor GNAME64290(G64290,G64291,G76237);
  xor GNAME64291(G64291,G77795,G76234);
  and GNAME64292(G64292,G77795,G76237);
  and GNAME64293(G64293,G76234,G76237);
  and GNAME64294(G64294,G77795,G76234);
  or GNAME64295(G64295,G64294,G64293,G64292);
  xor GNAME64305(G64305,G64306,G76243);
  xor GNAME64306(G64306,G77796,G76240);
  and GNAME64307(G64307,G77796,G76243);
  and GNAME64308(G64308,G76240,G76243);
  and GNAME64309(G64309,G77796,G76240);
  or GNAME64310(G64310,G64309,G64308,G64307);
  xor GNAME64320(G64320,G64321,G76249);
  xor GNAME64321(G64321,G77797,G76246);
  and GNAME64322(G64322,G77797,G76249);
  and GNAME64323(G64323,G76246,G76249);
  and GNAME64324(G64324,G77797,G76246);
  or GNAME64325(G64325,G64324,G64323,G64322);
  xor GNAME64335(G64335,G64336,G64475);
  xor GNAME64336(G64336,G76252,G75855);
  and GNAME64337(G64337,G76252,G64475);
  and GNAME64338(G64338,G75855,G64475);
  and GNAME64339(G64339,G76252,G75855);
  or GNAME64340(G64340,G64339,G64338,G64337);
  xor GNAME64350(G64350,G64351,G64490);
  xor GNAME64351(G64351,G76255,G75857);
  and GNAME64352(G64352,G76255,G64490);
  and GNAME64353(G64353,G75857,G64490);
  and GNAME64354(G64354,G76255,G75857);
  or GNAME64355(G64355,G64354,G64353,G64352);
  xor GNAME64365(G64365,G64366,G64505);
  xor GNAME64366(G64366,G76258,G75859);
  and GNAME64367(G64367,G76258,G64505);
  and GNAME64368(G64368,G75859,G64505);
  and GNAME64369(G64369,G76258,G75859);
  or GNAME64370(G64370,G64369,G64368,G64367);
  xor GNAME64380(G64380,G64381,G64335);
  xor GNAME64381(G64381,G63525,G64430);
  and GNAME64382(G64382,G63525,G64335);
  and GNAME64383(G64383,G64430,G64335);
  and GNAME64384(G64384,G63525,G64430);
  or GNAME64385(G64385,G64384,G64383,G64382);
  xor GNAME64395(G64395,G64396,G64350);
  xor GNAME64396(G64396,G63540,G64445);
  and GNAME64397(G64397,G63540,G64350);
  and GNAME64398(G64398,G64445,G64350);
  and GNAME64399(G64399,G63540,G64445);
  or GNAME64400(G64400,G64399,G64398,G64397);
  xor GNAME64410(G64410,G64411,G64365);
  xor GNAME64411(G64411,G63555,G64460);
  and GNAME64412(G64412,G63555,G64365);
  and GNAME64413(G64413,G64460,G64365);
  and GNAME64414(G64414,G63555,G64460);
  or GNAME64415(G64415,G64414,G64413,G64412);
  xor GNAME64425(G64425,G64426,G64520);
  xor GNAME64426(G64426,G76261,G63575);
  and GNAME64427(G64427,G76261,G64520);
  and GNAME64428(G64428,G63575,G64520);
  and GNAME64429(G64429,G76261,G63575);
  or GNAME64430(G64430,G64429,G64428,G64427);
  xor GNAME64440(G64440,G64441,G64535);
  xor GNAME64441(G64441,G76264,G63590);
  and GNAME64442(G64442,G76264,G64535);
  and GNAME64443(G64443,G63590,G64535);
  and GNAME64444(G64444,G76264,G63590);
  or GNAME64445(G64445,G64444,G64443,G64442);
  xor GNAME64455(G64455,G64456,G64550);
  xor GNAME64456(G64456,G76267,G63605);
  and GNAME64457(G64457,G76267,G64550);
  and GNAME64458(G64458,G63605,G64550);
  and GNAME64459(G64459,G76267,G63605);
  or GNAME64460(G64460,G64459,G64458,G64457);
  xor GNAME64470(G64470,G64471,G76273);
  xor GNAME64471(G64471,G77798,G76270);
  and GNAME64472(G64472,G77798,G76273);
  and GNAME64473(G64473,G76270,G76273);
  and GNAME64474(G64474,G77798,G76270);
  or GNAME64475(G64475,G64474,G64473,G64472);
  xor GNAME64485(G64485,G64486,G76279);
  xor GNAME64486(G64486,G77799,G76276);
  and GNAME64487(G64487,G77799,G76279);
  and GNAME64488(G64488,G76276,G76279);
  and GNAME64489(G64489,G77799,G76276);
  or GNAME64490(G64490,G64489,G64488,G64487);
  xor GNAME64500(G64500,G64501,G76285);
  xor GNAME64501(G64501,G77800,G76282);
  and GNAME64502(G64502,G77800,G76285);
  and GNAME64503(G64503,G76282,G76285);
  and GNAME64504(G64504,G77800,G76282);
  or GNAME64505(G64505,G64504,G64503,G64502);
  xor GNAME64515(G64515,G64516,G75861);
  xor GNAME64516(G64516,G76288,G76291);
  and GNAME64517(G64517,G76288,G75861);
  and GNAME64518(G64518,G76291,G75861);
  and GNAME64519(G64519,G76288,G76291);
  or GNAME64520(G64520,G64519,G64518,G64517);
  xor GNAME64530(G64530,G64531,G75863);
  xor GNAME64531(G64531,G76294,G76297);
  and GNAME64532(G64532,G76294,G75863);
  and GNAME64533(G64533,G76297,G75863);
  and GNAME64534(G64534,G76294,G76297);
  or GNAME64535(G64535,G64534,G64533,G64532);
  xor GNAME64545(G64545,G64546,G75865);
  xor GNAME64546(G64546,G76300,G76303);
  and GNAME64547(G64547,G76300,G75865);
  and GNAME64548(G64548,G76303,G75865);
  and GNAME64549(G64549,G76300,G76303);
  or GNAME64550(G64550,G64549,G64548,G64547);
  xor GNAME64560(G64560,G64561,G64515);
  xor GNAME64561(G64561,G64610,G63570);
  and GNAME64562(G64562,G64610,G64515);
  and GNAME64563(G64563,G63570,G64515);
  and GNAME64564(G64564,G64610,G63570);
  or GNAME64565(G64565,G64564,G64563,G64562);
  xor GNAME64575(G64575,G64576,G64530);
  xor GNAME64576(G64576,G64625,G63585);
  and GNAME64577(G64577,G64625,G64530);
  and GNAME64578(G64578,G63585,G64530);
  and GNAME64579(G64579,G64625,G63585);
  or GNAME64580(G64580,G64579,G64578,G64577);
  xor GNAME64590(G64590,G64591,G64545);
  xor GNAME64591(G64591,G64640,G63600);
  and GNAME64592(G64592,G64640,G64545);
  and GNAME64593(G64593,G63600,G64545);
  and GNAME64594(G64594,G64640,G63600);
  or GNAME64595(G64595,G64594,G64593,G64592);
  xor GNAME64605(G64605,G64606,G76309);
  xor GNAME64606(G64606,G77801,G76306);
  and GNAME64607(G64607,G77801,G76309);
  and GNAME64608(G64608,G76306,G76309);
  and GNAME64609(G64609,G77801,G76306);
  or GNAME64610(G64610,G64609,G64608,G64607);
  xor GNAME64620(G64620,G64621,G76315);
  xor GNAME64621(G64621,G77802,G76312);
  and GNAME64622(G64622,G77802,G76315);
  and GNAME64623(G64623,G76312,G76315);
  and GNAME64624(G64624,G77802,G76312);
  or GNAME64625(G64625,G64624,G64623,G64622);
  xor GNAME64635(G64635,G64636,G76321);
  xor GNAME64636(G64636,G77803,G76318);
  and GNAME64637(G64637,G77803,G76321);
  and GNAME64638(G64638,G76318,G76321);
  and GNAME64639(G64639,G77803,G76318);
  or GNAME64640(G64640,G64639,G64638,G64637);
  xor GNAME64650(G64650,G64651,G63620);
  xor GNAME64651(G64651,G76324,G76327);
  and GNAME64652(G64652,G76324,G63620);
  and GNAME64653(G64653,G76327,G63620);
  and GNAME64654(G64654,G76324,G76327);
  or GNAME64655(G64655,G64654,G64653,G64652);
  xor GNAME64665(G64665,G64666,G63635);
  xor GNAME64666(G64666,G76330,G76333);
  and GNAME64667(G64667,G76330,G63635);
  and GNAME64668(G64668,G76333,G63635);
  and GNAME64669(G64669,G76330,G76333);
  or GNAME64670(G64670,G64669,G64668,G64667);
  xor GNAME64680(G64680,G64681,G63650);
  xor GNAME64681(G64681,G76336,G76339);
  and GNAME64682(G64682,G76336,G63650);
  and GNAME64683(G64683,G76339,G63650);
  and GNAME64684(G64684,G76336,G76339);
  or GNAME64685(G64685,G64684,G64683,G64682);
  xor GNAME64695(G64695,G64696,G64790);
  xor GNAME64696(G64696,G63615,G64920);
  and GNAME64697(G64697,G63615,G64790);
  and GNAME64698(G64698,G64920,G64790);
  and GNAME64699(G64699,G63615,G64920);
  or GNAME64700(G64700,G64699,G64698,G64697);
  xor GNAME64710(G64710,G64711,G64805);
  xor GNAME64711(G64711,G63630,G64935);
  and GNAME64712(G64712,G63630,G64805);
  and GNAME64713(G64713,G64935,G64805);
  and GNAME64714(G64714,G63630,G64935);
  or GNAME64715(G64715,G64714,G64713,G64712);
  xor GNAME64725(G64725,G64726,G64820);
  xor GNAME64726(G64726,G63645,G64950);
  and GNAME64727(G64727,G63645,G64820);
  and GNAME64728(G64728,G64950,G64820);
  and GNAME64729(G64729,G63645,G64950);
  or GNAME64730(G64730,G64729,G64728,G64727);
  xor GNAME64740(G64740,G64741,G76345);
  xor GNAME64741(G64741,G77804,G76342);
  and GNAME64742(G64742,G77804,G76345);
  and GNAME64743(G64743,G76342,G76345);
  and GNAME64744(G64744,G77804,G76342);
  or GNAME64745(G64745,G64744,G64743,G64742);
  xor GNAME64755(G64755,G64756,G76351);
  xor GNAME64756(G64756,G77805,G76348);
  and GNAME64757(G64757,G77805,G76351);
  and GNAME64758(G64758,G76348,G76351);
  and GNAME64759(G64759,G77805,G76348);
  or GNAME64760(G64760,G64759,G64758,G64757);
  xor GNAME64770(G64770,G64771,G76357);
  xor GNAME64771(G64771,G77806,G76354);
  and GNAME64772(G64772,G77806,G76357);
  and GNAME64773(G64773,G76354,G76357);
  and GNAME64774(G64774,G77806,G76354);
  or GNAME64775(G64775,G64774,G64773,G64772);
  xor GNAME64785(G64785,G64786,G64740);
  xor GNAME64786(G64786,G63665,G64970);
  and GNAME64787(G64787,G63665,G64740);
  and GNAME64788(G64788,G64970,G64740);
  and GNAME64789(G64789,G63665,G64970);
  or GNAME64790(G64790,G64789,G64788,G64787);
  xor GNAME64800(G64800,G64801,G64755);
  xor GNAME64801(G64801,G63680,G64985);
  and GNAME64802(G64802,G63680,G64755);
  and GNAME64803(G64803,G64985,G64755);
  and GNAME64804(G64804,G63680,G64985);
  or GNAME64805(G64805,G64804,G64803,G64802);
  xor GNAME64815(G64815,G64816,G64770);
  xor GNAME64816(G64816,G63695,G65000);
  and GNAME64817(G64817,G63695,G64770);
  and GNAME64818(G64818,G65000,G64770);
  and GNAME64819(G64819,G63695,G65000);
  or GNAME64820(G64820,G64819,G64818,G64817);
  xor GNAME64830(G64830,G64831,G64880);
  xor GNAME64831(G64831,G76360,G64745);
  and GNAME64832(G64832,G76360,G64880);
  and GNAME64833(G64833,G64745,G64880);
  and GNAME64834(G64834,G76360,G64745);
  or GNAME64835(G64835,G64834,G64833,G64832);
  xor GNAME64845(G64845,G64846,G64895);
  xor GNAME64846(G64846,G76363,G64760);
  and GNAME64847(G64847,G76363,G64895);
  and GNAME64848(G64848,G64760,G64895);
  and GNAME64849(G64849,G76363,G64760);
  or GNAME64850(G64850,G64849,G64848,G64847);
  xor GNAME64860(G64860,G64861,G64910);
  xor GNAME64861(G64861,G76366,G64775);
  and GNAME64862(G64862,G76366,G64910);
  and GNAME64863(G64863,G64775,G64910);
  and GNAME64864(G64864,G76366,G64775);
  or GNAME64865(G64865,G64864,G64863,G64862);
  xor GNAME64875(G64875,G64876,G76375);
  xor GNAME64876(G64876,G76369,G76372);
  and GNAME64877(G64877,G76369,G76375);
  and GNAME64878(G64878,G76372,G76375);
  and GNAME64879(G64879,G76369,G76372);
  or GNAME64880(G64880,G64879,G64878,G64877);
  xor GNAME64890(G64890,G64891,G76384);
  xor GNAME64891(G64891,G76378,G76381);
  and GNAME64892(G64892,G76378,G76384);
  and GNAME64893(G64893,G76381,G76384);
  and GNAME64894(G64894,G76378,G76381);
  or GNAME64895(G64895,G64894,G64893,G64892);
  xor GNAME64905(G64905,G64906,G76393);
  xor GNAME64906(G64906,G76387,G76390);
  and GNAME64907(G64907,G76387,G76393);
  and GNAME64908(G64908,G76390,G76393);
  and GNAME64909(G64909,G76387,G76390);
  or GNAME64910(G64910,G64909,G64908,G64907);
  xor GNAME64920(G64920,G64921,G75867);
  xor GNAME64921(G64921,G76396,G76399);
  and GNAME64922(G64922,G76396,G75867);
  and GNAME64923(G64923,G76399,G75867);
  and GNAME64924(G64924,G76396,G76399);
  or GNAME64925(G64925,G64924,G64923,G64922);
  xor GNAME64935(G64935,G64936,G75869);
  xor GNAME64936(G64936,G76402,G76405);
  and GNAME64937(G64937,G76402,G75869);
  and GNAME64938(G64938,G76405,G75869);
  and GNAME64939(G64939,G76402,G76405);
  or GNAME64940(G64940,G64939,G64938,G64937);
  xor GNAME64950(G64950,G64951,G75871);
  xor GNAME64951(G64951,G76408,G76411);
  and GNAME64952(G64952,G76408,G75871);
  and GNAME64953(G64953,G76411,G75871);
  and GNAME64954(G64954,G76408,G76411);
  or GNAME64955(G64955,G64954,G64953,G64952);
  xor GNAME64965(G64965,G64966,G75873);
  xor GNAME64966(G64966,G76414,G76417);
  and GNAME64967(G64967,G76414,G75873);
  and GNAME64968(G64968,G76417,G75873);
  and GNAME64969(G64969,G76414,G76417);
  or GNAME64970(G64970,G64969,G64968,G64967);
  xor GNAME64980(G64980,G64981,G75875);
  xor GNAME64981(G64981,G76420,G76423);
  and GNAME64982(G64982,G76420,G75875);
  and GNAME64983(G64983,G76423,G75875);
  and GNAME64984(G64984,G76420,G76423);
  or GNAME64985(G64985,G64984,G64983,G64982);
  xor GNAME64995(G64995,G64996,G75877);
  xor GNAME64996(G64996,G76426,G76429);
  and GNAME64997(G64997,G76426,G75877);
  and GNAME64998(G64998,G76429,G75877);
  and GNAME64999(G64999,G76426,G76429);
  or GNAME65000(G65000,G64999,G64998,G64997);
  xor GNAME65010(G65010,G65011,G65060);
  xor GNAME65011(G65011,G76432,G76435);
  and GNAME65012(G65012,G76432,G65060);
  and GNAME65013(G65013,G76435,G65060);
  and GNAME65014(G65014,G76432,G76435);
  or GNAME65015(G65015,G65014,G65013,G65012);
  xor GNAME65025(G65025,G65026,G65075);
  xor GNAME65026(G65026,G76438,G76441);
  and GNAME65027(G65027,G76438,G65075);
  and GNAME65028(G65028,G76441,G65075);
  and GNAME65029(G65029,G76438,G76441);
  or GNAME65030(G65030,G65029,G65028,G65027);
  xor GNAME65040(G65040,G65041,G65090);
  xor GNAME65041(G65041,G76444,G76447);
  and GNAME65042(G65042,G76444,G65090);
  and GNAME65043(G65043,G76447,G65090);
  and GNAME65044(G65044,G76444,G76447);
  or GNAME65045(G65045,G65044,G65043,G65042);
  xor GNAME65055(G65055,G65056,G76453);
  xor GNAME65056(G65056,G77807,G76450);
  and GNAME65057(G65057,G77807,G76453);
  and GNAME65058(G65058,G76450,G76453);
  and GNAME65059(G65059,G77807,G76450);
  or GNAME65060(G65060,G65059,G65058,G65057);
  xor GNAME65070(G65070,G65071,G76459);
  xor GNAME65071(G65071,G77808,G76456);
  and GNAME65072(G65072,G77808,G76459);
  and GNAME65073(G65073,G76456,G76459);
  and GNAME65074(G65074,G77808,G76456);
  or GNAME65075(G65075,G65074,G65073,G65072);
  xor GNAME65085(G65085,G65086,G76465);
  xor GNAME65086(G65086,G77809,G76462);
  and GNAME65087(G65087,G77809,G76465);
  and GNAME65088(G65088,G76462,G76465);
  and GNAME65089(G65089,G77809,G76462);
  or GNAME65090(G65090,G65089,G65088,G65087);
  xor GNAME65100(G65100,G65101,G64965);
  xor GNAME65101(G65101,G65150,G63660);
  and GNAME65102(G65102,G65150,G64965);
  and GNAME65103(G65103,G63660,G64965);
  and GNAME65104(G65104,G65150,G63660);
  or GNAME65105(G65105,G65104,G65103,G65102);
  xor GNAME65115(G65115,G65116,G64980);
  xor GNAME65116(G65116,G65165,G63675);
  and GNAME65117(G65117,G65165,G64980);
  and GNAME65118(G65118,G63675,G64980);
  and GNAME65119(G65119,G65165,G63675);
  or GNAME65120(G65120,G65119,G65118,G65117);
  xor GNAME65130(G65130,G65131,G64995);
  xor GNAME65131(G65131,G65180,G63690);
  and GNAME65132(G65132,G65180,G64995);
  and GNAME65133(G65133,G63690,G64995);
  and GNAME65134(G65134,G65180,G63690);
  or GNAME65135(G65135,G65134,G65133,G65132);
  xor GNAME65145(G65145,G65146,G76474);
  xor GNAME65146(G65146,G76468,G76471);
  and GNAME65147(G65147,G76468,G76474);
  and GNAME65148(G65148,G76471,G76474);
  and GNAME65149(G65149,G76468,G76471);
  or GNAME65150(G65150,G65149,G65148,G65147);
  xor GNAME65160(G65160,G65161,G76483);
  xor GNAME65161(G65161,G76477,G76480);
  and GNAME65162(G65162,G76477,G76483);
  and GNAME65163(G65163,G76480,G76483);
  and GNAME65164(G65164,G76477,G76480);
  or GNAME65165(G65165,G65164,G65163,G65162);
  xor GNAME65175(G65175,G65176,G76492);
  xor GNAME65176(G65176,G76486,G76489);
  and GNAME65177(G65177,G76486,G76492);
  and GNAME65178(G65178,G76489,G76492);
  and GNAME65179(G65179,G76486,G76489);
  or GNAME65180(G65180,G65179,G65178,G65177);
  xor GNAME65190(G65190,G65191,G75879);
  xor GNAME65191(G65191,G76495,G76498);
  and GNAME65192(G65192,G76495,G75879);
  and GNAME65193(G65193,G76498,G75879);
  and GNAME65194(G65194,G76495,G76498);
  or GNAME65195(G65195,G65194,G65193,G65192);
  xor GNAME65205(G65205,G65206,G75881);
  xor GNAME65206(G65206,G76501,G76504);
  and GNAME65207(G65207,G76501,G75881);
  and GNAME65208(G65208,G76504,G75881);
  and GNAME65209(G65209,G76501,G76504);
  or GNAME65210(G65210,G65209,G65208,G65207);
  xor GNAME65220(G65220,G65221,G75883);
  xor GNAME65221(G65221,G76507,G76510);
  and GNAME65222(G65222,G76507,G75883);
  and GNAME65223(G65223,G76510,G75883);
  and GNAME65224(G65224,G76507,G76510);
  or GNAME65225(G65225,G65224,G65223,G65222);
  xor GNAME65235(G65235,G65236,G65195);
  xor GNAME65236(G65236,G76513,G63710);
  and GNAME65237(G65237,G76513,G65195);
  and GNAME65238(G65238,G63710,G65195);
  and GNAME65239(G65239,G76513,G63710);
  or GNAME65240(G65240,G65239,G65238,G65237);
  xor GNAME65250(G65250,G65251,G65345);
  xor GNAME65251(G65251,G63755,G65510);
  and GNAME65252(G65252,G63755,G65345);
  and GNAME65253(G65253,G65510,G65345);
  and GNAME65254(G65254,G63755,G65510);
  or GNAME65255(G65255,G65254,G65253,G65252);
  xor GNAME65265(G65265,G65266,G65210);
  xor GNAME65266(G65266,G76516,G63725);
  and GNAME65267(G65267,G76516,G65210);
  and GNAME65268(G65268,G63725,G65210);
  and GNAME65269(G65269,G76516,G63725);
  or GNAME65270(G65270,G65269,G65268,G65267);
  xor GNAME65280(G65280,G65281,G65225);
  xor GNAME65281(G65281,G76519,G63740);
  and GNAME65282(G65282,G76519,G65225);
  and GNAME65283(G65283,G63740,G65225);
  and GNAME65284(G65284,G76519,G63740);
  or GNAME65285(G65285,G65284,G65283,G65282);
  xor GNAME65295(G65295,G65296,G65390);
  xor GNAME65296(G65296,G63770,G65525);
  and GNAME65297(G65297,G63770,G65390);
  and GNAME65298(G65298,G65525,G65390);
  and GNAME65299(G65299,G63770,G65525);
  or GNAME65300(G65300,G65299,G65298,G65297);
  xor GNAME65310(G65310,G65311,G65405);
  xor GNAME65311(G65311,G63785,G65540);
  and GNAME65312(G65312,G63785,G65405);
  and GNAME65313(G65313,G65540,G65405);
  and GNAME65314(G65314,G63785,G65540);
  or GNAME65315(G65315,G65314,G65313,G65312);
  xor GNAME65325(G65325,G65326,G76528);
  xor GNAME65326(G65326,G76522,G76525);
  and GNAME65327(G65327,G76522,G76528);
  and GNAME65328(G65328,G76525,G76528);
  and GNAME65329(G65329,G76522,G76525);
  or GNAME65330(G65330,G65329,G65328,G65327);
  xor GNAME65340(G65340,G65341,G76537);
  xor GNAME65341(G65341,G76531,G76534);
  and GNAME65342(G65342,G76531,G76537);
  and GNAME65343(G65343,G76534,G76537);
  and GNAME65344(G65344,G76531,G76534);
  or GNAME65345(G65345,G65344,G65343,G65342);
  xor GNAME65355(G65355,G65356,G76546);
  xor GNAME65356(G65356,G76540,G76543);
  and GNAME65357(G65357,G76540,G76546);
  and GNAME65358(G65358,G76543,G76546);
  and GNAME65359(G65359,G76540,G76543);
  or GNAME65360(G65360,G65359,G65358,G65357);
  xor GNAME65370(G65370,G65371,G76555);
  xor GNAME65371(G65371,G76549,G76552);
  and GNAME65372(G65372,G76549,G76555);
  and GNAME65373(G65373,G76552,G76555);
  and GNAME65374(G65374,G76549,G76552);
  or GNAME65375(G65375,G65374,G65373,G65372);
  xor GNAME65385(G65385,G65386,G76564);
  xor GNAME65386(G65386,G76558,G76561);
  and GNAME65387(G65387,G76558,G76564);
  and GNAME65388(G65388,G76561,G76564);
  and GNAME65389(G65389,G76558,G76561);
  or GNAME65390(G65390,G65389,G65388,G65387);
  xor GNAME65400(G65400,G65401,G76573);
  xor GNAME65401(G65401,G76567,G76570);
  and GNAME65402(G65402,G76567,G76573);
  and GNAME65403(G65403,G76570,G76573);
  and GNAME65404(G65404,G76567,G76570);
  or GNAME65405(G65405,G65404,G65403,G65402);
  xor GNAME65415(G65415,G65416,G65190);
  xor GNAME65416(G65416,G63705,G65325);
  and GNAME65417(G65417,G63705,G65190);
  and GNAME65418(G65418,G65325,G65190);
  and GNAME65419(G65419,G63705,G65325);
  or GNAME65420(G65420,G65419,G65418,G65417);
  xor GNAME65430(G65430,G65431,G65505);
  xor GNAME65431(G65431,G63750,G65340);
  and GNAME65432(G65432,G63750,G65505);
  and GNAME65433(G65433,G65340,G65505);
  and GNAME65434(G65434,G63750,G65340);
  or GNAME65435(G65435,G65434,G65433,G65432);
  xor GNAME65445(G65445,G65446,G65205);
  xor GNAME65446(G65446,G63720,G65355);
  and GNAME65447(G65447,G63720,G65205);
  and GNAME65448(G65448,G65355,G65205);
  and GNAME65449(G65449,G63720,G65355);
  or GNAME65450(G65450,G65449,G65448,G65447);
  xor GNAME65460(G65460,G65461,G65520);
  xor GNAME65461(G65461,G63765,G65385);
  and GNAME65462(G65462,G63765,G65520);
  and GNAME65463(G65463,G65385,G65520);
  and GNAME65464(G65464,G63765,G65385);
  or GNAME65465(G65465,G65464,G65463,G65462);
  xor GNAME65475(G65475,G65476,G65220);
  xor GNAME65476(G65476,G63735,G65370);
  and GNAME65477(G65477,G63735,G65220);
  and GNAME65478(G65478,G65370,G65220);
  and GNAME65479(G65479,G63735,G65370);
  or GNAME65480(G65480,G65479,G65478,G65477);
  xor GNAME65490(G65490,G65491,G65535);
  xor GNAME65491(G65491,G63780,G65400);
  and GNAME65492(G65492,G63780,G65535);
  and GNAME65493(G65493,G65400,G65535);
  and GNAME65494(G65494,G63780,G65400);
  or GNAME65495(G65495,G65494,G65493,G65492);
  xor GNAME65505(G65505,G65506,G76582);
  xor GNAME65506(G65506,G76576,G76579);
  and GNAME65507(G65507,G76576,G76582);
  and GNAME65508(G65508,G76579,G76582);
  and GNAME65509(G65509,G76576,G76579);
  or GNAME65510(G65510,G65509,G65508,G65507);
  xor GNAME65520(G65520,G65521,G76591);
  xor GNAME65521(G65521,G76585,G76588);
  and GNAME65522(G65522,G76585,G76591);
  and GNAME65523(G65523,G76588,G76591);
  and GNAME65524(G65524,G76585,G76588);
  or GNAME65525(G65525,G65524,G65523,G65522);
  xor GNAME65535(G65535,G65536,G76600);
  xor GNAME65536(G65536,G76594,G76597);
  and GNAME65537(G65537,G76594,G76600);
  and GNAME65538(G65538,G76597,G76600);
  and GNAME65539(G65539,G76594,G76597);
  or GNAME65540(G65540,G65539,G65538,G65537);
  xor GNAME65550(G65550,G65551,G75885);
  xor GNAME65551(G65551,G76603,G76606);
  and GNAME65552(G65552,G76603,G75885);
  and GNAME65553(G65553,G76606,G75885);
  and GNAME65554(G65554,G76603,G76606);
  or GNAME65555(G65555,G65554,G65553,G65552);
  xor GNAME65565(G65565,G65566,G75887);
  xor GNAME65566(G65566,G76609,G76612);
  and GNAME65567(G65567,G76609,G75887);
  and GNAME65568(G65568,G76612,G75887);
  and GNAME65569(G65569,G76609,G76612);
  or GNAME65570(G65570,G65569,G65568,G65567);
  xor GNAME65580(G65580,G65581,G75889);
  xor GNAME65581(G65581,G76615,G76618);
  and GNAME65582(G65582,G76615,G75889);
  and GNAME65583(G65583,G76618,G75889);
  and GNAME65584(G65584,G76615,G76618);
  or GNAME65585(G65585,G65584,G65583,G65582);
  xor GNAME65595(G65595,G65596,G76627);
  xor GNAME65596(G65596,G76621,G76624);
  and GNAME65597(G65597,G76621,G76627);
  and GNAME65598(G65598,G76624,G76627);
  and GNAME65599(G65599,G76621,G76624);
  or GNAME65600(G65600,G65599,G65598,G65597);
  xor GNAME65610(G65610,G65611,G76636);
  xor GNAME65611(G65611,G76630,G76633);
  and GNAME65612(G65612,G76630,G76636);
  and GNAME65613(G65613,G76633,G76636);
  and GNAME65614(G65614,G76630,G76633);
  or GNAME65615(G65615,G65614,G65613,G65612);
  xor GNAME65625(G65625,G65626,G76645);
  xor GNAME65626(G65626,G76639,G76642);
  and GNAME65627(G65627,G76639,G76645);
  and GNAME65628(G65628,G76642,G76645);
  and GNAME65629(G65629,G76639,G76642);
  or GNAME65630(G65630,G65629,G65628,G65627);
  xor GNAME65640(G65640,G65641,G76648);
  xor GNAME65641(G65641,G75217,G76651);
  and GNAME65642(G65642,G75217,G76648);
  and GNAME65643(G65643,G76651,G76648);
  and GNAME65644(G65644,G75217,G76651);
  or GNAME65645(G65645,G65644,G65643,G65642);
  xor GNAME65655(G65655,G65656,G76654);
  xor GNAME65656(G65656,G75218,G76657);
  and GNAME65657(G65657,G75218,G76654);
  and GNAME65658(G65658,G76657,G76654);
  and GNAME65659(G65659,G75218,G76657);
  or GNAME65660(G65660,G65659,G65658,G65657);
  xor GNAME65670(G65670,G65671,G76660);
  xor GNAME65671(G65671,G75219,G76663);
  and GNAME65672(G65672,G75219,G76660);
  and GNAME65673(G65673,G76663,G76660);
  and GNAME65674(G65674,G75219,G76663);
  or GNAME65675(G65675,G65674,G65673,G65672);
  xor GNAME65685(G65685,G65686,G76669);
  xor GNAME65686(G65686,G77810,G76666);
  and GNAME65687(G65687,G77810,G76669);
  and GNAME65688(G65688,G76666,G76669);
  and GNAME65689(G65689,G77810,G76666);
  or GNAME65690(G65690,G65689,G65688,G65687);
  xor GNAME65700(G65700,G65701,G76675);
  xor GNAME65701(G65701,G77811,G76672);
  and GNAME65702(G65702,G77811,G76675);
  and GNAME65703(G65703,G76672,G76675);
  and GNAME65704(G65704,G77811,G76672);
  or GNAME65705(G65705,G65704,G65703,G65702);
  xor GNAME65715(G65715,G65716,G76681);
  xor GNAME65716(G65716,G77812,G76678);
  and GNAME65717(G65717,G77812,G76681);
  and GNAME65718(G65718,G76678,G76681);
  and GNAME65719(G65719,G77812,G76678);
  or GNAME65720(G65720,G65719,G65718,G65717);
  xor GNAME65730(G65730,G65731,G76690);
  xor GNAME65731(G65731,G76684,G76687);
  and GNAME65732(G65732,G76684,G76690);
  and GNAME65733(G65733,G76687,G76690);
  and GNAME65734(G65734,G76684,G76687);
  or GNAME65735(G65735,G65734,G65733,G65732);
  xor GNAME65745(G65745,G65746,G76699);
  xor GNAME65746(G65746,G76693,G76696);
  and GNAME65747(G65747,G76693,G76699);
  and GNAME65748(G65748,G76696,G76699);
  and GNAME65749(G65749,G76693,G76696);
  or GNAME65750(G65750,G65749,G65748,G65747);
  xor GNAME65760(G65760,G65761,G76708);
  xor GNAME65761(G65761,G76702,G76705);
  and GNAME65762(G65762,G76702,G76708);
  and GNAME65763(G65763,G76705,G76708);
  and GNAME65764(G65764,G76702,G76705);
  or GNAME65765(G65765,G65764,G65763,G65762);
  xor GNAME65775(G65775,G65776,G76717);
  xor GNAME65776(G65776,G76711,G76714);
  and GNAME65777(G65777,G76711,G76717);
  and GNAME65778(G65778,G76714,G76717);
  and GNAME65779(G65779,G76711,G76714);
  or GNAME65780(G65780,G65779,G65778,G65777);
  xor GNAME65790(G65790,G65791,G76726);
  xor GNAME65791(G65791,G76720,G76723);
  and GNAME65792(G65792,G76720,G76726);
  and GNAME65793(G65793,G76723,G76726);
  and GNAME65794(G65794,G76720,G76723);
  or GNAME65795(G65795,G65794,G65793,G65792);
  xor GNAME65805(G65805,G65806,G76735);
  xor GNAME65806(G65806,G76729,G76732);
  and GNAME65807(G65807,G76729,G76735);
  and GNAME65808(G65808,G76732,G76735);
  and GNAME65809(G65809,G76729,G76732);
  or GNAME65810(G65810,G65809,G65808,G65807);
  xor GNAME65820(G65820,G65821,G76744);
  xor GNAME65821(G65821,G76738,G76741);
  and GNAME65822(G65822,G76738,G76744);
  and GNAME65823(G65823,G76741,G76744);
  and GNAME65824(G65824,G76738,G76741);
  or GNAME65825(G65825,G65824,G65823,G65822);
  xor GNAME65835(G65835,G65836,G76753);
  xor GNAME65836(G65836,G76747,G76750);
  and GNAME65837(G65837,G76747,G76753);
  and GNAME65838(G65838,G76750,G76753);
  and GNAME65839(G65839,G76747,G76750);
  or GNAME65840(G65840,G65839,G65838,G65837);
  xor GNAME65850(G65850,G65851,G76762);
  xor GNAME65851(G65851,G76756,G76759);
  and GNAME65852(G65852,G76756,G76762);
  and GNAME65853(G65853,G76759,G76762);
  and GNAME65854(G65854,G76756,G76759);
  or GNAME65855(G65855,G65854,G65853,G65852);
  xor GNAME65865(G65865,G65866,G76771);
  xor GNAME65866(G65866,G76765,G76768);
  and GNAME65867(G65867,G76765,G76771);
  and GNAME65868(G65868,G76768,G76771);
  and GNAME65869(G65869,G76765,G76768);
  or GNAME65870(G65870,G65869,G65868,G65867);
  xor GNAME65880(G65880,G65881,G76780);
  xor GNAME65881(G65881,G76774,G76777);
  and GNAME65882(G65882,G76774,G76780);
  and GNAME65883(G65883,G76777,G76780);
  and GNAME65884(G65884,G76774,G76777);
  or GNAME65885(G65885,G65884,G65883,G65882);
  xor GNAME65895(G65895,G65896,G76789);
  xor GNAME65896(G65896,G76783,G76786);
  and GNAME65897(G65897,G76783,G76789);
  and GNAME65898(G65898,G76786,G76789);
  and GNAME65899(G65899,G76783,G76786);
  or GNAME65900(G65900,G65899,G65898,G65897);
  xor GNAME65910(G65910,G65911,G76792);
  xor GNAME65911(G65911,G75220,G76795);
  and GNAME65912(G65912,G75220,G76792);
  and GNAME65913(G65913,G76795,G76792);
  and GNAME65914(G65914,G75220,G76795);
  or GNAME65915(G65915,G65914,G65913,G65912);
  xor GNAME65925(G65925,G65926,G76798);
  xor GNAME65926(G65926,G75221,G76801);
  and GNAME65927(G65927,G75221,G76798);
  and GNAME65928(G65928,G76801,G76798);
  and GNAME65929(G65929,G75221,G76801);
  or GNAME65930(G65930,G65929,G65928,G65927);
  xor GNAME65940(G65940,G65941,G76804);
  xor GNAME65941(G65941,G75222,G76807);
  and GNAME65942(G65942,G75222,G76804);
  and GNAME65943(G65943,G76807,G76804);
  and GNAME65944(G65944,G75222,G76807);
  or GNAME65945(G65945,G65944,G65943,G65942);
  xor GNAME65955(G65955,G65956,G76810);
  xor GNAME65956(G65956,G75223,G76813);
  and GNAME65957(G65957,G75223,G76810);
  and GNAME65958(G65958,G76813,G76810);
  and GNAME65959(G65959,G75223,G76813);
  or GNAME65960(G65960,G65959,G65958,G65957);
  xor GNAME65970(G65970,G65971,G76816);
  xor GNAME65971(G65971,G75224,G76819);
  and GNAME65972(G65972,G75224,G76816);
  and GNAME65973(G65973,G76819,G76816);
  and GNAME65974(G65974,G75224,G76819);
  or GNAME65975(G65975,G65974,G65973,G65972);
  xor GNAME65985(G65985,G65986,G76822);
  xor GNAME65986(G65986,G75225,G76825);
  and GNAME65987(G65987,G75225,G76822);
  and GNAME65988(G65988,G76825,G76822);
  and GNAME65989(G65989,G75225,G76825);
  or GNAME65990(G65990,G65989,G65988,G65987);
  xor GNAME66000(G66000,G66001,G76834);
  xor GNAME66001(G66001,G76828,G76831);
  and GNAME66002(G66002,G76828,G76834);
  and GNAME66003(G66003,G76831,G76834);
  and GNAME66004(G66004,G76828,G76831);
  or GNAME66005(G66005,G66004,G66003,G66002);
  xor GNAME66015(G66015,G66016,G76843);
  xor GNAME66016(G66016,G76837,G76840);
  and GNAME66017(G66017,G76837,G76843);
  and GNAME66018(G66018,G76840,G76843);
  and GNAME66019(G66019,G76837,G76840);
  or GNAME66020(G66020,G66019,G66018,G66017);
  xor GNAME66030(G66030,G66031,G76852);
  xor GNAME66031(G66031,G76846,G76849);
  and GNAME66032(G66032,G76846,G76852);
  and GNAME66033(G66033,G76849,G76852);
  and GNAME66034(G66034,G76846,G76849);
  or GNAME66035(G66035,G66034,G66033,G66032);
  xor GNAME66045(G66045,G66046,G76861);
  xor GNAME66046(G66046,G76855,G76858);
  and GNAME66047(G66047,G76855,G76861);
  and GNAME66048(G66048,G76858,G76861);
  and GNAME66049(G66049,G76855,G76858);
  or GNAME66050(G66050,G66049,G66048,G66047);
  xor GNAME66060(G66060,G66061,G76870);
  xor GNAME66061(G66061,G76864,G76867);
  and GNAME66062(G66062,G76864,G76870);
  and GNAME66063(G66063,G76867,G76870);
  and GNAME66064(G66064,G76864,G76867);
  or GNAME66065(G66065,G66064,G66063,G66062);
  xor GNAME66075(G66075,G66076,G76879);
  xor GNAME66076(G66076,G76873,G76876);
  and GNAME66077(G66077,G76873,G76879);
  and GNAME66078(G66078,G76876,G76879);
  and GNAME66079(G66079,G76873,G76876);
  or GNAME66080(G66080,G66079,G66078,G66077);
  xor GNAME66090(G66090,G66091,G76888);
  xor GNAME66091(G66091,G76882,G76885);
  and GNAME66092(G66092,G76882,G76888);
  and GNAME66093(G66093,G76885,G76888);
  and GNAME66094(G66094,G76882,G76885);
  or GNAME66095(G66095,G66094,G66093,G66092);
  xor GNAME66105(G66105,G66106,G76897);
  xor GNAME66106(G66106,G76891,G76894);
  and GNAME66107(G66107,G76891,G76897);
  and GNAME66108(G66108,G76894,G76897);
  and GNAME66109(G66109,G76891,G76894);
  or GNAME66110(G66110,G66109,G66108,G66107);
  xor GNAME66120(G66120,G66121,G76906);
  xor GNAME66121(G66121,G76900,G76903);
  and GNAME66122(G66122,G76900,G76906);
  and GNAME66123(G66123,G76903,G76906);
  and GNAME66124(G66124,G76900,G76903);
  or GNAME66125(G66125,G66124,G66123,G66122);
  xor GNAME66135(G66135,G66136,G76915);
  xor GNAME66136(G66136,G76909,G76912);
  and GNAME66137(G66137,G76909,G76915);
  and GNAME66138(G66138,G76912,G76915);
  and GNAME66139(G66139,G76909,G76912);
  or GNAME66140(G66140,G66139,G66138,G66137);
  xor GNAME66150(G66150,G66151,G76924);
  xor GNAME66151(G66151,G76918,G76921);
  and GNAME66152(G66152,G76918,G76924);
  and GNAME66153(G66153,G76921,G76924);
  and GNAME66154(G66154,G76918,G76921);
  or GNAME66155(G66155,G66154,G66153,G66152);
  xor GNAME66165(G66165,G66166,G76933);
  xor GNAME66166(G66166,G76927,G76930);
  and GNAME66167(G66167,G76927,G76933);
  and GNAME66168(G66168,G76930,G76933);
  and GNAME66169(G66169,G76927,G76930);
  or GNAME66170(G66170,G66169,G66168,G66167);
  xor GNAME66180(G66180,G66181,G76936);
  xor GNAME66181(G66181,G75226,G76939);
  and GNAME66182(G66182,G75226,G76936);
  and GNAME66183(G66183,G76939,G76936);
  and GNAME66184(G66184,G75226,G76939);
  or GNAME66185(G66185,G66184,G66183,G66182);
  xor GNAME66195(G66195,G66196,G76942);
  xor GNAME66196(G66196,G75227,G76945);
  and GNAME66197(G66197,G75227,G76942);
  and GNAME66198(G66198,G76945,G76942);
  and GNAME66199(G66199,G75227,G76945);
  or GNAME66200(G66200,G66199,G66198,G66197);
  xor GNAME66210(G66210,G66211,G76948);
  xor GNAME66211(G66211,G75228,G76951);
  and GNAME66212(G66212,G75228,G76948);
  and GNAME66213(G66213,G76951,G76948);
  and GNAME66214(G66214,G75228,G76951);
  or GNAME66215(G66215,G66214,G66213,G66212);
  xor GNAME66225(G66225,G66226,G76954);
  xor GNAME66226(G66226,G75229,G76957);
  and GNAME66227(G66227,G75229,G76954);
  and GNAME66228(G66228,G76957,G76954);
  and GNAME66229(G66229,G75229,G76957);
  or GNAME66230(G66230,G66229,G66228,G66227);
  xor GNAME66240(G66240,G66241,G76960);
  xor GNAME66241(G66241,G75230,G76963);
  and GNAME66242(G66242,G75230,G76960);
  and GNAME66243(G66243,G76963,G76960);
  and GNAME66244(G66244,G75230,G76963);
  or GNAME66245(G66245,G66244,G66243,G66242);
  xor GNAME66255(G66255,G66256,G76966);
  xor GNAME66256(G66256,G75231,G76969);
  and GNAME66257(G66257,G75231,G76966);
  and GNAME66258(G66258,G76969,G76966);
  and GNAME66259(G66259,G75231,G76969);
  or GNAME66260(G66260,G66259,G66258,G66257);
  xor GNAME66270(G66270,G66271,G76978);
  xor GNAME66271(G66271,G76972,G76975);
  and GNAME66272(G66272,G76972,G76978);
  and GNAME66273(G66273,G76975,G76978);
  and GNAME66274(G66274,G76972,G76975);
  or GNAME66275(G66275,G66274,G66273,G66272);
  xor GNAME66285(G66285,G66286,G76987);
  xor GNAME66286(G66286,G76981,G76984);
  and GNAME66287(G66287,G76981,G76987);
  and GNAME66288(G66288,G76984,G76987);
  and GNAME66289(G66289,G76981,G76984);
  or GNAME66290(G66290,G66289,G66288,G66287);
  xor GNAME66300(G66300,G66301,G76996);
  xor GNAME66301(G66301,G76990,G76993);
  and GNAME66302(G66302,G76990,G76996);
  and GNAME66303(G66303,G76993,G76996);
  and GNAME66304(G66304,G76990,G76993);
  or GNAME66305(G66305,G66304,G66303,G66302);
  xor GNAME66315(G66315,G66316,G77005);
  xor GNAME66316(G66316,G76999,G77002);
  and GNAME66317(G66317,G76999,G77005);
  and GNAME66318(G66318,G77002,G77005);
  and GNAME66319(G66319,G76999,G77002);
  or GNAME66320(G66320,G66319,G66318,G66317);
  xor GNAME66330(G66330,G66331,G77014);
  xor GNAME66331(G66331,G77008,G77011);
  and GNAME66332(G66332,G77008,G77014);
  and GNAME66333(G66333,G77011,G77014);
  and GNAME66334(G66334,G77008,G77011);
  or GNAME66335(G66335,G66334,G66333,G66332);
  xor GNAME66345(G66345,G66346,G77023);
  xor GNAME66346(G66346,G77017,G77020);
  and GNAME66347(G66347,G77017,G77023);
  and GNAME66348(G66348,G77020,G77023);
  and GNAME66349(G66349,G77017,G77020);
  or GNAME66350(G66350,G66349,G66348,G66347);
  xor GNAME66360(G66360,G66361,G77032);
  xor GNAME66361(G66361,G77026,G77029);
  and GNAME66362(G66362,G77026,G77032);
  and GNAME66363(G66363,G77029,G77032);
  and GNAME66364(G66364,G77026,G77029);
  or GNAME66365(G66365,G66364,G66363,G66362);
  xor GNAME66375(G66375,G66376,G77041);
  xor GNAME66376(G66376,G77035,G77038);
  and GNAME66377(G66377,G77035,G77041);
  and GNAME66378(G66378,G77038,G77041);
  and GNAME66379(G66379,G77035,G77038);
  or GNAME66380(G66380,G66379,G66378,G66377);
  xor GNAME66390(G66390,G66391,G77050);
  xor GNAME66391(G66391,G77044,G77047);
  and GNAME66392(G66392,G77044,G77050);
  and GNAME66393(G66393,G77047,G77050);
  and GNAME66394(G66394,G77044,G77047);
  or GNAME66395(G66395,G66394,G66393,G66392);
  xor GNAME66405(G66405,G66406,G77059);
  xor GNAME66406(G66406,G77053,G77056);
  and GNAME66407(G66407,G77053,G77059);
  and GNAME66408(G66408,G77056,G77059);
  and GNAME66409(G66409,G77053,G77056);
  or GNAME66410(G66410,G66409,G66408,G66407);
  xor GNAME66420(G66420,G66421,G77068);
  xor GNAME66421(G66421,G77062,G77065);
  and GNAME66422(G66422,G77062,G77068);
  and GNAME66423(G66423,G77065,G77068);
  and GNAME66424(G66424,G77062,G77065);
  or GNAME66425(G66425,G66424,G66423,G66422);
  xor GNAME66435(G66435,G66436,G77077);
  xor GNAME66436(G66436,G77071,G77074);
  and GNAME66437(G66437,G77071,G77077);
  and GNAME66438(G66438,G77074,G77077);
  and GNAME66439(G66439,G77071,G77074);
  or GNAME66440(G66440,G66439,G66438,G66437);
  xor GNAME66450(G66450,G66451,G77080);
  xor GNAME66451(G66451,G75232,G77083);
  and GNAME66452(G66452,G75232,G77080);
  and GNAME66453(G66453,G77083,G77080);
  and GNAME66454(G66454,G75232,G77083);
  or GNAME66455(G66455,G66454,G66453,G66452);
  xor GNAME66465(G66465,G66466,G77086);
  xor GNAME66466(G66466,G75233,G77089);
  and GNAME66467(G66467,G75233,G77086);
  and GNAME66468(G66468,G77089,G77086);
  and GNAME66469(G66469,G75233,G77089);
  or GNAME66470(G66470,G66469,G66468,G66467);
  xor GNAME66480(G66480,G66481,G77092);
  xor GNAME66481(G66481,G75234,G77095);
  and GNAME66482(G66482,G75234,G77092);
  and GNAME66483(G66483,G77095,G77092);
  and GNAME66484(G66484,G75234,G77095);
  or GNAME66485(G66485,G66484,G66483,G66482);
  xor GNAME66495(G66495,G66496,G77098);
  xor GNAME66496(G66496,G75235,G77101);
  and GNAME66497(G66497,G75235,G77098);
  and GNAME66498(G66498,G77101,G77098);
  and GNAME66499(G66499,G75235,G77101);
  or GNAME66500(G66500,G66499,G66498,G66497);
  xor GNAME66510(G66510,G66511,G77104);
  xor GNAME66511(G66511,G75236,G77107);
  and GNAME66512(G66512,G75236,G77104);
  and GNAME66513(G66513,G77107,G77104);
  and GNAME66514(G66514,G75236,G77107);
  or GNAME66515(G66515,G66514,G66513,G66512);
  xor GNAME66525(G66525,G66526,G77110);
  xor GNAME66526(G66526,G75237,G77113);
  and GNAME66527(G66527,G75237,G77110);
  and GNAME66528(G66528,G77113,G77110);
  and GNAME66529(G66529,G75237,G77113);
  or GNAME66530(G66530,G66529,G66528,G66527);
  xor GNAME66540(G66540,G66541,G77122);
  xor GNAME66541(G66541,G77116,G77119);
  and GNAME66542(G66542,G77116,G77122);
  and GNAME66543(G66543,G77119,G77122);
  and GNAME66544(G66544,G77116,G77119);
  or GNAME66545(G66545,G66544,G66543,G66542);
  xor GNAME66555(G66555,G66556,G77131);
  xor GNAME66556(G66556,G77125,G77128);
  and GNAME66557(G66557,G77125,G77131);
  and GNAME66558(G66558,G77128,G77131);
  and GNAME66559(G66559,G77125,G77128);
  or GNAME66560(G66560,G66559,G66558,G66557);
  xor GNAME66570(G66570,G66571,G77140);
  xor GNAME66571(G66571,G77134,G77137);
  and GNAME66572(G66572,G77134,G77140);
  and GNAME66573(G66573,G77137,G77140);
  and GNAME66574(G66574,G77134,G77137);
  or GNAME66575(G66575,G66574,G66573,G66572);
  xor GNAME66585(G66585,G66586,G77149);
  xor GNAME66586(G66586,G77143,G77146);
  and GNAME66587(G66587,G77143,G77149);
  and GNAME66588(G66588,G77146,G77149);
  and GNAME66589(G66589,G77143,G77146);
  or GNAME66590(G66590,G66589,G66588,G66587);
  xor GNAME66600(G66600,G66601,G77158);
  xor GNAME66601(G66601,G77152,G77155);
  and GNAME66602(G66602,G77152,G77158);
  and GNAME66603(G66603,G77155,G77158);
  and GNAME66604(G66604,G77152,G77155);
  or GNAME66605(G66605,G66604,G66603,G66602);
  xor GNAME66615(G66615,G66616,G77167);
  xor GNAME66616(G66616,G77161,G77164);
  and GNAME66617(G66617,G77161,G77167);
  and GNAME66618(G66618,G77164,G77167);
  and GNAME66619(G66619,G77161,G77164);
  or GNAME66620(G66620,G66619,G66618,G66617);
  xor GNAME66630(G66630,G66631,G66695);
  xor GNAME66631(G66631,G63800,G66875);
  and GNAME66632(G66632,G63800,G66695);
  and GNAME66633(G66633,G66875,G66695);
  and GNAME66634(G66634,G63800,G66875);
  or GNAME66635(G66635,G66634,G66633,G66632);
  xor GNAME66645(G66645,G66646,G66740);
  xor GNAME66646(G66646,G63815,G66920);
  and GNAME66647(G66647,G63815,G66740);
  and GNAME66648(G66648,G66920,G66740);
  and GNAME66649(G66649,G63815,G66920);
  or GNAME66650(G66650,G66649,G66648,G66647);
  xor GNAME66660(G66660,G66661,G66755);
  xor GNAME66661(G66661,G63830,G66935);
  and GNAME66662(G66662,G63830,G66755);
  and GNAME66663(G66663,G66935,G66755);
  and GNAME66664(G66664,G63830,G66935);
  or GNAME66665(G66665,G66664,G66663,G66662);
  xor GNAME66675(G66675,G66676,G77176);
  xor GNAME66676(G66676,G77170,G77173);
  and GNAME66677(G66677,G77170,G77176);
  and GNAME66678(G66678,G77173,G77176);
  and GNAME66679(G66679,G77170,G77173);
  or GNAME66680(G66680,G66679,G66678,G66677);
  xor GNAME66690(G66690,G66691,G77185);
  xor GNAME66691(G66691,G77179,G77182);
  and GNAME66692(G66692,G77179,G77185);
  and GNAME66693(G66693,G77182,G77185);
  and GNAME66694(G66694,G77179,G77182);
  or GNAME66695(G66695,G66694,G66693,G66692);
  xor GNAME66705(G66705,G66706,G77194);
  xor GNAME66706(G66706,G77188,G77191);
  and GNAME66707(G66707,G77188,G77194);
  and GNAME66708(G66708,G77191,G77194);
  and GNAME66709(G66709,G77188,G77191);
  or GNAME66710(G66710,G66709,G66708,G66707);
  xor GNAME66720(G66720,G66721,G77203);
  xor GNAME66721(G66721,G77197,G77200);
  and GNAME66722(G66722,G77197,G77203);
  and GNAME66723(G66723,G77200,G77203);
  and GNAME66724(G66724,G77197,G77200);
  or GNAME66725(G66725,G66724,G66723,G66722);
  xor GNAME66735(G66735,G66736,G77212);
  xor GNAME66736(G66736,G77206,G77209);
  and GNAME66737(G66737,G77206,G77212);
  and GNAME66738(G66738,G77209,G77212);
  and GNAME66739(G66739,G77206,G77209);
  or GNAME66740(G66740,G66739,G66738,G66737);
  xor GNAME66750(G66750,G66751,G77221);
  xor GNAME66751(G66751,G77215,G77218);
  and GNAME66752(G66752,G77215,G77221);
  and GNAME66753(G66753,G77218,G77221);
  and GNAME66754(G66754,G77215,G77218);
  or GNAME66755(G66755,G66754,G66753,G66752);
  xor GNAME66765(G66765,G66766,G66870);
  xor GNAME66766(G66766,G63795,G66690);
  and GNAME66767(G66767,G63795,G66870);
  and GNAME66768(G66768,G66690,G66870);
  and GNAME66769(G66769,G63795,G66690);
  or GNAME66770(G66770,G66769,G66768,G66767);
  xor GNAME66780(G66780,G66781,G66915);
  xor GNAME66781(G66781,G63810,G66735);
  and GNAME66782(G66782,G63810,G66915);
  and GNAME66783(G66783,G66735,G66915);
  and GNAME66784(G66784,G63810,G66735);
  or GNAME66785(G66785,G66784,G66783,G66782);
  xor GNAME66795(G66795,G66796,G66930);
  xor GNAME66796(G66796,G63825,G66750);
  and GNAME66797(G66797,G63825,G66930);
  and GNAME66798(G66798,G66750,G66930);
  and GNAME66799(G66799,G63825,G66750);
  or GNAME66800(G66800,G66799,G66798,G66797);
  xor GNAME66810(G66810,G66811,G77224);
  xor GNAME66811(G66811,G75238,G77227);
  and GNAME66812(G66812,G75238,G77224);
  and GNAME66813(G66813,G77227,G77224);
  and GNAME66814(G66814,G75238,G77227);
  or GNAME66815(G66815,G66814,G66813,G66812);
  xor GNAME66825(G66825,G66826,G77230);
  xor GNAME66826(G66826,G75239,G77233);
  and GNAME66827(G66827,G75239,G77230);
  and GNAME66828(G66828,G77233,G77230);
  and GNAME66829(G66829,G75239,G77233);
  or GNAME66830(G66830,G66829,G66828,G66827);
  xor GNAME66840(G66840,G66841,G77236);
  xor GNAME66841(G66841,G75240,G77239);
  and GNAME66842(G66842,G75240,G77236);
  and GNAME66843(G66843,G77239,G77236);
  and GNAME66844(G66844,G75240,G77239);
  or GNAME66845(G66845,G66844,G66843,G66842);
  xor GNAME66855(G66855,G66856,G77248);
  xor GNAME66856(G66856,G77242,G77245);
  and GNAME66857(G66857,G77242,G77248);
  and GNAME66858(G66858,G77245,G77248);
  and GNAME66859(G66859,G77242,G77245);
  or GNAME66860(G66860,G66859,G66858,G66857);
  xor GNAME66870(G66870,G66871,G77257);
  xor GNAME66871(G66871,G77251,G77254);
  and GNAME66872(G66872,G77251,G77257);
  and GNAME66873(G66873,G77254,G77257);
  and GNAME66874(G66874,G77251,G77254);
  or GNAME66875(G66875,G66874,G66873,G66872);
  xor GNAME66885(G66885,G66886,G77266);
  xor GNAME66886(G66886,G77260,G77263);
  and GNAME66887(G66887,G77260,G77266);
  and GNAME66888(G66888,G77263,G77266);
  and GNAME66889(G66889,G77260,G77263);
  or GNAME66890(G66890,G66889,G66888,G66887);
  xor GNAME66900(G66900,G66901,G77275);
  xor GNAME66901(G66901,G77269,G77272);
  and GNAME66902(G66902,G77269,G77275);
  and GNAME66903(G66903,G77272,G77275);
  and GNAME66904(G66904,G77269,G77272);
  or GNAME66905(G66905,G66904,G66903,G66902);
  xor GNAME66915(G66915,G66916,G77284);
  xor GNAME66916(G66916,G77278,G77281);
  and GNAME66917(G66917,G77278,G77284);
  and GNAME66918(G66918,G77281,G77284);
  and GNAME66919(G66919,G77278,G77281);
  or GNAME66920(G66920,G66919,G66918,G66917);
  xor GNAME66930(G66930,G66931,G77293);
  xor GNAME66931(G66931,G77287,G77290);
  and GNAME66932(G66932,G77287,G77293);
  and GNAME66933(G66933,G77290,G77293);
  and GNAME66934(G66934,G77287,G77290);
  or GNAME66935(G66935,G66934,G66933,G66932);
  xor GNAME66945(G66945,G66946,G77302);
  xor GNAME66946(G66946,G77296,G77299);
  and GNAME66947(G66947,G77296,G77302);
  and GNAME66948(G66948,G77299,G77302);
  and GNAME66949(G66949,G77296,G77299);
  or GNAME66950(G66950,G66949,G66948,G66947);
  xor GNAME66960(G66960,G66961,G77311);
  xor GNAME66961(G66961,G77305,G77308);
  and GNAME66962(G66962,G77305,G77311);
  and GNAME66963(G66963,G77308,G77311);
  and GNAME66964(G66964,G77305,G77308);
  or GNAME66965(G66965,G66964,G66963,G66962);
  xor GNAME66975(G66975,G66976,G77320);
  xor GNAME66976(G66976,G77314,G77317);
  and GNAME66977(G66977,G77314,G77320);
  and GNAME66978(G66978,G77317,G77320);
  and GNAME66979(G66979,G77314,G77317);
  or GNAME66980(G66980,G66979,G66978,G66977);
  xor GNAME66990(G66990,G66991,G66950);
  xor GNAME66991(G66991,G74381,G67175);
  and GNAME66992(G66992,G74381,G66950);
  and GNAME66993(G66993,G67175,G66950);
  and GNAME66994(G66994,G74381,G67175);
  or GNAME66995(G66995,G66994,G66993,G66992);
  xor GNAME67005(G67005,G67006,G66965);
  xor GNAME67006(G67006,G74387,G67205);
  and GNAME67007(G67007,G74387,G66965);
  and GNAME67008(G67008,G67205,G66965);
  and GNAME67009(G67009,G74387,G67205);
  or GNAME67010(G67010,G67009,G67008,G67007);
  xor GNAME67020(G67020,G67021,G66980);
  xor GNAME67021(G67021,G74393,G67220);
  and GNAME67022(G67022,G74393,G66980);
  and GNAME67023(G67023,G67220,G66980);
  and GNAME67024(G67024,G74393,G67220);
  or GNAME67025(G67025,G67024,G67023,G67022);
  xor GNAME67035(G67035,G67036,G74363);
  xor GNAME67036(G67036,G77323,G77326);
  and GNAME67037(G67037,G77323,G74363);
  and GNAME67038(G67038,G77326,G74363);
  and GNAME67039(G67039,G77323,G77326);
  or GNAME67040(G67040,G67039,G67038,G67037);
  xor GNAME67050(G67050,G67051,G74369);
  xor GNAME67051(G67051,G77329,G77332);
  and GNAME67052(G67052,G77329,G74369);
  and GNAME67053(G67053,G77332,G74369);
  and GNAME67054(G67054,G77329,G77332);
  or GNAME67055(G67055,G67054,G67053,G67052);
  xor GNAME67065(G67065,G67066,G74375);
  xor GNAME67066(G67066,G77335,G77338);
  and GNAME67067(G67067,G77335,G74375);
  and GNAME67068(G67068,G77338,G74375);
  and GNAME67069(G67069,G77335,G77338);
  or GNAME67070(G67070,G67069,G67068,G67067);
  xor GNAME67080(G67080,G67081,G63845);
  xor GNAME67081(G67081,G77341,G74380);
  and GNAME67082(G67082,G77341,G63845);
  and GNAME67083(G67083,G74380,G63845);
  and GNAME67084(G67084,G77341,G74380);
  or GNAME67085(G67085,G67084,G67083,G67082);
  xor GNAME67095(G67095,G67096,G63860);
  xor GNAME67096(G67096,G77344,G74386);
  and GNAME67097(G67097,G77344,G63860);
  and GNAME67098(G67098,G74386,G63860);
  and GNAME67099(G67099,G77344,G74386);
  or GNAME67100(G67100,G67099,G67098,G67097);
  xor GNAME67110(G67110,G67111,G63875);
  xor GNAME67111(G67111,G77347,G74392);
  and GNAME67112(G67112,G77347,G63875);
  and GNAME67113(G67113,G74392,G63875);
  and GNAME67114(G67114,G77347,G74392);
  or GNAME67115(G67115,G67114,G67113,G67112);
  xor GNAME67125(G67125,G67126,G63840);
  xor GNAME67126(G67126,G67310,G67535);
  and GNAME67127(G67127,G67310,G63840);
  and GNAME67128(G67128,G67535,G63840);
  and GNAME67129(G67129,G67310,G67535);
  or GNAME67130(G67130,G67129,G67128,G67127);
  xor GNAME67140(G67140,G67141,G63855);
  xor GNAME67141(G67141,G67340,G67550);
  and GNAME67142(G67142,G67340,G63855);
  and GNAME67143(G67143,G67550,G63855);
  and GNAME67144(G67144,G67340,G67550);
  or GNAME67145(G67145,G67144,G67143,G67142);
  xor GNAME67155(G67155,G67156,G63870);
  xor GNAME67156(G67156,G67355,G67565);
  and GNAME67157(G67157,G67355,G63870);
  and GNAME67158(G67158,G67565,G63870);
  and GNAME67159(G67159,G67355,G67565);
  or GNAME67160(G67160,G67159,G67158,G67157);
  xor GNAME67170(G67170,G67171,G77353);
  xor GNAME67171(G67171,G77350,G77356);
  and GNAME67172(G67172,G77350,G77353);
  and GNAME67173(G67173,G77356,G77353);
  and GNAME67174(G67174,G77350,G77356);
  or GNAME67175(G67175,G67174,G67173,G67172);
  xor GNAME67185(G67185,G67186,G77365);
  xor GNAME67186(G67186,G77359,G77362);
  and GNAME67187(G67187,G77359,G77365);
  and GNAME67188(G67188,G77362,G77365);
  and GNAME67189(G67189,G77359,G77362);
  or GNAME67190(G67190,G67189,G67188,G67187);
  xor GNAME67200(G67200,G67201,G77371);
  xor GNAME67201(G67201,G77368,G77374);
  and GNAME67202(G67202,G77368,G77371);
  and GNAME67203(G67203,G77374,G77371);
  and GNAME67204(G67204,G77368,G77374);
  or GNAME67205(G67205,G67204,G67203,G67202);
  xor GNAME67215(G67215,G67216,G77380);
  xor GNAME67216(G67216,G77377,G77383);
  and GNAME67217(G67217,G77377,G77380);
  and GNAME67218(G67218,G77383,G77380);
  and GNAME67219(G67219,G77377,G77383);
  or GNAME67220(G67220,G67219,G67218,G67217);
  xor GNAME67230(G67230,G67231,G77392);
  xor GNAME67231(G67231,G77386,G77389);
  and GNAME67232(G67232,G77386,G77392);
  and GNAME67233(G67233,G77389,G77392);
  and GNAME67234(G67234,G77386,G77389);
  or GNAME67235(G67235,G67234,G67233,G67232);
  xor GNAME67245(G67245,G67246,G77401);
  xor GNAME67246(G67246,G77395,G77398);
  and GNAME67247(G67247,G77395,G77401);
  and GNAME67248(G67248,G77398,G77401);
  and GNAME67249(G67249,G77395,G77398);
  or GNAME67250(G67250,G67249,G67248,G67247);
  xor GNAME67260(G67260,G67261,G67460);
  xor GNAME67261(G67261,G63885,G67320);
  and GNAME67262(G67262,G63885,G67460);
  and GNAME67263(G67263,G67320,G67460);
  and GNAME67264(G67264,G63885,G67320);
  or GNAME67265(G67265,G67264,G67263,G67262);
  xor GNAME67275(G67275,G67276,G67505);
  xor GNAME67276(G67276,G63900,G67365);
  and GNAME67277(G67277,G63900,G67505);
  and GNAME67278(G67278,G67365,G67505);
  and GNAME67279(G67279,G63900,G67365);
  or GNAME67280(G67280,G67279,G67278,G67277);
  xor GNAME67290(G67290,G67291,G67520);
  xor GNAME67291(G67291,G63915,G67380);
  and GNAME67292(G67292,G63915,G67520);
  and GNAME67293(G67293,G67380,G67520);
  and GNAME67294(G67294,G63915,G67380);
  or GNAME67295(G67295,G67294,G67293,G67292);
  xor GNAME67305(G67305,G67306,G77410);
  xor GNAME67306(G67306,G77404,G77407);
  and GNAME67307(G67307,G77404,G77410);
  and GNAME67308(G67308,G77407,G77410);
  and GNAME67309(G67309,G77404,G77407);
  or GNAME67310(G67310,G67309,G67308,G67307);
  xor GNAME67320(G67320,G67321,G77419);
  xor GNAME67321(G67321,G77413,G77416);
  and GNAME67322(G67322,G77413,G77419);
  and GNAME67323(G67323,G77416,G77419);
  and GNAME67324(G67324,G77413,G77416);
  or GNAME67325(G67325,G67324,G67323,G67322);
  xor GNAME67335(G67335,G67336,G77428);
  xor GNAME67336(G67336,G77422,G77425);
  and GNAME67337(G67337,G77422,G77428);
  and GNAME67338(G67338,G77425,G77428);
  and GNAME67339(G67339,G77422,G77425);
  or GNAME67340(G67340,G67339,G67338,G67337);
  xor GNAME67350(G67350,G67351,G77437);
  xor GNAME67351(G67351,G77431,G77434);
  and GNAME67352(G67352,G77431,G77437);
  and GNAME67353(G67353,G77434,G77437);
  and GNAME67354(G67354,G77431,G77434);
  or GNAME67355(G67355,G67354,G67353,G67352);
  xor GNAME67365(G67365,G67366,G77446);
  xor GNAME67366(G67366,G77440,G77443);
  and GNAME67367(G67367,G77440,G77446);
  and GNAME67368(G67368,G77443,G77446);
  and GNAME67369(G67369,G77440,G77443);
  or GNAME67370(G67370,G67369,G67368,G67367);
  xor GNAME67380(G67380,G67381,G77455);
  xor GNAME67381(G67381,G77449,G77452);
  and GNAME67382(G67382,G77449,G77455);
  and GNAME67383(G67383,G77452,G77455);
  and GNAME67384(G67384,G77449,G77452);
  or GNAME67385(G67385,G67384,G67383,G67382);
  xor GNAME67395(G67395,G67396,G67325);
  xor GNAME67396(G67396,G74362,G63890);
  and GNAME67397(G67397,G74362,G67325);
  and GNAME67398(G67398,G63890,G67325);
  and GNAME67399(G67399,G74362,G63890);
  or GNAME67400(G67400,G67399,G67398,G67397);
  xor GNAME67410(G67410,G67411,G67370);
  xor GNAME67411(G67411,G74368,G63905);
  and GNAME67412(G67412,G74368,G67370);
  and GNAME67413(G67413,G63905,G67370);
  and GNAME67414(G67414,G74368,G63905);
  or GNAME67415(G67415,G67414,G67413,G67412);
  xor GNAME67425(G67425,G67426,G67385);
  xor GNAME67426(G67426,G74374,G63920);
  and GNAME67427(G67427,G74374,G67385);
  and GNAME67428(G67428,G63920,G67385);
  and GNAME67429(G67429,G74374,G63920);
  or GNAME67430(G67430,G67429,G67428,G67427);
  xor GNAME67440(G67440,G67441,G67580);
  xor GNAME67441(G67441,G77458,G74399);
  and GNAME67442(G67442,G77458,G67580);
  and GNAME67443(G67443,G74399,G67580);
  and GNAME67444(G67444,G77458,G74399);
  or GNAME67445(G67445,G67444,G67443,G67442);
  xor GNAME67455(G67455,G67456,G74398);
  xor GNAME67456(G67456,G77461,G77464);
  and GNAME67457(G67457,G77461,G74398);
  and GNAME67458(G67458,G77464,G74398);
  and GNAME67459(G67459,G77461,G77464);
  or GNAME67460(G67460,G67459,G67458,G67457);
  xor GNAME67470(G67470,G67471,G67595);
  xor GNAME67471(G67471,G77467,G74405);
  and GNAME67472(G67472,G77467,G67595);
  and GNAME67473(G67473,G74405,G67595);
  and GNAME67474(G67474,G77467,G74405);
  or GNAME67475(G67475,G67474,G67473,G67472);
  xor GNAME67485(G67485,G67486,G67610);
  xor GNAME67486(G67486,G77470,G74411);
  and GNAME67487(G67487,G77470,G67610);
  and GNAME67488(G67488,G74411,G67610);
  and GNAME67489(G67489,G77470,G74411);
  or GNAME67490(G67490,G67489,G67488,G67487);
  xor GNAME67500(G67500,G67501,G74404);
  xor GNAME67501(G67501,G77473,G77476);
  and GNAME67502(G67502,G77473,G74404);
  and GNAME67503(G67503,G77476,G74404);
  and GNAME67504(G67504,G77473,G77476);
  or GNAME67505(G67505,G67504,G67503,G67502);
  xor GNAME67515(G67515,G67516,G74410);
  xor GNAME67516(G67516,G77479,G77482);
  and GNAME67517(G67517,G77479,G74410);
  and GNAME67518(G67518,G77482,G74410);
  and GNAME67519(G67519,G77479,G77482);
  or GNAME67520(G67520,G67519,G67518,G67517);
  xor GNAME67530(G67530,G67531,G77488);
  xor GNAME67531(G67531,G77485,G77491);
  and GNAME67532(G67532,G77485,G77488);
  and GNAME67533(G67533,G77491,G77488);
  and GNAME67534(G67534,G77485,G77491);
  or GNAME67535(G67535,G67534,G67533,G67532);
  xor GNAME67545(G67545,G67546,G77497);
  xor GNAME67546(G67546,G77494,G77500);
  and GNAME67547(G67547,G77494,G77497);
  and GNAME67548(G67548,G77500,G77497);
  and GNAME67549(G67549,G77494,G77500);
  or GNAME67550(G67550,G67549,G67548,G67547);
  xor GNAME67560(G67560,G67561,G77506);
  xor GNAME67561(G67561,G77503,G77509);
  and GNAME67562(G67562,G77503,G77506);
  and GNAME67563(G67563,G77509,G77506);
  and GNAME67564(G67564,G77503,G77509);
  or GNAME67565(G67565,G67564,G67563,G67562);
  xor GNAME67575(G67575,G67576,G77515);
  xor GNAME67576(G67576,G77512,G77518);
  and GNAME67577(G67577,G77512,G77515);
  and GNAME67578(G67578,G77518,G77515);
  and GNAME67579(G67579,G77512,G77518);
  or GNAME67580(G67580,G67579,G67578,G67577);
  xor GNAME67590(G67590,G67591,G77524);
  xor GNAME67591(G67591,G77521,G77527);
  and GNAME67592(G67592,G77521,G77524);
  and GNAME67593(G67593,G77527,G77524);
  and GNAME67594(G67594,G77521,G77527);
  or GNAME67595(G67595,G67594,G67593,G67592);
  xor GNAME67605(G67605,G67606,G77533);
  xor GNAME67606(G67606,G77530,G77536);
  and GNAME67607(G67607,G77530,G77533);
  and GNAME67608(G67608,G77536,G77533);
  and GNAME67609(G67609,G77530,G77536);
  or GNAME67610(G67610,G67609,G67608,G67607);
  xor GNAME67620(G67620,G67621,G67575);
  xor GNAME67621(G67621,G63935,G67760);
  and GNAME67622(G67622,G63935,G67575);
  and GNAME67623(G67623,G67760,G67575);
  and GNAME67624(G67624,G63935,G67760);
  or GNAME67625(G67625,G67624,G67623,G67622);
  xor GNAME67635(G67635,G67636,G63930);
  xor GNAME67636(G67636,G74417,G67715);
  and GNAME67637(G67637,G74417,G63930);
  and GNAME67638(G67638,G67715,G63930);
  and GNAME67639(G67639,G74417,G67715);
  or GNAME67640(G67640,G67639,G67638,G67637);
  xor GNAME67650(G67650,G67651,G67590);
  xor GNAME67651(G67651,G63950,G67775);
  and GNAME67652(G67652,G63950,G67590);
  and GNAME67653(G67653,G67775,G67590);
  and GNAME67654(G67654,G63950,G67775);
  or GNAME67655(G67655,G67654,G67653,G67652);
  xor GNAME67665(G67665,G67666,G67605);
  xor GNAME67666(G67666,G63965,G67790);
  and GNAME67667(G67667,G63965,G67605);
  and GNAME67668(G67668,G67790,G67605);
  and GNAME67669(G67669,G63965,G67790);
  or GNAME67670(G67670,G67669,G67668,G67667);
  xor GNAME67680(G67680,G67681,G63945);
  xor GNAME67681(G67681,G74423,G67730);
  and GNAME67682(G67682,G74423,G63945);
  and GNAME67683(G67683,G67730,G63945);
  and GNAME67684(G67684,G74423,G67730);
  or GNAME67685(G67685,G67684,G67683,G67682);
  xor GNAME67695(G67695,G67696,G63960);
  xor GNAME67696(G67696,G74429,G67745);
  and GNAME67697(G67697,G74429,G63960);
  and GNAME67698(G67698,G67745,G63960);
  and GNAME67699(G67699,G74429,G67745);
  or GNAME67700(G67700,G67699,G67698,G67697);
  xor GNAME67710(G67710,G67711,G77542);
  xor GNAME67711(G67711,G77539,G77545);
  and GNAME67712(G67712,G77539,G77542);
  and GNAME67713(G67713,G77545,G77542);
  and GNAME67714(G67714,G77539,G77545);
  or GNAME67715(G67715,G67714,G67713,G67712);
  xor GNAME67725(G67725,G67726,G77551);
  xor GNAME67726(G67726,G77548,G77554);
  and GNAME67727(G67727,G77548,G77551);
  and GNAME67728(G67728,G77554,G77551);
  and GNAME67729(G67729,G77548,G77554);
  or GNAME67730(G67730,G67729,G67728,G67727);
  xor GNAME67740(G67740,G67741,G77560);
  xor GNAME67741(G67741,G77557,G77563);
  and GNAME67742(G67742,G77557,G77560);
  and GNAME67743(G67743,G77563,G77560);
  and GNAME67744(G67744,G77557,G77563);
  or GNAME67745(G67745,G67744,G67743,G67742);
  xor GNAME67755(G67755,G67756,G77572);
  xor GNAME67756(G67756,G77566,G77569);
  and GNAME67757(G67757,G77566,G77572);
  and GNAME67758(G67758,G77569,G77572);
  and GNAME67759(G67759,G77566,G77569);
  or GNAME67760(G67760,G67759,G67758,G67757);
  xor GNAME67770(G67770,G67771,G77581);
  xor GNAME67771(G67771,G77575,G77578);
  and GNAME67772(G67772,G77575,G77581);
  and GNAME67773(G67773,G77578,G77581);
  and GNAME67774(G67774,G77575,G77578);
  or GNAME67775(G67775,G67774,G67773,G67772);
  xor GNAME67785(G67785,G67786,G77590);
  xor GNAME67786(G67786,G77584,G77587);
  and GNAME67787(G67787,G77584,G77590);
  and GNAME67788(G67788,G77587,G77590);
  and GNAME67789(G67789,G77584,G77587);
  or GNAME67790(G67790,G67789,G67788,G67787);
  xor GNAME67800(G67800,G67801,G77596);
  xor GNAME67801(G67801,G77593,G77599);
  and GNAME67802(G67802,G77593,G77596);
  and GNAME67803(G67803,G77599,G77596);
  and GNAME67804(G67804,G77593,G77599);
  or GNAME67805(G67805,G67804,G67803,G67802);
  xor GNAME67815(G67815,G67816,G77605);
  xor GNAME67816(G67816,G77602,G77608);
  and GNAME67817(G67817,G77602,G77605);
  and GNAME67818(G67818,G77608,G77605);
  and GNAME67819(G67819,G77602,G77608);
  or GNAME67820(G67820,G67819,G67818,G67817);
  xor GNAME67830(G67830,G67831,G77614);
  xor GNAME67831(G67831,G77611,G77617);
  and GNAME67832(G67832,G77611,G77614);
  and GNAME67833(G67833,G77617,G77614);
  and GNAME67834(G67834,G77611,G77617);
  or GNAME67835(G67835,G67834,G67833,G67832);
  xor GNAME67845(G67845,G67846,G74435);
  xor GNAME67846(G67846,G77620,G77623);
  and GNAME67847(G67847,G77620,G74435);
  and GNAME67848(G67848,G77623,G74435);
  and GNAME67849(G67849,G77620,G77623);
  or GNAME67850(G67850,G67849,G67848,G67847);
  xor GNAME67860(G67860,G67861,G74441);
  xor GNAME67861(G67861,G77626,G77629);
  and GNAME67862(G67862,G77626,G74441);
  and GNAME67863(G67863,G77629,G74441);
  and GNAME67864(G67864,G77626,G77629);
  or GNAME67865(G67865,G67864,G67863,G67862);
  xor GNAME67875(G67875,G67876,G74447);
  xor GNAME67876(G67876,G77632,G77635);
  and GNAME67877(G67877,G77632,G74447);
  and GNAME67878(G67878,G77635,G74447);
  and GNAME67879(G67879,G77632,G77635);
  or GNAME67880(G67880,G67879,G67878,G67877);
  xor GNAME67890(G67890,G67891,G63980);
  xor GNAME67891(G67891,G77638,G74416);
  and GNAME67892(G67892,G77638,G63980);
  and GNAME67893(G67893,G74416,G63980);
  and GNAME67894(G67894,G77638,G74416);
  or GNAME67895(G67895,G67894,G67893,G67892);
  xor GNAME67905(G67905,G67906,G63995);
  xor GNAME67906(G67906,G77641,G74422);
  and GNAME67907(G67907,G77641,G63995);
  and GNAME67908(G67908,G74422,G63995);
  and GNAME67909(G67909,G77641,G74422);
  or GNAME67910(G67910,G67909,G67908,G67907);
  xor GNAME67920(G67920,G67921,G64010);
  xor GNAME67921(G67921,G77644,G74428);
  and GNAME67922(G67922,G77644,G64010);
  and GNAME67923(G67923,G74428,G64010);
  and GNAME67924(G67924,G77644,G74428);
  or GNAME67925(G67925,G67924,G67923,G67922);
  xor GNAME67935(G67935,G67936,G67800);
  xor GNAME67936(G67936,G74434,G64025);
  and GNAME67937(G67937,G74434,G67800);
  and GNAME67938(G67938,G64025,G67800);
  and GNAME67939(G67939,G74434,G64025);
  or GNAME67940(G67940,G67939,G67938,G67937);
  xor GNAME67950(G67950,G67951,G67845);
  xor GNAME67951(G67951,G67805,G63975);
  and GNAME67952(G67952,G67805,G67845);
  and GNAME67953(G67953,G63975,G67845);
  and GNAME67954(G67954,G67805,G63975);
  or GNAME67955(G67955,G67954,G67953,G67952);
  xor GNAME67965(G67965,G67966,G67860);
  xor GNAME67966(G67966,G67820,G63990);
  and GNAME67967(G67967,G67820,G67860);
  and GNAME67968(G67968,G63990,G67860);
  and GNAME67969(G67969,G67820,G63990);
  or GNAME67970(G67970,G67969,G67968,G67967);
  xor GNAME67980(G67980,G67981,G67875);
  xor GNAME67981(G67981,G67835,G64005);
  and GNAME67982(G67982,G67835,G67875);
  and GNAME67983(G67983,G64005,G67875);
  and GNAME67984(G67984,G67835,G64005);
  or GNAME67985(G67985,G67984,G67983,G67982);
  xor GNAME67995(G67995,G67996,G67815);
  xor GNAME67996(G67996,G74440,G64040);
  and GNAME67997(G67997,G74440,G67815);
  and GNAME67998(G67998,G64040,G67815);
  and GNAME67999(G67999,G74440,G64040);
  or GNAME68000(G68000,G67999,G67998,G67997);
  xor GNAME68010(G68010,G68011,G67830);
  xor GNAME68011(G68011,G74446,G64055);
  and GNAME68012(G68012,G74446,G67830);
  and GNAME68013(G68013,G64055,G67830);
  and GNAME68014(G68014,G74446,G64055);
  or GNAME68015(G68015,G68014,G68013,G68012);
  xor GNAME68025(G68025,G68026,G64020);
  xor GNAME68026(G68026,G77647,G74471);
  and GNAME68027(G68027,G77647,G64020);
  and GNAME68028(G68028,G74471,G64020);
  and GNAME68029(G68029,G77647,G74471);
  or GNAME68030(G68030,G68029,G68028,G68027);
  xor GNAME68040(G68040,G68041,G75133);
  xor GNAME68041(G68041,G68030,G67935);
  and GNAME68042(G68042,G68030,G75133);
  and GNAME68043(G68043,G67935,G75133);
  and GNAME68044(G68044,G68030,G67935);
  or GNAME68045(G68045,G68044,G68043,G68042);
  xor GNAME68055(G68055,G68056,G64035);
  xor GNAME68056(G68056,G77650,G74477);
  and GNAME68057(G68057,G77650,G64035);
  and GNAME68058(G68058,G74477,G64035);
  and GNAME68059(G68059,G77650,G74477);
  or GNAME68060(G68060,G68059,G68058,G68057);
  xor GNAME68070(G68070,G68071,G75153);
  xor GNAME68071(G68071,G68060,G67995);
  and GNAME68072(G68072,G68060,G75153);
  and GNAME68073(G68073,G67995,G75153);
  and GNAME68074(G68074,G68060,G67995);
  or GNAME68075(G68075,G68074,G68073,G68072);
  xor GNAME68085(G68085,G68086,G64050);
  xor GNAME68086(G68086,G77653,G74483);
  and GNAME68087(G68087,G77653,G64050);
  and GNAME68088(G68088,G74483,G64050);
  and GNAME68089(G68089,G77653,G74483);
  or GNAME68090(G68090,G68089,G68088,G68087);
  xor GNAME68100(G68100,G68101,G75173);
  xor GNAME68101(G68101,G68090,G68010);
  and GNAME68102(G68102,G68090,G75173);
  and GNAME68103(G68103,G68010,G75173);
  and GNAME68104(G68104,G68090,G68010);
  or GNAME68105(G68105,G68104,G68103,G68102);
  xor GNAME68115(G68115,G68116,G64565);
  xor GNAME68116(G68116,G64470,G64425);
  and GNAME68117(G68117,G64470,G64565);
  and GNAME68118(G68118,G64425,G64565);
  and GNAME68119(G68119,G64470,G64425);
  or GNAME68120(G68120,G68119,G68118,G68117);
  xor GNAME68130(G68130,G68131,G64580);
  xor GNAME68131(G68131,G64485,G64440);
  and GNAME68132(G68132,G64485,G64580);
  and GNAME68133(G68133,G64440,G64580);
  and GNAME68134(G68134,G64485,G64440);
  or GNAME68135(G68135,G68134,G68133,G68132);
  xor GNAME68145(G68145,G68146,G64595);
  xor GNAME68146(G68146,G64500,G64455);
  and GNAME68147(G68147,G64500,G64595);
  and GNAME68148(G68148,G64455,G64595);
  and GNAME68149(G68149,G64500,G64455);
  or GNAME68150(G68150,G68149,G68148,G68147);
  xor GNAME68160(G68160,G68161,G68210);
  xor GNAME68161(G68161,G64655,G64560);
  and GNAME68162(G68162,G64655,G68210);
  and GNAME68163(G68163,G64560,G68210);
  and GNAME68164(G68164,G64655,G64560);
  or GNAME68165(G68165,G68164,G68163,G68162);
  xor GNAME68175(G68175,G68176,G68225);
  xor GNAME68176(G68176,G64670,G64575);
  and GNAME68177(G68177,G64670,G68225);
  and GNAME68178(G68178,G64575,G68225);
  and GNAME68179(G68179,G64670,G64575);
  or GNAME68180(G68180,G68179,G68178,G68177);
  xor GNAME68190(G68190,G68191,G68240);
  xor GNAME68191(G68191,G64685,G64590);
  and GNAME68192(G68192,G64685,G68240);
  and GNAME68193(G68193,G64590,G68240);
  and GNAME68194(G68194,G64685,G64590);
  or GNAME68195(G68195,G68194,G68193,G68192);
  xor GNAME68205(G68205,G68206,G64835);
  xor GNAME68206(G68206,G64925,G64605);
  and GNAME68207(G68207,G64925,G64835);
  and GNAME68208(G68208,G64605,G64835);
  and GNAME68209(G68209,G64925,G64605);
  or GNAME68210(G68210,G68209,G68208,G68207);
  xor GNAME68220(G68220,G68221,G64850);
  xor GNAME68221(G68221,G64940,G64620);
  and GNAME68222(G68222,G64940,G64850);
  and GNAME68223(G68223,G64620,G64850);
  and GNAME68224(G68224,G64940,G64620);
  or GNAME68225(G68225,G68224,G68223,G68222);
  xor GNAME68235(G68235,G68236,G64865);
  xor GNAME68236(G68236,G64955,G64635);
  and GNAME68237(G68237,G64955,G64865);
  and GNAME68238(G68238,G64635,G64865);
  and GNAME68239(G68239,G64955,G64635);
  or GNAME68240(G68240,G68239,G68238,G68237);
  xor GNAME68250(G68250,G68251,G68205);
  xor GNAME68251(G68251,G64650,G64700);
  and GNAME68252(G68252,G64650,G68205);
  and GNAME68253(G68253,G64700,G68205);
  and GNAME68254(G68254,G64650,G64700);
  or GNAME68255(G68255,G68254,G68253,G68252);
  xor GNAME68265(G68265,G68266,G64695);
  xor GNAME68266(G68266,G64830,G68345);
  and GNAME68267(G68267,G64830,G64695);
  and GNAME68268(G68268,G68345,G64695);
  and GNAME68269(G68269,G64830,G68345);
  or GNAME68270(G68270,G68269,G68268,G68267);
  xor GNAME68280(G68280,G68281,G68220);
  xor GNAME68281(G68281,G64665,G64715);
  and GNAME68282(G68282,G64665,G68220);
  and GNAME68283(G68283,G64715,G68220);
  and GNAME68284(G68284,G64665,G64715);
  or GNAME68285(G68285,G68284,G68283,G68282);
  xor GNAME68295(G68295,G68296,G68235);
  xor GNAME68296(G68296,G64680,G64730);
  and GNAME68297(G68297,G64680,G68235);
  and GNAME68298(G68298,G64730,G68235);
  and GNAME68299(G68299,G64680,G64730);
  or GNAME68300(G68300,G68299,G68298,G68297);
  xor GNAME68310(G68310,G68311,G64710);
  xor GNAME68311(G68311,G64845,G68375);
  and GNAME68312(G68312,G64845,G64710);
  and GNAME68313(G68313,G68375,G64710);
  and GNAME68314(G68314,G64845,G68375);
  or GNAME68315(G68315,G68314,G68313,G68312);
  xor GNAME68325(G68325,G68326,G64725);
  xor GNAME68326(G68326,G64860,G68405);
  and GNAME68327(G68327,G64860,G64725);
  and GNAME68328(G68328,G68405,G64725);
  and GNAME68329(G68329,G64860,G68405);
  or GNAME68330(G68330,G68329,G68328,G68327);
  xor GNAME68340(G68340,G68341,G65105);
  xor GNAME68341(G68341,G64875,G65015);
  and GNAME68342(G68342,G64875,G65105);
  and GNAME68343(G68343,G65015,G65105);
  and GNAME68344(G68344,G64875,G65015);
  or GNAME68345(G68345,G68344,G68343,G68342);
  xor GNAME68355(G68355,G68356,G68525);
  xor GNAME68356(G68356,G65240,G65010);
  and GNAME68357(G68357,G65240,G68525);
  and GNAME68358(G68358,G65010,G68525);
  and GNAME68359(G68359,G65240,G65010);
  or GNAME68360(G68360,G68359,G68358,G68357);
  xor GNAME68370(G68370,G68371,G65120);
  xor GNAME68371(G68371,G64890,G65030);
  and GNAME68372(G68372,G64890,G65120);
  and GNAME68373(G68373,G65030,G65120);
  and GNAME68374(G68374,G64890,G65030);
  or GNAME68375(G68375,G68374,G68373,G68372);
  xor GNAME68385(G68385,G68386,G68540);
  xor GNAME68386(G68386,G65270,G65025);
  and GNAME68387(G68387,G65270,G68540);
  and GNAME68388(G68388,G65025,G68540);
  and GNAME68389(G68389,G65270,G65025);
  or GNAME68390(G68390,G68389,G68388,G68387);
  xor GNAME68400(G68400,G68401,G65135);
  xor GNAME68401(G68401,G64905,G65045);
  and GNAME68402(G68402,G64905,G65135);
  and GNAME68403(G68403,G65045,G65135);
  and GNAME68404(G68404,G64905,G65045);
  or GNAME68405(G68405,G68404,G68403,G68402);
  xor GNAME68415(G68415,G68416,G68555);
  xor GNAME68416(G68416,G65285,G65040);
  and GNAME68417(G68417,G65285,G68555);
  and GNAME68418(G68418,G65040,G68555);
  and GNAME68419(G68419,G65285,G65040);
  or GNAME68420(G68420,G68419,G68418,G68417);
  xor GNAME68430(G68430,G68431,G68340);
  xor GNAME68431(G68431,G64785,G68360);
  and GNAME68432(G68432,G64785,G68340);
  and GNAME68433(G68433,G68360,G68340);
  and GNAME68434(G68434,G64785,G68360);
  or GNAME68435(G68435,G68434,G68433,G68432);
  xor GNAME68445(G68445,G68446,G68355);
  xor GNAME68446(G68446,G65100,G68570);
  and GNAME68447(G68447,G65100,G68355);
  and GNAME68448(G68448,G68570,G68355);
  and GNAME68449(G68449,G65100,G68570);
  or GNAME68450(G68450,G68449,G68448,G68447);
  xor GNAME68460(G68460,G68461,G68370);
  xor GNAME68461(G68461,G64800,G68390);
  and GNAME68462(G68462,G64800,G68370);
  and GNAME68463(G68463,G68390,G68370);
  and GNAME68464(G68464,G64800,G68390);
  or GNAME68465(G68465,G68464,G68463,G68462);
  xor GNAME68475(G68475,G68476,G68400);
  xor GNAME68476(G68476,G64815,G68420);
  and GNAME68477(G68477,G64815,G68400);
  and GNAME68478(G68478,G68420,G68400);
  and GNAME68479(G68479,G64815,G68420);
  or GNAME68480(G68480,G68479,G68478,G68477);
  xor GNAME68490(G68490,G68491,G68385);
  xor GNAME68491(G68491,G65115,G68600);
  and GNAME68492(G68492,G65115,G68385);
  and GNAME68493(G68493,G68600,G68385);
  and GNAME68494(G68494,G65115,G68600);
  or GNAME68495(G68495,G68494,G68493,G68492);
  xor GNAME68505(G68505,G68506,G68415);
  xor GNAME68506(G68506,G65130,G68630);
  and GNAME68507(G68507,G65130,G68415);
  and GNAME68508(G68508,G68630,G68415);
  and GNAME68509(G68509,G65130,G68630);
  or GNAME68510(G68510,G68509,G68508,G68507);
  xor GNAME68520(G68520,G68521,G65145);
  xor GNAME68521(G68521,G65330,G65055);
  and GNAME68522(G68522,G65330,G65145);
  and GNAME68523(G68523,G65055,G65145);
  and GNAME68524(G68524,G65330,G65055);
  or GNAME68525(G68525,G68524,G68523,G68522);
  xor GNAME68535(G68535,G68536,G65160);
  xor GNAME68536(G68536,G65360,G65070);
  and GNAME68537(G68537,G65360,G65160);
  and GNAME68538(G68538,G65070,G65160);
  and GNAME68539(G68539,G65360,G65070);
  or GNAME68540(G68540,G68539,G68538,G68537);
  xor GNAME68550(G68550,G68551,G65175);
  xor GNAME68551(G68551,G65375,G65085);
  and GNAME68552(G68552,G65375,G65175);
  and GNAME68553(G68553,G65085,G65175);
  and GNAME68554(G68554,G65375,G65085);
  or GNAME68555(G68555,G68554,G68553,G68552);
  xor GNAME68565(G68565,G68566,G65420);
  xor GNAME68566(G68566,G65255,G65235);
  and GNAME68567(G68567,G65255,G65420);
  and GNAME68568(G68568,G65235,G65420);
  and GNAME68569(G68569,G65255,G65235);
  or GNAME68570(G68570,G68569,G68568,G68567);
  xor GNAME68580(G68580,G68581,G65435);
  xor GNAME68581(G68581,G68705,G65250);
  and GNAME68582(G68582,G68705,G65435);
  and GNAME68583(G68583,G65250,G65435);
  and GNAME68584(G68584,G68705,G65250);
  or GNAME68585(G68585,G68584,G68583,G68582);
  xor GNAME68595(G68595,G68596,G65450);
  xor GNAME68596(G68596,G65300,G65265);
  and GNAME68597(G68597,G65300,G65450);
  and GNAME68598(G68598,G65265,G65450);
  and GNAME68599(G68599,G65300,G65265);
  or GNAME68600(G68600,G68599,G68598,G68597);
  xor GNAME68610(G68610,G68611,G65465);
  xor GNAME68611(G68611,G68720,G65295);
  and GNAME68612(G68612,G68720,G65465);
  and GNAME68613(G68613,G65295,G65465);
  and GNAME68614(G68614,G68720,G65295);
  or GNAME68615(G68615,G68614,G68613,G68612);
  xor GNAME68625(G68625,G68626,G65480);
  xor GNAME68626(G68626,G65315,G65280);
  and GNAME68627(G68627,G65315,G65480);
  and GNAME68628(G68628,G65280,G65480);
  and GNAME68629(G68629,G65315,G65280);
  or GNAME68630(G68630,G68629,G68628,G68627);
  xor GNAME68640(G68640,G68641,G65495);
  xor GNAME68641(G68641,G68735,G65310);
  and GNAME68642(G68642,G68735,G65495);
  and GNAME68643(G68643,G65310,G65495);
  and GNAME68644(G68644,G68735,G65310);
  or GNAME68645(G68645,G68644,G68643,G68642);
  xor GNAME68655(G68655,G68656,G68580);
  xor GNAME68656(G68656,G65415,G70505);
  and GNAME68657(G68657,G65415,G68580);
  and GNAME68658(G68658,G70505,G68580);
  and GNAME68659(G68659,G65415,G70505);
  or GNAME68660(G68660,G68659,G68658,G68657);
  xor GNAME68670(G68670,G68671,G68610);
  xor GNAME68671(G68671,G65445,G70535);
  and GNAME68672(G68672,G65445,G68610);
  and GNAME68673(G68673,G70535,G68610);
  and GNAME68674(G68674,G65445,G70535);
  or GNAME68675(G68675,G68674,G68673,G68672);
  xor GNAME68685(G68685,G68686,G68640);
  xor GNAME68686(G68686,G65475,G70565);
  and GNAME68687(G68687,G65475,G68640);
  and GNAME68688(G68688,G70565,G68640);
  and GNAME68689(G68689,G65475,G70565);
  or GNAME68690(G68690,G68689,G68688,G68687);
  xor GNAME68700(G68700,G68701,G65555);
  xor GNAME68701(G68701,G65690,G65735);
  and GNAME68702(G68702,G65690,G65555);
  and GNAME68703(G68703,G65735,G65555);
  and GNAME68704(G68704,G65690,G65735);
  or GNAME68705(G68705,G68704,G68703,G68702);
  xor GNAME68715(G68715,G68716,G65570);
  xor GNAME68716(G68716,G65705,G65765);
  and GNAME68717(G68717,G65705,G65570);
  and GNAME68718(G68718,G65765,G65570);
  and GNAME68719(G68719,G65705,G65765);
  or GNAME68720(G68720,G68719,G68718,G68717);
  xor GNAME68730(G68730,G68731,G65585);
  xor GNAME68731(G68731,G65720,G65780);
  and GNAME68732(G68732,G65720,G65585);
  and GNAME68733(G68733,G65780,G65585);
  and GNAME68734(G68734,G65720,G65780);
  or GNAME68735(G68735,G68734,G68733,G68732);
  xor GNAME68745(G68745,G68746,G70500);
  xor GNAME68746(G68746,G65430,G70520);
  and GNAME68747(G68747,G65430,G70500);
  and GNAME68748(G68748,G70520,G70500);
  and GNAME68749(G68749,G65430,G70520);
  or GNAME68750(G68750,G68749,G68748,G68747);
  xor GNAME68760(G68760,G68761,G70530);
  xor GNAME68761(G68761,G65460,G70550);
  and GNAME68762(G68762,G65460,G70530);
  and GNAME68763(G68763,G70550,G70530);
  and GNAME68764(G68764,G65460,G70550);
  or GNAME68765(G68765,G68764,G68763,G68762);
  xor GNAME68775(G68775,G68776,G70560);
  xor GNAME68776(G68776,G65490,G70580);
  and GNAME68777(G68777,G65490,G70560);
  and GNAME68778(G68778,G70580,G70560);
  and GNAME68779(G68779,G65490,G70580);
  or GNAME68780(G68780,G68779,G68778,G68777);
  xor GNAME68790(G68790,G68791,G65600);
  xor GNAME68791(G68791,G65645,G65750);
  and GNAME68792(G68792,G65645,G65600);
  and GNAME68793(G68793,G65750,G65600);
  and GNAME68794(G68794,G65645,G65750);
  or GNAME68795(G68795,G68794,G68793,G68792);
  xor GNAME68805(G68805,G68806,G65615);
  xor GNAME68806(G68806,G65660,G65795);
  and GNAME68807(G68807,G65660,G65615);
  and GNAME68808(G68808,G65795,G65615);
  and GNAME68809(G68809,G65660,G65795);
  or GNAME68810(G68810,G68809,G68808,G68807);
  xor GNAME68820(G68820,G68821,G65630);
  xor GNAME68821(G68821,G65675,G65810);
  and GNAME68822(G68822,G65675,G65630);
  and GNAME68823(G68823,G65810,G65630);
  and GNAME68824(G68824,G65675,G65810);
  or GNAME68825(G68825,G68824,G68823,G68822);
  xor GNAME68835(G68835,G68836,G65730);
  xor GNAME68836(G68836,G65685,G65550);
  and GNAME68837(G68837,G65685,G65730);
  and GNAME68838(G68838,G65550,G65730);
  and GNAME68839(G68839,G65685,G65550);
  or GNAME68840(G68840,G68839,G68838,G68837);
  xor GNAME68850(G68850,G68851,G65745);
  xor GNAME68851(G68851,G65640,G65595);
  and GNAME68852(G68852,G65640,G65745);
  and GNAME68853(G68853,G65595,G65745);
  and GNAME68854(G68854,G65640,G65595);
  or GNAME68855(G68855,G68854,G68853,G68852);
  xor GNAME68865(G68865,G68866,G65760);
  xor GNAME68866(G68866,G65700,G65565);
  and GNAME68867(G68867,G65700,G65760);
  and GNAME68868(G68868,G65565,G65760);
  and GNAME68869(G68869,G65700,G65565);
  or GNAME68870(G68870,G68869,G68868,G68867);
  xor GNAME68880(G68880,G68881,G65790);
  xor GNAME68881(G68881,G65655,G65610);
  and GNAME68882(G68882,G65655,G65790);
  and GNAME68883(G68883,G65610,G65790);
  and GNAME68884(G68884,G65655,G65610);
  or GNAME68885(G68885,G68884,G68883,G68882);
  xor GNAME68895(G68895,G68896,G65775);
  xor GNAME68896(G68896,G65715,G65580);
  and GNAME68897(G68897,G65715,G65775);
  and GNAME68898(G68898,G65580,G65775);
  and GNAME68899(G68899,G65715,G65580);
  or GNAME68900(G68900,G68899,G68898,G68897);
  xor GNAME68910(G68910,G68911,G65805);
  xor GNAME68911(G68911,G65670,G65625);
  and GNAME68912(G68912,G65670,G65805);
  and GNAME68913(G68913,G65625,G65805);
  and GNAME68914(G68914,G65670,G65625);
  or GNAME68915(G68915,G68914,G68913,G68912);
  xor GNAME68925(G68925,G68926,G65825);
  xor GNAME68926(G68926,G65915,G66005);
  and GNAME68927(G68927,G65915,G65825);
  and GNAME68928(G68928,G66005,G65825);
  and GNAME68929(G68929,G65915,G66005);
  or GNAME68930(G68930,G68929,G68928,G68927);
  xor GNAME68940(G68940,G68941,G65840);
  xor GNAME68941(G68941,G65930,G66020);
  and GNAME68942(G68942,G65930,G65840);
  and GNAME68943(G68943,G66020,G65840);
  and GNAME68944(G68944,G65930,G66020);
  or GNAME68945(G68945,G68944,G68943,G68942);
  xor GNAME68955(G68955,G68956,G65855);
  xor GNAME68956(G68956,G65945,G66035);
  and GNAME68957(G68957,G65945,G65855);
  and GNAME68958(G68958,G66035,G65855);
  and GNAME68959(G68959,G65945,G66035);
  or GNAME68960(G68960,G68959,G68958,G68957);
  xor GNAME68970(G68970,G68971,G65870);
  xor GNAME68971(G68971,G65960,G66050);
  and GNAME68972(G68972,G65960,G65870);
  and GNAME68973(G68973,G66050,G65870);
  and GNAME68974(G68974,G65960,G66050);
  or GNAME68975(G68975,G68974,G68973,G68972);
  xor GNAME68985(G68985,G68986,G65885);
  xor GNAME68986(G68986,G65975,G66065);
  and GNAME68987(G68987,G65975,G65885);
  and GNAME68988(G68988,G66065,G65885);
  and GNAME68989(G68989,G65975,G66065);
  or GNAME68990(G68990,G68989,G68988,G68987);
  xor GNAME69000(G69000,G69001,G65900);
  xor GNAME69001(G69001,G65990,G66080);
  and GNAME69002(G69002,G65990,G65900);
  and GNAME69003(G69003,G66080,G65900);
  and GNAME69004(G69004,G65990,G66080);
  or GNAME69005(G69005,G69004,G69003,G69002);
  xor GNAME69015(G69015,G69016,G66000);
  xor GNAME69016(G69016,G65910,G65820);
  and GNAME69017(G69017,G65910,G66000);
  and GNAME69018(G69018,G65820,G66000);
  and GNAME69019(G69019,G65910,G65820);
  or GNAME69020(G69020,G69019,G69018,G69017);
  xor GNAME69030(G69030,G69031,G66015);
  xor GNAME69031(G69031,G65925,G65835);
  and GNAME69032(G69032,G65925,G66015);
  and GNAME69033(G69033,G65835,G66015);
  and GNAME69034(G69034,G65925,G65835);
  or GNAME69035(G69035,G69034,G69033,G69032);
  xor GNAME69045(G69045,G69046,G66030);
  xor GNAME69046(G69046,G65940,G65850);
  and GNAME69047(G69047,G65940,G66030);
  and GNAME69048(G69048,G65850,G66030);
  and GNAME69049(G69049,G65940,G65850);
  or GNAME69050(G69050,G69049,G69048,G69047);
  xor GNAME69060(G69060,G69061,G66060);
  xor GNAME69061(G69061,G65970,G65880);
  and GNAME69062(G69062,G65970,G66060);
  and GNAME69063(G69063,G65880,G66060);
  and GNAME69064(G69064,G65970,G65880);
  or GNAME69065(G69065,G69064,G69063,G69062);
  xor GNAME69075(G69075,G69076,G66045);
  xor GNAME69076(G69076,G65955,G65865);
  and GNAME69077(G69077,G65955,G66045);
  and GNAME69078(G69078,G65865,G66045);
  and GNAME69079(G69079,G65955,G65865);
  or GNAME69080(G69080,G69079,G69078,G69077);
  xor GNAME69090(G69090,G69091,G66075);
  xor GNAME69091(G69091,G65985,G65895);
  and GNAME69092(G69092,G65985,G66075);
  and GNAME69093(G69093,G65895,G66075);
  and GNAME69094(G69094,G65985,G65895);
  or GNAME69095(G69095,G69094,G69093,G69092);
  xor GNAME69105(G69105,G69106,G66095);
  xor GNAME69106(G69106,G66185,G66275);
  and GNAME69107(G69107,G66185,G66095);
  and GNAME69108(G69108,G66275,G66095);
  and GNAME69109(G69109,G66185,G66275);
  or GNAME69110(G69110,G69109,G69108,G69107);
  xor GNAME69120(G69120,G69121,G66110);
  xor GNAME69121(G69121,G66200,G66290);
  and GNAME69122(G69122,G66200,G66110);
  and GNAME69123(G69123,G66290,G66110);
  and GNAME69124(G69124,G66200,G66290);
  or GNAME69125(G69125,G69124,G69123,G69122);
  xor GNAME69135(G69135,G69136,G66125);
  xor GNAME69136(G69136,G66215,G66305);
  and GNAME69137(G69137,G66215,G66125);
  and GNAME69138(G69138,G66305,G66125);
  and GNAME69139(G69139,G66215,G66305);
  or GNAME69140(G69140,G69139,G69138,G69137);
  xor GNAME69150(G69150,G69151,G66140);
  xor GNAME69151(G69151,G66230,G66320);
  and GNAME69152(G69152,G66230,G66140);
  and GNAME69153(G69153,G66320,G66140);
  and GNAME69154(G69154,G66230,G66320);
  or GNAME69155(G69155,G69154,G69153,G69152);
  xor GNAME69165(G69165,G69166,G66155);
  xor GNAME69166(G69166,G66245,G66335);
  and GNAME69167(G69167,G66245,G66155);
  and GNAME69168(G69168,G66335,G66155);
  and GNAME69169(G69169,G66245,G66335);
  or GNAME69170(G69170,G69169,G69168,G69167);
  xor GNAME69180(G69180,G69181,G66170);
  xor GNAME69181(G69181,G66260,G66350);
  and GNAME69182(G69182,G66260,G66170);
  and GNAME69183(G69183,G66350,G66170);
  and GNAME69184(G69184,G66260,G66350);
  or GNAME69185(G69185,G69184,G69183,G69182);
  xor GNAME69195(G69195,G69196,G66270);
  xor GNAME69196(G69196,G66180,G66090);
  and GNAME69197(G69197,G66180,G66270);
  and GNAME69198(G69198,G66090,G66270);
  and GNAME69199(G69199,G66180,G66090);
  or GNAME69200(G69200,G69199,G69198,G69197);
  xor GNAME69210(G69210,G69211,G66285);
  xor GNAME69211(G69211,G66195,G66105);
  and GNAME69212(G69212,G66195,G66285);
  and GNAME69213(G69213,G66105,G66285);
  and GNAME69214(G69214,G66195,G66105);
  or GNAME69215(G69215,G69214,G69213,G69212);
  xor GNAME69225(G69225,G69226,G66300);
  xor GNAME69226(G69226,G66210,G66120);
  and GNAME69227(G69227,G66210,G66300);
  and GNAME69228(G69228,G66120,G66300);
  and GNAME69229(G69229,G66210,G66120);
  or GNAME69230(G69230,G69229,G69228,G69227);
  xor GNAME69240(G69240,G69241,G66330);
  xor GNAME69241(G69241,G66240,G66150);
  and GNAME69242(G69242,G66240,G66330);
  and GNAME69243(G69243,G66150,G66330);
  and GNAME69244(G69244,G66240,G66150);
  or GNAME69245(G69245,G69244,G69243,G69242);
  xor GNAME69255(G69255,G69256,G66315);
  xor GNAME69256(G69256,G66225,G66135);
  and GNAME69257(G69257,G66225,G66315);
  and GNAME69258(G69258,G66135,G66315);
  and GNAME69259(G69259,G66225,G66135);
  or GNAME69260(G69260,G69259,G69258,G69257);
  xor GNAME69270(G69270,G69271,G66345);
  xor GNAME69271(G69271,G66255,G66165);
  and GNAME69272(G69272,G66255,G66345);
  and GNAME69273(G69273,G66165,G66345);
  and GNAME69274(G69274,G66255,G66165);
  or GNAME69275(G69275,G69274,G69273,G69272);
  xor GNAME69285(G69285,G69286,G66365);
  xor GNAME69286(G69286,G66455,G66545);
  and GNAME69287(G69287,G66455,G66365);
  and GNAME69288(G69288,G66545,G66365);
  and GNAME69289(G69289,G66455,G66545);
  or GNAME69290(G69290,G69289,G69288,G69287);
  xor GNAME69300(G69300,G69301,G66380);
  xor GNAME69301(G69301,G66470,G66560);
  and GNAME69302(G69302,G66470,G66380);
  and GNAME69303(G69303,G66560,G66380);
  and GNAME69304(G69304,G66470,G66560);
  or GNAME69305(G69305,G69304,G69303,G69302);
  xor GNAME69315(G69315,G69316,G66395);
  xor GNAME69316(G69316,G66485,G66575);
  and GNAME69317(G69317,G66485,G66395);
  and GNAME69318(G69318,G66575,G66395);
  and GNAME69319(G69319,G66485,G66575);
  or GNAME69320(G69320,G69319,G69318,G69317);
  xor GNAME69330(G69330,G69331,G66410);
  xor GNAME69331(G69331,G66500,G66590);
  and GNAME69332(G69332,G66500,G66410);
  and GNAME69333(G69333,G66590,G66410);
  and GNAME69334(G69334,G66500,G66590);
  or GNAME69335(G69335,G69334,G69333,G69332);
  xor GNAME69345(G69345,G69346,G66425);
  xor GNAME69346(G69346,G66515,G66605);
  and GNAME69347(G69347,G66515,G66425);
  and GNAME69348(G69348,G66605,G66425);
  and GNAME69349(G69349,G66515,G66605);
  or GNAME69350(G69350,G69349,G69348,G69347);
  xor GNAME69360(G69360,G69361,G66440);
  xor GNAME69361(G69361,G66530,G66620);
  and GNAME69362(G69362,G66530,G66440);
  and GNAME69363(G69363,G66620,G66440);
  and GNAME69364(G69364,G66530,G66620);
  or GNAME69365(G69365,G69364,G69363,G69362);
  xor GNAME69375(G69375,G69376,G66540);
  xor GNAME69376(G69376,G66450,G66360);
  and GNAME69377(G69377,G66450,G66540);
  and GNAME69378(G69378,G66360,G66540);
  and GNAME69379(G69379,G66450,G66360);
  or GNAME69380(G69380,G69379,G69378,G69377);
  xor GNAME69390(G69390,G69391,G66555);
  xor GNAME69391(G69391,G66465,G66375);
  and GNAME69392(G69392,G66465,G66555);
  and GNAME69393(G69393,G66375,G66555);
  and GNAME69394(G69394,G66465,G66375);
  or GNAME69395(G69395,G69394,G69393,G69392);
  xor GNAME69405(G69405,G69406,G66570);
  xor GNAME69406(G69406,G66480,G66390);
  and GNAME69407(G69407,G66480,G66570);
  and GNAME69408(G69408,G66390,G66570);
  and GNAME69409(G69409,G66480,G66390);
  or GNAME69410(G69410,G69409,G69408,G69407);
  xor GNAME69420(G69420,G69421,G66600);
  xor GNAME69421(G69421,G66510,G66420);
  and GNAME69422(G69422,G66510,G66600);
  and GNAME69423(G69423,G66420,G66600);
  and GNAME69424(G69424,G66510,G66420);
  or GNAME69425(G69425,G69424,G69423,G69422);
  xor GNAME69435(G69435,G69436,G66585);
  xor GNAME69436(G69436,G66495,G66405);
  and GNAME69437(G69437,G66495,G66585);
  and GNAME69438(G69438,G66405,G66585);
  and GNAME69439(G69439,G66495,G66405);
  or GNAME69440(G69440,G69439,G69438,G69437);
  xor GNAME69450(G69450,G69451,G66615);
  xor GNAME69451(G69451,G66525,G66435);
  and GNAME69452(G69452,G66525,G66615);
  and GNAME69453(G69453,G66435,G66615);
  and GNAME69454(G69454,G66525,G66435);
  or GNAME69455(G69455,G69454,G69453,G69452);
  xor GNAME69465(G69465,G69466,G69605);
  xor GNAME69466(G69466,G66635,G69555);
  and GNAME69467(G69467,G66635,G69605);
  and GNAME69468(G69468,G69555,G69605);
  and GNAME69469(G69469,G66635,G69555);
  or GNAME69470(G69470,G69469,G69468,G69467);
  xor GNAME69480(G69480,G69481,G66770);
  xor GNAME69481(G69481,G66995,G66630);
  and GNAME69482(G69482,G66995,G66770);
  and GNAME69483(G69483,G66630,G66770);
  and GNAME69484(G69484,G66995,G66630);
  or GNAME69485(G69485,G69484,G69483,G69482);
  xor GNAME69495(G69495,G69496,G69620);
  xor GNAME69496(G69496,G66650,G69570);
  and GNAME69497(G69497,G66650,G69620);
  and GNAME69498(G69498,G69570,G69620);
  and GNAME69499(G69499,G66650,G69570);
  or GNAME69500(G69500,G69499,G69498,G69497);
  xor GNAME69510(G69510,G69511,G66785);
  xor GNAME69511(G69511,G67010,G66645);
  and GNAME69512(G69512,G67010,G66785);
  and GNAME69513(G69513,G66645,G66785);
  and GNAME69514(G69514,G67010,G66645);
  or GNAME69515(G69515,G69514,G69513,G69512);
  xor GNAME69525(G69525,G69526,G69635);
  xor GNAME69526(G69526,G66665,G69585);
  and GNAME69527(G69527,G66665,G69635);
  and GNAME69528(G69528,G69585,G69635);
  and GNAME69529(G69529,G66665,G69585);
  or GNAME69530(G69530,G69529,G69528,G69527);
  xor GNAME69540(G69540,G69541,G66800);
  xor GNAME69541(G69541,G67025,G66660);
  and GNAME69542(G69542,G67025,G66800);
  and GNAME69543(G69543,G66660,G66800);
  and GNAME69544(G69544,G67025,G66660);
  or GNAME69545(G69545,G69544,G69543,G69542);
  xor GNAME69555(G69555,G69556,G66680);
  xor GNAME69556(G69556,G66815,G66860);
  and GNAME69557(G69557,G66815,G66680);
  and GNAME69558(G69558,G66860,G66680);
  and GNAME69559(G69559,G66815,G66860);
  or GNAME69560(G69560,G69559,G69558,G69557);
  xor GNAME69570(G69570,G69571,G66710);
  xor GNAME69571(G69571,G66830,G66890);
  and GNAME69572(G69572,G66830,G66710);
  and GNAME69573(G69573,G66890,G66710);
  and GNAME69574(G69574,G66830,G66890);
  or GNAME69575(G69575,G69574,G69573,G69572);
  xor GNAME69585(G69585,G69586,G66725);
  xor GNAME69586(G69586,G66845,G66905);
  and GNAME69587(G69587,G66845,G66725);
  and GNAME69588(G69588,G66905,G66725);
  and GNAME69589(G69589,G66845,G66905);
  or GNAME69590(G69590,G69589,G69588,G69587);
  xor GNAME69600(G69600,G69601,G66855);
  xor GNAME69601(G69601,G66810,G66675);
  and GNAME69602(G69602,G66810,G66855);
  and GNAME69603(G69603,G66675,G66855);
  and GNAME69604(G69604,G66810,G66675);
  or GNAME69605(G69605,G69604,G69603,G69602);
  xor GNAME69615(G69615,G69616,G66885);
  xor GNAME69616(G69616,G66825,G66705);
  and GNAME69617(G69617,G66825,G66885);
  and GNAME69618(G69618,G66705,G66885);
  and GNAME69619(G69619,G66825,G66705);
  or GNAME69620(G69620,G69619,G69618,G69617);
  xor GNAME69630(G69630,G69631,G66900);
  xor GNAME69631(G69631,G66840,G66720);
  and GNAME69632(G69632,G66840,G66900);
  and GNAME69633(G69633,G66720,G66900);
  and GNAME69634(G69634,G66840,G66720);
  or GNAME69635(G69635,G69634,G69633,G69632);
  xor GNAME69645(G69645,G69646,G66990);
  xor GNAME69646(G69646,G67085,G69785);
  and GNAME69647(G69647,G67085,G66990);
  and GNAME69648(G69648,G69785,G66990);
  and GNAME69649(G69649,G67085,G69785);
  or GNAME69650(G69650,G69649,G69648,G69647);
  xor GNAME69660(G69660,G69661,G67130);
  xor GNAME69661(G69661,G67170,G67080);
  and GNAME69662(G69662,G67170,G67130);
  and GNAME69663(G69663,G67080,G67130);
  and GNAME69664(G69664,G67170,G67080);
  or GNAME69665(G69665,G69664,G69663,G69662);
  xor GNAME69675(G69675,G69676,G67005);
  xor GNAME69676(G69676,G67100,G69800);
  and GNAME69677(G69677,G67100,G67005);
  and GNAME69678(G69678,G69800,G67005);
  and GNAME69679(G69679,G67100,G69800);
  or GNAME69680(G69680,G69679,G69678,G69677);
  xor GNAME69690(G69690,G69691,G67145);
  xor GNAME69691(G69691,G67200,G67095);
  and GNAME69692(G69692,G67200,G67145);
  and GNAME69693(G69693,G67095,G67145);
  and GNAME69694(G69694,G67200,G67095);
  or GNAME69695(G69695,G69694,G69693,G69692);
  xor GNAME69705(G69705,G69706,G67020);
  xor GNAME69706(G69706,G67115,G69815);
  and GNAME69707(G69707,G67115,G67020);
  and GNAME69708(G69708,G69815,G67020);
  and GNAME69709(G69709,G67115,G69815);
  or GNAME69710(G69710,G69709,G69708,G69707);
  xor GNAME69720(G69720,G69721,G67160);
  xor GNAME69721(G69721,G67215,G67110);
  and GNAME69722(G69722,G67215,G67160);
  and GNAME69723(G69723,G67110,G67160);
  and GNAME69724(G69724,G67215,G67110);
  or GNAME69725(G69725,G69724,G69723,G69722);
  xor GNAME69735(G69735,G69736,G69645);
  xor GNAME69736(G69736,G66765,G69665);
  and GNAME69737(G69737,G66765,G69645);
  and GNAME69738(G69738,G69665,G69645);
  and GNAME69739(G69739,G66765,G69665);
  or GNAME69740(G69740,G69739,G69738,G69737);
  xor GNAME69750(G69750,G69751,G69675);
  xor GNAME69751(G69751,G66780,G69695);
  and GNAME69752(G69752,G66780,G69675);
  and GNAME69753(G69753,G69695,G69675);
  and GNAME69754(G69754,G66780,G69695);
  or GNAME69755(G69755,G69754,G69753,G69752);
  xor GNAME69765(G69765,G69766,G69705);
  xor GNAME69766(G69766,G66795,G69725);
  and GNAME69767(G69767,G66795,G69705);
  and GNAME69768(G69768,G69725,G69705);
  and GNAME69769(G69769,G66795,G69725);
  or GNAME69770(G69770,G69769,G69768,G69767);
  xor GNAME69780(G69780,G69781,G66945);
  xor GNAME69781(G69781,G67190,G67040);
  and GNAME69782(G69782,G67190,G66945);
  and GNAME69783(G69783,G67040,G66945);
  and GNAME69784(G69784,G67190,G67040);
  or GNAME69785(G69785,G69784,G69783,G69782);
  xor GNAME69795(G69795,G69796,G66960);
  xor GNAME69796(G69796,G67235,G67055);
  and GNAME69797(G69797,G67235,G66960);
  and GNAME69798(G69798,G67055,G66960);
  and GNAME69799(G69799,G67235,G67055);
  or GNAME69800(G69800,G69799,G69798,G69797);
  xor GNAME69810(G69810,G69811,G66975);
  xor GNAME69811(G69811,G67250,G67070);
  and GNAME69812(G69812,G67250,G66975);
  and GNAME69813(G69813,G67070,G66975);
  and GNAME69814(G69814,G67250,G67070);
  or GNAME69815(G69815,G69814,G69813,G69812);
  xor GNAME69825(G69825,G69826,G67400);
  xor GNAME69826(G69826,G67185,G67035);
  and GNAME69827(G69827,G67185,G67400);
  and GNAME69828(G69828,G67035,G67400);
  and GNAME69829(G69829,G67185,G67035);
  or GNAME69830(G69830,G69829,G69828,G69827);
  xor GNAME69840(G69840,G69841,G67445);
  xor GNAME69841(G69841,G67530,G67305);
  and GNAME69842(G69842,G67530,G67445);
  and GNAME69843(G69843,G67305,G67445);
  and GNAME69844(G69844,G67530,G67305);
  or GNAME69845(G69845,G69844,G69843,G69842);
  xor GNAME69855(G69855,G69856,G67415);
  xor GNAME69856(G69856,G67230,G67050);
  and GNAME69857(G69857,G67230,G67415);
  and GNAME69858(G69858,G67050,G67415);
  and GNAME69859(G69859,G67230,G67050);
  or GNAME69860(G69860,G69859,G69858,G69857);
  xor GNAME69870(G69870,G69871,G67475);
  xor GNAME69871(G69871,G67545,G67335);
  and GNAME69872(G69872,G67545,G67475);
  and GNAME69873(G69873,G67335,G67475);
  and GNAME69874(G69874,G67545,G67335);
  or GNAME69875(G69875,G69874,G69873,G69872);
  xor GNAME69885(G69885,G69886,G67430);
  xor GNAME69886(G69886,G67245,G67065);
  and GNAME69887(G69887,G67245,G67430);
  and GNAME69888(G69888,G67065,G67430);
  and GNAME69889(G69889,G67245,G67065);
  or GNAME69890(G69890,G69889,G69888,G69887);
  xor GNAME69900(G69900,G69901,G67490);
  xor GNAME69901(G69901,G67560,G67350);
  and GNAME69902(G69902,G67560,G67490);
  and GNAME69903(G69903,G67350,G67490);
  and GNAME69904(G69904,G67560,G67350);
  or GNAME69905(G69905,G69904,G69903,G69902);
  xor GNAME69915(G69915,G69916,G69825);
  xor GNAME69916(G69916,G67125,G69845);
  and GNAME69917(G69917,G67125,G69825);
  and GNAME69918(G69918,G69845,G69825);
  and GNAME69919(G69919,G67125,G69845);
  or GNAME69920(G69920,G69919,G69918,G69917);
  xor GNAME69930(G69930,G69931,G69840);
  xor GNAME69931(G69931,G67395,G67265);
  and GNAME69932(G69932,G67395,G69840);
  and GNAME69933(G69933,G67265,G69840);
  and GNAME69934(G69934,G67395,G67265);
  or GNAME69935(G69935,G69934,G69933,G69932);
  xor GNAME69945(G69945,G69946,G67260);
  xor GNAME69946(G69946,G67440,G67625);
  and GNAME69947(G69947,G67440,G67260);
  and GNAME69948(G69948,G67625,G67260);
  and GNAME69949(G69949,G67440,G67625);
  or GNAME69950(G69950,G69949,G69948,G69947);
  xor GNAME69960(G69960,G69961,G69855);
  xor GNAME69961(G69961,G67140,G69875);
  and GNAME69962(G69962,G67140,G69855);
  and GNAME69963(G69963,G69875,G69855);
  and GNAME69964(G69964,G67140,G69875);
  or GNAME69965(G69965,G69964,G69963,G69962);
  xor GNAME69975(G69975,G69976,G69885);
  xor GNAME69976(G69976,G67155,G69905);
  and GNAME69977(G69977,G67155,G69885);
  and GNAME69978(G69978,G69905,G69885);
  and GNAME69979(G69979,G67155,G69905);
  or GNAME69980(G69980,G69979,G69978,G69977);
  xor GNAME69990(G69990,G69991,G69870);
  xor GNAME69991(G69991,G67410,G67280);
  and GNAME69992(G69992,G67410,G69870);
  and GNAME69993(G69993,G67280,G69870);
  and GNAME69994(G69994,G67410,G67280);
  or GNAME69995(G69995,G69994,G69993,G69992);
  xor GNAME70005(G70005,G70006,G67275);
  xor GNAME70006(G70006,G67470,G67655);
  and GNAME70007(G70007,G67470,G67275);
  and GNAME70008(G70008,G67655,G67275);
  and GNAME70009(G70009,G67470,G67655);
  or GNAME70010(G70010,G70009,G70008,G70007);
  xor GNAME70020(G70020,G70021,G69900);
  xor GNAME70021(G70021,G67425,G67295);
  and GNAME70022(G70022,G67425,G69900);
  and GNAME70023(G70023,G67295,G69900);
  and GNAME70024(G70024,G67425,G67295);
  or GNAME70025(G70025,G70024,G70023,G70022);
  xor GNAME70035(G70035,G70036,G67290);
  xor GNAME70036(G70036,G67485,G67670);
  and GNAME70037(G70037,G67485,G67290);
  and GNAME70038(G70038,G67670,G67290);
  and GNAME70039(G70039,G67485,G67670);
  or GNAME70040(G70040,G70039,G70038,G70037);
  xor GNAME70050(G70050,G70051,G67620);
  xor GNAME70051(G70051,G67455,G67640);
  and GNAME70052(G70052,G67455,G67620);
  and GNAME70053(G70053,G67640,G67620);
  and GNAME70054(G70054,G67455,G67640);
  or GNAME70055(G70055,G70054,G70053,G70052);
  xor GNAME70065(G70065,G70066,G67635);
  xor GNAME70066(G70066,G67755,G67895);
  and GNAME70067(G70067,G67755,G67635);
  and GNAME70068(G70068,G67895,G67635);
  and GNAME70069(G70069,G67755,G67895);
  or GNAME70070(G70070,G70069,G70068,G70067);
  xor GNAME70080(G70080,G70081,G67650);
  xor GNAME70081(G70081,G67500,G67685);
  and GNAME70082(G70082,G67500,G67650);
  and GNAME70083(G70083,G67685,G67650);
  and GNAME70084(G70084,G67500,G67685);
  or GNAME70085(G70085,G70084,G70083,G70082);
  xor GNAME70095(G70095,G70096,G67680);
  xor GNAME70096(G70096,G67770,G67910);
  and GNAME70097(G70097,G67770,G67680);
  and GNAME70098(G70098,G67910,G67680);
  and GNAME70099(G70099,G67770,G67910);
  or GNAME70100(G70100,G70099,G70098,G70097);
  xor GNAME70110(G70110,G70111,G67665);
  xor GNAME70111(G70111,G67515,G67700);
  and GNAME70112(G70112,G67515,G67665);
  and GNAME70113(G70113,G67700,G67665);
  and GNAME70114(G70114,G67515,G67700);
  or GNAME70115(G70115,G70114,G70113,G70112);
  xor GNAME70125(G70125,G70126,G67695);
  xor GNAME70126(G70126,G67785,G67925);
  and GNAME70127(G70127,G67785,G67695);
  and GNAME70128(G70128,G67925,G67695);
  and GNAME70129(G70129,G67785,G67925);
  or GNAME70130(G70130,G70129,G70128,G70127);
  xor GNAME70140(G70140,G70141,G67890);
  xor GNAME70141(G70141,G67850,G67710);
  and GNAME70142(G70142,G67850,G67890);
  and GNAME70143(G70143,G67710,G67890);
  and GNAME70144(G70144,G67850,G67710);
  or GNAME70145(G70145,G70144,G70143,G70142);
  xor GNAME70155(G70155,G70156,G67905);
  xor GNAME70156(G70156,G67865,G67725);
  and GNAME70157(G70157,G67865,G67905);
  and GNAME70158(G70158,G67725,G67905);
  and GNAME70159(G70159,G67865,G67725);
  or GNAME70160(G70160,G70159,G70158,G70157);
  xor GNAME70170(G70170,G70171,G67920);
  xor GNAME70171(G70171,G67880,G67740);
  and GNAME70172(G70172,G67880,G67920);
  and GNAME70173(G70173,G67740,G67920);
  and GNAME70174(G70174,G67880,G67740);
  or GNAME70175(G70175,G70174,G70173,G70172);
  xor GNAME70185(G70185,G70186,G70205);
  xor GNAME70186(G70186,G64200,G64250);
  and GNAME70187(G70187,G64200,G70205);
  and GNAME70188(G70188,G64250,G70205);
  and GNAME70189(G70189,G64200,G64250);
  or GNAME70190(G70190,G70189,G70188,G70187);
  xor GNAME70200(G70200,G70201,G70220);
  xor GNAME70201(G70201,G64385,G64245);
  and GNAME70202(G70202,G64385,G70220);
  and GNAME70203(G70203,G64245,G70220);
  and GNAME70204(G70204,G64385,G64245);
  or GNAME70205(G70205,G70204,G70203,G70202);
  xor GNAME70215(G70215,G70216,G71315);
  xor GNAME70216(G70216,G68120,G64380);
  and GNAME70217(G70217,G68120,G71315);
  and GNAME70218(G70218,G64380,G71315);
  and GNAME70219(G70219,G68120,G64380);
  or GNAME70220(G70220,G70219,G70218,G70217);
  xor GNAME70230(G70230,G70231,G70265);
  xor GNAME70231(G70231,G64215,G64265);
  and GNAME70232(G70232,G64215,G70265);
  and GNAME70233(G70233,G64265,G70265);
  and GNAME70234(G70234,G64215,G64265);
  or GNAME70235(G70235,G70234,G70233,G70232);
  xor GNAME70245(G70245,G70246,G70295);
  xor GNAME70246(G70246,G64230,G64280);
  and GNAME70247(G70247,G64230,G70295);
  and GNAME70248(G70248,G64280,G70295);
  and GNAME70249(G70249,G64230,G64280);
  or GNAME70250(G70250,G70249,G70248,G70247);
  xor GNAME70260(G70260,G70261,G70280);
  xor GNAME70261(G70261,G64400,G64260);
  and GNAME70262(G70262,G64400,G70280);
  and GNAME70263(G70263,G64260,G70280);
  and GNAME70264(G70264,G64400,G64260);
  or GNAME70265(G70265,G70264,G70263,G70262);
  xor GNAME70275(G70275,G70276,G71450);
  xor GNAME70276(G70276,G68135,G64395);
  and GNAME70277(G70277,G68135,G71450);
  and GNAME70278(G70278,G64395,G71450);
  and GNAME70279(G70279,G68135,G64395);
  or GNAME70280(G70280,G70279,G70278,G70277);
  xor GNAME70290(G70290,G70291,G70310);
  xor GNAME70291(G70291,G64415,G64275);
  and GNAME70292(G70292,G64415,G70310);
  and GNAME70293(G70293,G64275,G70310);
  and GNAME70294(G70294,G64415,G64275);
  or GNAME70295(G70295,G70294,G70293,G70292);
  xor GNAME70305(G70305,G70306,G71480);
  xor GNAME70306(G70306,G68150,G64410);
  and GNAME70307(G70307,G68150,G71480);
  and GNAME70308(G70308,G64410,G71480);
  and GNAME70309(G70309,G68150,G64410);
  or GNAME70310(G70310,G70309,G70308,G70307);
  xor GNAME70320(G70320,G70321,G70340);
  xor GNAME70321(G70321,G67955,G70140);
  and GNAME70322(G70322,G67955,G70340);
  and GNAME70323(G70323,G70140,G70340);
  and GNAME70324(G70324,G67955,G70140);
  or GNAME70325(G70325,G70324,G70323,G70322);
  xor GNAME70335(G70335,G70336,G68045);
  xor GNAME70336(G70336,G67940,G67950);
  and GNAME70337(G70337,G67940,G68045);
  and GNAME70338(G70338,G67950,G68045);
  and GNAME70339(G70339,G67940,G67950);
  or GNAME70340(G70340,G70339,G70338,G70337);
  xor GNAME70350(G70350,G70351,G70385);
  xor GNAME70351(G70351,G67970,G70155);
  and GNAME70352(G70352,G67970,G70385);
  and GNAME70353(G70353,G70155,G70385);
  and GNAME70354(G70354,G67970,G70155);
  or GNAME70355(G70355,G70354,G70353,G70352);
  xor GNAME70365(G70365,G70366,G70400);
  xor GNAME70366(G70366,G67985,G70170);
  and GNAME70367(G70367,G67985,G70400);
  and GNAME70368(G70368,G70170,G70400);
  and GNAME70369(G70369,G67985,G70170);
  or GNAME70370(G70370,G70369,G70368,G70367);
  xor GNAME70380(G70380,G70381,G68075);
  xor GNAME70381(G70381,G68000,G67965);
  and GNAME70382(G70382,G68000,G68075);
  and GNAME70383(G70383,G67965,G68075);
  and GNAME70384(G70384,G68000,G67965);
  or GNAME70385(G70385,G70384,G70383,G70382);
  xor GNAME70395(G70395,G70396,G68105);
  xor GNAME70396(G70396,G68015,G67980);
  and GNAME70397(G70397,G68015,G68105);
  and GNAME70398(G70398,G67980,G68105);
  and GNAME70399(G70399,G68015,G67980);
  or GNAME70400(G70400,G70399,G70398,G70397);
  xor GNAME70410(G70410,G70411,G70190);
  xor GNAME70411(G70411,G64205,G64155);
  and GNAME70412(G70412,G64205,G70190);
  and GNAME70413(G70413,G64155,G70190);
  and GNAME70414(G70414,G64205,G64155);
  or GNAME70415(G70415,G70414,G70413,G70412);
  xor GNAME70425(G70425,G70426,G70235);
  xor GNAME70426(G70426,G64220,G64170);
  and GNAME70427(G70427,G64220,G70235);
  and GNAME70428(G70428,G64170,G70235);
  and GNAME70429(G70429,G64220,G64170);
  or GNAME70430(G70430,G70429,G70428,G70427);
  xor GNAME70440(G70440,G70441,G70250);
  xor GNAME70441(G70441,G64235,G64185);
  and GNAME70442(G70442,G64235,G70250);
  and GNAME70443(G70443,G64185,G70250);
  and GNAME70444(G70444,G64235,G64185);
  or GNAME70445(G70445,G70444,G70443,G70442);
  xor GNAME70455(G70455,G70456,G68565);
  xor GNAME70456(G70456,G68520,G68585);
  and GNAME70457(G70457,G68520,G68565);
  and GNAME70458(G70458,G68585,G68565);
  and GNAME70459(G70459,G68520,G68585);
  or GNAME70460(G70460,G70459,G70458,G70457);
  xor GNAME70470(G70470,G70471,G68595);
  xor GNAME70471(G70471,G68535,G68615);
  and GNAME70472(G70472,G68535,G68595);
  and GNAME70473(G70473,G68615,G68595);
  and GNAME70474(G70474,G68535,G68615);
  or GNAME70475(G70475,G70474,G70473,G70472);
  xor GNAME70485(G70485,G70486,G68625);
  xor GNAME70486(G70486,G68550,G68645);
  and GNAME70487(G70487,G68550,G68625);
  and GNAME70488(G70488,G68645,G68625);
  and GNAME70489(G70489,G68550,G68645);
  or GNAME70490(G70490,G70489,G70488,G70487);
  xor GNAME70500(G70500,G70501,G68700);
  xor GNAME70501(G70501,G68795,G68840);
  and GNAME70502(G70502,G68795,G68700);
  and GNAME70503(G70503,G68840,G68700);
  and GNAME70504(G70504,G68795,G68840);
  or GNAME70505(G70505,G70504,G70503,G70502);
  xor GNAME70515(G70515,G70516,G68855);
  xor GNAME70516(G70516,G68930,G68790);
  and GNAME70517(G70517,G68930,G68855);
  and GNAME70518(G70518,G68790,G68855);
  and GNAME70519(G70519,G68930,G68790);
  or GNAME70520(G70520,G70519,G70518,G70517);
  xor GNAME70530(G70530,G70531,G68715);
  xor GNAME70531(G70531,G68810,G68870);
  and GNAME70532(G70532,G68810,G68715);
  and GNAME70533(G70533,G68870,G68715);
  and GNAME70534(G70534,G68810,G68870);
  or GNAME70535(G70535,G70534,G70533,G70532);
  xor GNAME70545(G70545,G70546,G68885);
  xor GNAME70546(G70546,G68960,G68805);
  and GNAME70547(G70547,G68960,G68885);
  and GNAME70548(G70548,G68805,G68885);
  and GNAME70549(G70549,G68960,G68805);
  or GNAME70550(G70550,G70549,G70548,G70547);
  xor GNAME70560(G70560,G70561,G68730);
  xor GNAME70561(G70561,G68825,G68900);
  and GNAME70562(G70562,G68825,G68730);
  and GNAME70563(G70563,G68900,G68730);
  and GNAME70564(G70564,G68825,G68900);
  or GNAME70565(G70565,G70564,G70563,G70562);
  xor GNAME70575(G70575,G70576,G68915);
  xor GNAME70576(G70576,G68975,G68820);
  and GNAME70577(G70577,G68975,G68915);
  and GNAME70578(G70578,G68820,G68915);
  and GNAME70579(G70579,G68975,G68820);
  or GNAME70580(G70580,G70579,G70578,G70577);
  xor GNAME70590(G70590,G70591,G70515);
  xor GNAME70591(G70591,G68835,G70640);
  and GNAME70592(G70592,G68835,G70515);
  and GNAME70593(G70593,G70640,G70515);
  and GNAME70594(G70594,G68835,G70640);
  or GNAME70595(G70595,G70594,G70593,G70592);
  xor GNAME70605(G70605,G70606,G70545);
  xor GNAME70606(G70606,G68865,G70670);
  and GNAME70607(G70607,G68865,G70545);
  and GNAME70608(G70608,G70670,G70545);
  and GNAME70609(G70609,G68865,G70670);
  or GNAME70610(G70610,G70609,G70608,G70607);
  xor GNAME70620(G70620,G70621,G70575);
  xor GNAME70621(G70621,G68895,G70700);
  and GNAME70622(G70622,G68895,G70575);
  and GNAME70623(G70623,G70700,G70575);
  and GNAME70624(G70624,G68895,G70700);
  or GNAME70625(G70625,G70624,G70623,G70622);
  xor GNAME70635(G70635,G70636,G69020);
  xor GNAME70636(G70636,G68945,G68925);
  and GNAME70637(G70637,G68945,G69020);
  and GNAME70638(G70638,G68925,G69020);
  and GNAME70639(G70639,G68945,G68925);
  or GNAME70640(G70640,G70639,G70638,G70637);
  xor GNAME70650(G70650,G70651,G69035);
  xor GNAME70651(G70651,G69110,G68940);
  and GNAME70652(G70652,G69110,G69035);
  and GNAME70653(G70653,G68940,G69035);
  and GNAME70654(G70654,G69110,G68940);
  or GNAME70655(G70655,G70654,G70653,G70652);
  xor GNAME70665(G70665,G70666,G69050);
  xor GNAME70666(G70666,G68990,G68955);
  and GNAME70667(G70667,G68990,G69050);
  and GNAME70668(G70668,G68955,G69050);
  and GNAME70669(G70669,G68990,G68955);
  or GNAME70670(G70670,G70669,G70668,G70667);
  xor GNAME70680(G70680,G70681,G69065);
  xor GNAME70681(G70681,G69140,G68985);
  and GNAME70682(G70682,G69140,G69065);
  and GNAME70683(G70683,G68985,G69065);
  and GNAME70684(G70684,G69140,G68985);
  or GNAME70685(G70685,G70684,G70683,G70682);
  xor GNAME70695(G70695,G70696,G69080);
  xor GNAME70696(G70696,G69005,G68970);
  and GNAME70697(G70697,G69005,G69080);
  and GNAME70698(G70698,G68970,G69080);
  and GNAME70699(G70699,G69005,G68970);
  or GNAME70700(G70700,G70699,G70698,G70697);
  xor GNAME70710(G70710,G70711,G69095);
  xor GNAME70711(G70711,G69155,G69000);
  and GNAME70712(G70712,G69155,G69095);
  and GNAME70713(G70713,G69000,G69095);
  and GNAME70714(G70714,G69155,G69000);
  or GNAME70715(G70715,G70714,G70713,G70712);
  xor GNAME70725(G70725,G70726,G70635);
  xor GNAME70726(G70726,G68850,G70655);
  and GNAME70727(G70727,G68850,G70635);
  and GNAME70728(G70728,G70655,G70635);
  and GNAME70729(G70729,G68850,G70655);
  or GNAME70730(G70730,G70729,G70728,G70727);
  xor GNAME70740(G70740,G70741,G70650);
  xor GNAME70741(G70741,G69015,G70820);
  and GNAME70742(G70742,G69015,G70650);
  and GNAME70743(G70743,G70820,G70650);
  and GNAME70744(G70744,G69015,G70820);
  or GNAME70745(G70745,G70744,G70743,G70742);
  xor GNAME70755(G70755,G70756,G70665);
  xor GNAME70756(G70756,G68880,G70685);
  and GNAME70757(G70757,G68880,G70665);
  and GNAME70758(G70758,G70685,G70665);
  and GNAME70759(G70759,G68880,G70685);
  or GNAME70760(G70760,G70759,G70758,G70757);
  xor GNAME70770(G70770,G70771,G70695);
  xor GNAME70771(G70771,G68910,G70715);
  and GNAME70772(G70772,G68910,G70695);
  and GNAME70773(G70773,G70715,G70695);
  and GNAME70774(G70774,G68910,G70715);
  or GNAME70775(G70775,G70774,G70773,G70772);
  xor GNAME70785(G70785,G70786,G70680);
  xor GNAME70786(G70786,G69045,G70850);
  and GNAME70787(G70787,G69045,G70680);
  and GNAME70788(G70788,G70850,G70680);
  and GNAME70789(G70789,G69045,G70850);
  or GNAME70790(G70790,G70789,G70788,G70787);
  xor GNAME70800(G70800,G70801,G70710);
  xor GNAME70801(G70801,G69075,G70880);
  and GNAME70802(G70802,G69075,G70710);
  and GNAME70803(G70803,G70880,G70710);
  and GNAME70804(G70804,G69075,G70880);
  or GNAME70805(G70805,G70804,G70803,G70802);
  xor GNAME70815(G70815,G70816,G69200);
  xor GNAME70816(G70816,G69125,G69105);
  and GNAME70817(G70817,G69125,G69200);
  and GNAME70818(G70818,G69105,G69200);
  and GNAME70819(G70819,G69125,G69105);
  or GNAME70820(G70820,G70819,G70818,G70817);
  xor GNAME70830(G70830,G70831,G69215);
  xor GNAME70831(G70831,G69290,G69120);
  and GNAME70832(G70832,G69290,G69215);
  and GNAME70833(G70833,G69120,G69215);
  and GNAME70834(G70834,G69290,G69120);
  or GNAME70835(G70835,G70834,G70833,G70832);
  xor GNAME70845(G70845,G70846,G69230);
  xor GNAME70846(G70846,G69170,G69135);
  and GNAME70847(G70847,G69170,G69230);
  and GNAME70848(G70848,G69135,G69230);
  and GNAME70849(G70849,G69170,G69135);
  or GNAME70850(G70850,G70849,G70848,G70847);
  xor GNAME70860(G70860,G70861,G69245);
  xor GNAME70861(G70861,G69320,G69165);
  and GNAME70862(G70862,G69320,G69245);
  and GNAME70863(G70863,G69165,G69245);
  and GNAME70864(G70864,G69320,G69165);
  or GNAME70865(G70865,G70864,G70863,G70862);
  xor GNAME70875(G70875,G70876,G69260);
  xor GNAME70876(G70876,G69185,G69150);
  and GNAME70877(G70877,G69185,G69260);
  and GNAME70878(G70878,G69150,G69260);
  and GNAME70879(G70879,G69185,G69150);
  or GNAME70880(G70880,G70879,G70878,G70877);
  xor GNAME70890(G70890,G70891,G69275);
  xor GNAME70891(G70891,G69335,G69180);
  and GNAME70892(G70892,G69335,G69275);
  and GNAME70893(G70893,G69180,G69275);
  and GNAME70894(G70894,G69335,G69180);
  or GNAME70895(G70895,G70894,G70893,G70892);
  xor GNAME70905(G70905,G70906,G70815);
  xor GNAME70906(G70906,G69030,G70835);
  and GNAME70907(G70907,G69030,G70815);
  and GNAME70908(G70908,G70835,G70815);
  and GNAME70909(G70909,G69030,G70835);
  or GNAME70910(G70910,G70909,G70908,G70907);
  xor GNAME70920(G70920,G70921,G70830);
  xor GNAME70921(G70921,G69195,G71000);
  and GNAME70922(G70922,G69195,G70830);
  and GNAME70923(G70923,G71000,G70830);
  and GNAME70924(G70924,G69195,G71000);
  or GNAME70925(G70925,G70924,G70923,G70922);
  xor GNAME70935(G70935,G70936,G70845);
  xor GNAME70936(G70936,G69060,G70865);
  and GNAME70937(G70937,G69060,G70845);
  and GNAME70938(G70938,G70865,G70845);
  and GNAME70939(G70939,G69060,G70865);
  or GNAME70940(G70940,G70939,G70938,G70937);
  xor GNAME70950(G70950,G70951,G70875);
  xor GNAME70951(G70951,G69090,G70895);
  and GNAME70952(G70952,G69090,G70875);
  and GNAME70953(G70953,G70895,G70875);
  and GNAME70954(G70954,G69090,G70895);
  or GNAME70955(G70955,G70954,G70953,G70952);
  xor GNAME70965(G70965,G70966,G70860);
  xor GNAME70966(G70966,G69225,G71030);
  and GNAME70967(G70967,G69225,G70860);
  and GNAME70968(G70968,G71030,G70860);
  and GNAME70969(G70969,G69225,G71030);
  or GNAME70970(G70970,G70969,G70968,G70967);
  xor GNAME70980(G70980,G70981,G70890);
  xor GNAME70981(G70981,G69255,G71060);
  and GNAME70982(G70982,G69255,G70890);
  and GNAME70983(G70983,G71060,G70890);
  and GNAME70984(G70984,G69255,G71060);
  or GNAME70985(G70985,G70984,G70983,G70982);
  xor GNAME70995(G70995,G70996,G69380);
  xor GNAME70996(G70996,G69305,G69285);
  and GNAME70997(G70997,G69305,G69380);
  and GNAME70998(G70998,G69285,G69380);
  and GNAME70999(G70999,G69305,G69285);
  or GNAME71000(G71000,G70999,G70998,G70997);
  xor GNAME71010(G71010,G71011,G69395);
  xor GNAME71011(G71011,G69560,G69300);
  and GNAME71012(G71012,G69560,G69395);
  and GNAME71013(G71013,G69300,G69395);
  and GNAME71014(G71014,G69560,G69300);
  or GNAME71015(G71015,G71014,G71013,G71012);
  xor GNAME71025(G71025,G71026,G69410);
  xor GNAME71026(G71026,G69350,G69315);
  and GNAME71027(G71027,G69350,G69410);
  and GNAME71028(G71028,G69315,G69410);
  and GNAME71029(G71029,G69350,G69315);
  or GNAME71030(G71030,G71029,G71028,G71027);
  xor GNAME71040(G71040,G71041,G69425);
  xor GNAME71041(G71041,G69575,G69345);
  and GNAME71042(G71042,G69575,G69425);
  and GNAME71043(G71043,G69345,G69425);
  and GNAME71044(G71044,G69575,G69345);
  or GNAME71045(G71045,G71044,G71043,G71042);
  xor GNAME71055(G71055,G71056,G69440);
  xor GNAME71056(G71056,G69365,G69330);
  and GNAME71057(G71057,G69365,G69440);
  and GNAME71058(G71058,G69330,G69440);
  and GNAME71059(G71059,G69365,G69330);
  or GNAME71060(G71060,G71059,G71058,G71057);
  xor GNAME71070(G71070,G71071,G69455);
  xor GNAME71071(G71071,G69590,G69360);
  and GNAME71072(G71072,G69590,G69455);
  and GNAME71073(G71073,G69360,G69455);
  and GNAME71074(G71074,G69590,G69360);
  or GNAME71075(G71075,G71074,G71073,G71072);
  xor GNAME71085(G71085,G71086,G70995);
  xor GNAME71086(G71086,G69210,G71015);
  and GNAME71087(G71087,G69210,G70995);
  and GNAME71088(G71088,G71015,G70995);
  and GNAME71089(G71089,G69210,G71015);
  or GNAME71090(G71090,G71089,G71088,G71087);
  xor GNAME71100(G71100,G71101,G71010);
  xor GNAME71101(G71101,G69375,G69470);
  and GNAME71102(G71102,G69375,G71010);
  and GNAME71103(G71103,G69470,G71010);
  and GNAME71104(G71104,G69375,G69470);
  or GNAME71105(G71105,G71104,G71103,G71102);
  xor GNAME71115(G71115,G71116,G71025);
  xor GNAME71116(G71116,G69240,G71045);
  and GNAME71117(G71117,G69240,G71025);
  and GNAME71118(G71118,G71045,G71025);
  and GNAME71119(G71119,G69240,G71045);
  or GNAME71120(G71120,G71119,G71118,G71117);
  xor GNAME71130(G71130,G71131,G71055);
  xor GNAME71131(G71131,G69270,G71075);
  and GNAME71132(G71132,G69270,G71055);
  and GNAME71133(G71133,G71075,G71055);
  and GNAME71134(G71134,G69270,G71075);
  or GNAME71135(G71135,G71134,G71133,G71132);
  xor GNAME71145(G71145,G71146,G71040);
  xor GNAME71146(G71146,G69405,G69500);
  and GNAME71147(G71147,G69405,G71040);
  and GNAME71148(G71148,G69500,G71040);
  and GNAME71149(G71149,G69405,G69500);
  or GNAME71150(G71150,G71149,G71148,G71147);
  xor GNAME71160(G71160,G71161,G71070);
  xor GNAME71161(G71161,G69435,G69530);
  and GNAME71162(G71162,G69435,G71070);
  and GNAME71163(G71163,G69530,G71070);
  and GNAME71164(G71164,G69435,G69530);
  or GNAME71165(G71165,G71164,G71163,G71162);
  xor GNAME71175(G71175,G71176,G69465);
  xor GNAME71176(G71176,G69390,G69485);
  and GNAME71177(G71177,G69390,G69465);
  and GNAME71178(G71178,G69485,G69465);
  and GNAME71179(G71179,G69390,G69485);
  or GNAME71180(G71180,G71179,G71178,G71177);
  xor GNAME71190(G71190,G71191,G69480);
  xor GNAME71191(G71191,G69600,G69650);
  and GNAME71192(G71192,G69600,G69480);
  and GNAME71193(G71193,G69650,G69480);
  and GNAME71194(G71194,G69600,G69650);
  or GNAME71195(G71195,G71194,G71193,G71192);
  xor GNAME71205(G71205,G71206,G69495);
  xor GNAME71206(G71206,G69420,G69515);
  and GNAME71207(G71207,G69420,G69495);
  and GNAME71208(G71208,G69515,G69495);
  and GNAME71209(G71209,G69420,G69515);
  or GNAME71210(G71210,G71209,G71208,G71207);
  xor GNAME71220(G71220,G71221,G69525);
  xor GNAME71221(G71221,G69450,G69545);
  and GNAME71222(G71222,G69450,G69525);
  and GNAME71223(G71223,G69545,G69525);
  and GNAME71224(G71224,G69450,G69545);
  or GNAME71225(G71225,G71224,G71223,G71222);
  xor GNAME71235(G71235,G71236,G69510);
  xor GNAME71236(G71236,G69615,G69680);
  and GNAME71237(G71237,G69615,G69510);
  and GNAME71238(G71238,G69680,G69510);
  and GNAME71239(G71239,G69615,G69680);
  or GNAME71240(G71240,G71239,G71238,G71237);
  xor GNAME71250(G71250,G71251,G69540);
  xor GNAME71251(G71251,G69630,G69710);
  and GNAME71252(G71252,G69630,G69540);
  and GNAME71253(G71253,G69710,G69540);
  and GNAME71254(G71254,G69630,G69710);
  or GNAME71255(G71255,G71254,G71253,G71252);
  xor GNAME71265(G71265,G71266,G69660);
  xor GNAME71266(G71266,G69780,G69830);
  and GNAME71267(G71267,G69780,G69660);
  and GNAME71268(G71268,G69830,G69660);
  and GNAME71269(G71269,G69780,G69830);
  or GNAME71270(G71270,G71269,G71268,G71267);
  xor GNAME71280(G71280,G71281,G69690);
  xor GNAME71281(G71281,G69795,G69860);
  and GNAME71282(G71282,G69795,G69690);
  and GNAME71283(G71283,G69860,G69690);
  and GNAME71284(G71284,G69795,G69860);
  or GNAME71285(G71285,G71284,G71283,G71282);
  xor GNAME71295(G71295,G71296,G69720);
  xor GNAME71296(G71296,G69810,G69890);
  and GNAME71297(G71297,G69810,G69720);
  and GNAME71298(G71298,G69890,G69720);
  and GNAME71299(G71299,G69810,G69890);
  or GNAME71300(G71300,G71299,G71298,G71297);
  xor GNAME71310(G71310,G71311,G71330);
  xor GNAME71311(G71311,G68115,G68165);
  and GNAME71312(G71312,G68115,G71330);
  and GNAME71313(G71313,G68165,G71330);
  and GNAME71314(G71314,G68115,G68165);
  or GNAME71315(G71315,G71314,G71313,G71312);
  xor GNAME71325(G71325,G71326,G71345);
  xor GNAME71326(G71326,G68160,G68255);
  and GNAME71327(G71327,G68160,G71345);
  and GNAME71328(G71328,G68255,G71345);
  and GNAME71329(G71329,G68160,G68255);
  or GNAME71330(G71330,G71329,G71328,G71327);
  xor GNAME71340(G71340,G71341,G71360);
  xor GNAME71341(G71341,G68270,G68250);
  and GNAME71342(G71342,G68270,G71360);
  and GNAME71343(G71343,G68250,G71360);
  and GNAME71344(G71344,G68270,G68250);
  or GNAME71345(G71345,G71344,G71343,G71342);
  xor GNAME71355(G71355,G71356,G71375);
  xor GNAME71356(G71356,G68435,G68265);
  and GNAME71357(G71357,G68435,G71375);
  and GNAME71358(G71358,G68265,G71375);
  and GNAME71359(G71359,G68435,G68265);
  or GNAME71360(G71360,G71359,G71358,G71357);
  xor GNAME71370(G71370,G71371,G71390);
  xor GNAME71371(G71371,G68450,G68430);
  and GNAME71372(G71372,G68450,G71390);
  and GNAME71373(G71373,G68430,G71390);
  and GNAME71374(G71374,G68450,G68430);
  or GNAME71375(G71375,G71374,G71373,G71372);
  xor GNAME71385(G71385,G71386,G71405);
  xor GNAME71386(G71386,G70460,G68445);
  and GNAME71387(G71387,G70460,G71405);
  and GNAME71388(G71388,G68445,G71405);
  and GNAME71389(G71389,G70460,G68445);
  or GNAME71390(G71390,G71389,G71388,G71387);
  xor GNAME71400(G71400,G71401,G71420);
  xor GNAME71401(G71401,G68660,G70455);
  and GNAME71402(G71402,G68660,G71420);
  and GNAME71403(G71403,G70455,G71420);
  and GNAME71404(G71404,G68660,G70455);
  or GNAME71405(G71405,G71404,G71403,G71402);
  xor GNAME71415(G71415,G71416,G71435);
  xor GNAME71416(G71416,G68750,G68655);
  and GNAME71417(G71417,G68750,G71435);
  and GNAME71418(G71418,G68655,G71435);
  and GNAME71419(G71419,G68750,G68655);
  or GNAME71420(G71420,G71419,G71418,G71417);
  xor GNAME71430(G71430,G71431,G72080);
  xor GNAME71431(G71431,G70595,G68745);
  and GNAME71432(G71432,G70595,G72080);
  and GNAME71433(G71433,G68745,G72080);
  and GNAME71434(G71434,G70595,G68745);
  or GNAME71435(G71435,G71434,G71433,G71432);
  xor GNAME71445(G71445,G71446,G71465);
  xor GNAME71446(G71446,G68130,G68180);
  and GNAME71447(G71447,G68130,G71465);
  and GNAME71448(G71448,G68180,G71465);
  and GNAME71449(G71449,G68130,G68180);
  or GNAME71450(G71450,G71449,G71448,G71447);
  xor GNAME71460(G71460,G71461,G71510);
  xor GNAME71461(G71461,G68175,G68285);
  and GNAME71462(G71462,G68175,G71510);
  and GNAME71463(G71463,G68285,G71510);
  and GNAME71464(G71464,G68175,G68285);
  or GNAME71465(G71465,G71464,G71463,G71462);
  xor GNAME71475(G71475,G71476,G71495);
  xor GNAME71476(G71476,G68145,G68195);
  and GNAME71477(G71477,G68145,G71495);
  and GNAME71478(G71478,G68195,G71495);
  and GNAME71479(G71479,G68145,G68195);
  or GNAME71480(G71480,G71479,G71478,G71477);
  xor GNAME71490(G71490,G71491,G71555);
  xor GNAME71491(G71491,G68190,G68300);
  and GNAME71492(G71492,G68190,G71555);
  and GNAME71493(G71493,G68300,G71555);
  and GNAME71494(G71494,G68190,G68300);
  or GNAME71495(G71495,G71494,G71493,G71492);
  xor GNAME71505(G71505,G71506,G71525);
  xor GNAME71506(G71506,G68315,G68280);
  and GNAME71507(G71507,G68315,G71525);
  and GNAME71508(G71508,G68280,G71525);
  and GNAME71509(G71509,G68315,G68280);
  or GNAME71510(G71510,G71509,G71508,G71507);
  xor GNAME71520(G71520,G71521,G71585);
  xor GNAME71521(G71521,G68465,G68310);
  and GNAME71522(G71522,G68465,G71585);
  and GNAME71523(G71523,G68310,G71585);
  and GNAME71524(G71524,G68465,G68310);
  or GNAME71525(G71525,G71524,G71523,G71522);
  xor GNAME71535(G71535,G71536,G71615);
  xor GNAME71536(G71536,G69740,G71190);
  and GNAME71537(G71537,G69740,G71615);
  and GNAME71538(G71538,G71190,G71615);
  and GNAME71539(G71539,G69740,G71190);
  or GNAME71540(G71540,G71539,G71538,G71537);
  xor GNAME71550(G71550,G71551,G71570);
  xor GNAME71551(G71551,G68330,G68295);
  and GNAME71552(G71552,G68330,G71570);
  and GNAME71553(G71553,G68295,G71570);
  and GNAME71554(G71554,G68330,G68295);
  or GNAME71555(G71555,G71554,G71553,G71552);
  xor GNAME71565(G71565,G71566,G71675);
  xor GNAME71566(G71566,G68480,G68325);
  and GNAME71567(G71567,G68480,G71675);
  and GNAME71568(G71568,G68325,G71675);
  and GNAME71569(G71569,G68480,G68325);
  or GNAME71570(G71570,G71569,G71568,G71567);
  xor GNAME71580(G71580,G71581,G71600);
  xor GNAME71581(G71581,G68495,G68460);
  and GNAME71582(G71582,G68495,G71600);
  and GNAME71583(G71583,G68460,G71600);
  and GNAME71584(G71584,G68495,G68460);
  or GNAME71585(G71585,G71584,G71583,G71582);
  xor GNAME71595(G71595,G71596,G71705);
  xor GNAME71596(G71596,G70475,G68490);
  and GNAME71597(G71597,G70475,G71705);
  and GNAME71598(G71598,G68490,G71705);
  and GNAME71599(G71599,G70475,G68490);
  or GNAME71600(G71600,G71599,G71598,G71597);
  xor GNAME71610(G71610,G71611,G71630);
  xor GNAME71611(G71611,G71270,G69735);
  and GNAME71612(G71612,G71270,G71630);
  and GNAME71613(G71613,G69735,G71630);
  and GNAME71614(G71614,G71270,G69735);
  or GNAME71615(G71615,G71614,G71613,G71612);
  xor GNAME71625(G71625,G71626,G71645);
  xor GNAME71626(G71626,G69920,G71265);
  and GNAME71627(G71627,G69920,G71645);
  and GNAME71628(G71628,G71265,G71645);
  and GNAME71629(G71629,G69920,G71265);
  or GNAME71630(G71630,G71629,G71628,G71627);
  xor GNAME71640(G71640,G71641,G71660);
  xor GNAME71641(G71641,G69935,G69915);
  and GNAME71642(G71642,G69935,G71660);
  and GNAME71643(G71643,G69915,G71660);
  and GNAME71644(G71644,G69935,G69915);
  or GNAME71645(G71645,G71644,G71643,G71642);
  xor GNAME71655(G71655,G71656,G71735);
  xor GNAME71656(G71656,G69950,G69930);
  and GNAME71657(G71657,G69950,G71735);
  and GNAME71658(G71658,G69930,G71735);
  and GNAME71659(G71659,G69950,G69930);
  or GNAME71660(G71660,G71659,G71658,G71657);
  xor GNAME71670(G71670,G71671,G71690);
  xor GNAME71671(G71671,G68510,G68475);
  and GNAME71672(G71672,G68510,G71690);
  and GNAME71673(G71673,G68475,G71690);
  and GNAME71674(G71674,G68510,G68475);
  or GNAME71675(G71675,G71674,G71673,G71672);
  xor GNAME71685(G71685,G71686,G71780);
  xor GNAME71686(G71686,G70490,G68505);
  and GNAME71687(G71687,G70490,G71780);
  and GNAME71688(G71688,G68505,G71780);
  and GNAME71689(G71689,G70490,G68505);
  or GNAME71690(G71690,G71689,G71688,G71687);
  xor GNAME71700(G71700,G71701,G71720);
  xor GNAME71701(G71701,G68675,G70470);
  and GNAME71702(G71702,G68675,G71720);
  and GNAME71703(G71703,G70470,G71720);
  and GNAME71704(G71704,G68675,G70470);
  or GNAME71705(G71705,G71704,G71703,G71702);
  xor GNAME71715(G71715,G71716,G71810);
  xor GNAME71716(G71716,G68765,G68670);
  and GNAME71717(G71717,G68765,G71810);
  and GNAME71718(G71718,G68670,G71810);
  and GNAME71719(G71719,G68765,G68670);
  or GNAME71720(G71720,G71719,G71718,G71717);
  xor GNAME71730(G71730,G71731,G71750);
  xor GNAME71731(G71731,G70055,G69945);
  and GNAME71732(G71732,G70055,G71750);
  and GNAME71733(G71733,G69945,G71750);
  and GNAME71734(G71734,G70055,G69945);
  or GNAME71735(G71735,G71734,G71733,G71732);
  xor GNAME71745(G71745,G71746,G71765);
  xor GNAME71746(G71746,G70070,G70050);
  and GNAME71747(G71747,G70070,G71765);
  and GNAME71748(G71748,G70050,G71765);
  and GNAME71749(G71749,G70070,G70050);
  or GNAME71750(G71750,G71749,G71748,G71747);
  xor GNAME71760(G71760,G71761,G70325);
  xor GNAME71761(G71761,G70145,G70065);
  and GNAME71762(G71762,G70145,G70325);
  and GNAME71763(G71763,G70065,G70325);
  and GNAME71764(G71764,G70145,G70065);
  or GNAME71765(G71765,G71764,G71763,G71762);
  xor GNAME71775(G71775,G71776,G71795);
  xor GNAME71776(G71776,G68690,G70485);
  and GNAME71777(G71777,G68690,G71795);
  and GNAME71778(G71778,G70485,G71795);
  and GNAME71779(G71779,G68690,G70485);
  or GNAME71780(G71780,G71779,G71778,G71777);
  xor GNAME71790(G71790,G71791,G71825);
  xor GNAME71791(G71791,G68780,G68685);
  and GNAME71792(G71792,G68780,G71825);
  and GNAME71793(G71793,G68685,G71825);
  and GNAME71794(G71794,G68780,G68685);
  or GNAME71795(G71795,G71794,G71793,G71792);
  xor GNAME71805(G71805,G71806,G72200);
  xor GNAME71806(G71806,G70610,G68760);
  and GNAME71807(G71807,G70610,G72200);
  and GNAME71808(G71808,G68760,G72200);
  and GNAME71809(G71809,G70610,G68760);
  or GNAME71810(G71810,G71809,G71808,G71807);
  xor GNAME71820(G71820,G71821,G72215);
  xor GNAME71821(G71821,G70625,G68775);
  and GNAME71822(G71822,G70625,G72215);
  and GNAME71823(G71823,G68775,G72215);
  and GNAME71824(G71824,G70625,G68775);
  or GNAME71825(G71825,G71824,G71823,G71822);
  xor GNAME71835(G71835,G71836,G71870);
  xor GNAME71836(G71836,G69755,G71235);
  and GNAME71837(G71837,G69755,G71870);
  and GNAME71838(G71838,G71235,G71870);
  and GNAME71839(G71839,G69755,G71235);
  or GNAME71840(G71840,G71839,G71838,G71837);
  xor GNAME71850(G71850,G71851,G71900);
  xor GNAME71851(G71851,G69770,G71250);
  and GNAME71852(G71852,G69770,G71900);
  and GNAME71853(G71853,G71250,G71900);
  and GNAME71854(G71854,G69770,G71250);
  or GNAME71855(G71855,G71854,G71853,G71852);
  xor GNAME71865(G71865,G71866,G71885);
  xor GNAME71866(G71866,G71285,G69750);
  and GNAME71867(G71867,G71285,G71885);
  and GNAME71868(G71868,G69750,G71885);
  and GNAME71869(G71869,G71285,G69750);
  or GNAME71870(G71870,G71869,G71868,G71867);
  xor GNAME71880(G71880,G71881,G71930);
  xor GNAME71881(G71881,G69965,G71280);
  and GNAME71882(G71882,G69965,G71930);
  and GNAME71883(G71883,G71280,G71930);
  and GNAME71884(G71884,G69965,G71280);
  or GNAME71885(G71885,G71884,G71883,G71882);
  xor GNAME71895(G71895,G71896,G71915);
  xor GNAME71896(G71896,G71300,G69765);
  and GNAME71897(G71897,G71300,G71915);
  and GNAME71898(G71898,G69765,G71915);
  and GNAME71899(G71899,G71300,G69765);
  or GNAME71900(G71900,G71899,G71898,G71897);
  xor GNAME71910(G71910,G71911,G71960);
  xor GNAME71911(G71911,G69980,G71295);
  and GNAME71912(G71912,G69980,G71960);
  and GNAME71913(G71913,G71295,G71960);
  and GNAME71914(G71914,G69980,G71295);
  or GNAME71915(G71915,G71914,G71913,G71912);
  xor GNAME71925(G71925,G71926,G71945);
  xor GNAME71926(G71926,G69995,G69960);
  and GNAME71927(G71927,G69995,G71945);
  and GNAME71928(G71928,G69960,G71945);
  and GNAME71929(G71929,G69995,G69960);
  or GNAME71930(G71930,G71929,G71928,G71927);
  xor GNAME71940(G71940,G71941,G71990);
  xor GNAME71941(G71941,G70010,G69990);
  and GNAME71942(G71942,G70010,G71990);
  and GNAME71943(G71943,G69990,G71990);
  and GNAME71944(G71944,G70010,G69990);
  or GNAME71945(G71945,G71944,G71943,G71942);
  xor GNAME71955(G71955,G71956,G71975);
  xor GNAME71956(G71956,G70025,G69975);
  and GNAME71957(G71957,G70025,G71975);
  and GNAME71958(G71958,G69975,G71975);
  and GNAME71959(G71959,G70025,G69975);
  or GNAME71960(G71960,G71959,G71958,G71957);
  xor GNAME71970(G71970,G71971,G72020);
  xor GNAME71971(G71971,G70040,G70020);
  and GNAME71972(G71972,G70040,G72020);
  and GNAME71973(G71973,G70020,G72020);
  and GNAME71974(G71974,G70040,G70020);
  or GNAME71975(G71975,G71974,G71973,G71972);
  xor GNAME71985(G71985,G71986,G72005);
  xor GNAME71986(G71986,G70085,G70005);
  and GNAME71987(G71987,G70085,G72005);
  and GNAME71988(G71988,G70005,G72005);
  and GNAME71989(G71989,G70085,G70005);
  or GNAME71990(G71990,G71989,G71988,G71987);
  xor GNAME72000(G72000,G72001,G72050);
  xor GNAME72001(G72001,G70100,G70080);
  and GNAME72002(G72002,G70100,G72050);
  and GNAME72003(G72003,G70080,G72050);
  and GNAME72004(G72004,G70100,G70080);
  or GNAME72005(G72005,G72004,G72003,G72002);
  xor GNAME72015(G72015,G72016,G72035);
  xor GNAME72016(G72016,G70115,G70035);
  and GNAME72017(G72017,G70115,G72035);
  and GNAME72018(G72018,G70035,G72035);
  and GNAME72019(G72019,G70115,G70035);
  or GNAME72020(G72020,G72019,G72018,G72017);
  xor GNAME72030(G72030,G72031,G72065);
  xor GNAME72031(G72031,G70130,G70110);
  and GNAME72032(G72032,G70130,G72065);
  and GNAME72033(G72033,G70110,G72065);
  and GNAME72034(G72034,G70130,G70110);
  or GNAME72035(G72035,G72034,G72033,G72032);
  xor GNAME72045(G72045,G72046,G70355);
  xor GNAME72046(G72046,G70160,G70095);
  and GNAME72047(G72047,G70160,G70355);
  and GNAME72048(G72048,G70095,G70355);
  and GNAME72049(G72049,G70160,G70095);
  or GNAME72050(G72050,G72049,G72048,G72047);
  xor GNAME72060(G72060,G72061,G70370);
  xor GNAME72061(G72061,G70175,G70125);
  and GNAME72062(G72062,G70175,G70370);
  and GNAME72063(G72063,G70125,G70370);
  and GNAME72064(G72064,G70175,G70125);
  or GNAME72065(G72065,G72064,G72063,G72062);
  xor GNAME72075(G72075,G72076,G72095);
  xor GNAME72076(G72076,G70730,G70590);
  and GNAME72077(G72077,G70730,G72095);
  and GNAME72078(G72078,G70590,G72095);
  and GNAME72079(G72079,G70730,G70590);
  or GNAME72080(G72080,G72079,G72078,G72077);
  xor GNAME72090(G72090,G72091,G72110);
  xor GNAME72091(G72091,G70745,G70725);
  and GNAME72092(G72092,G70745,G72110);
  and GNAME72093(G72093,G70725,G72110);
  and GNAME72094(G72094,G70745,G70725);
  or GNAME72095(G72095,G72094,G72093,G72092);
  xor GNAME72105(G72105,G72106,G72125);
  xor GNAME72106(G72106,G70910,G70740);
  and GNAME72107(G72107,G70910,G72125);
  and GNAME72108(G72108,G70740,G72125);
  and GNAME72109(G72109,G70910,G70740);
  or GNAME72110(G72110,G72109,G72108,G72107);
  xor GNAME72120(G72120,G72121,G72140);
  xor GNAME72121(G72121,G70925,G70905);
  and GNAME72122(G72122,G70925,G72140);
  and GNAME72123(G72123,G70905,G72140);
  and GNAME72124(G72124,G70925,G70905);
  or GNAME72125(G72125,G72124,G72123,G72122);
  xor GNAME72135(G72135,G72136,G72155);
  xor GNAME72136(G72136,G71090,G70920);
  and GNAME72137(G72137,G71090,G72155);
  and GNAME72138(G72138,G70920,G72155);
  and GNAME72139(G72139,G71090,G70920);
  or GNAME72140(G72140,G72139,G72138,G72137);
  xor GNAME72150(G72150,G72151,G72170);
  xor GNAME72151(G72151,G71105,G71085);
  and GNAME72152(G72152,G71105,G72170);
  and GNAME72153(G72153,G71085,G72170);
  and GNAME72154(G72154,G71105,G71085);
  or GNAME72155(G72155,G72154,G72153,G72152);
  xor GNAME72165(G72165,G72166,G72185);
  xor GNAME72166(G72166,G71180,G71100);
  and GNAME72167(G72167,G71180,G72185);
  and GNAME72168(G72168,G71100,G72185);
  and GNAME72169(G72169,G71180,G71100);
  or GNAME72170(G72170,G72169,G72168,G72167);
  xor GNAME72180(G72180,G72181,G71540);
  xor GNAME72181(G72181,G71195,G71175);
  and GNAME72182(G72182,G71195,G71540);
  and GNAME72183(G72183,G71175,G71540);
  and GNAME72184(G72184,G71195,G71175);
  or GNAME72185(G72185,G72184,G72183,G72182);
  xor GNAME72195(G72195,G72196,G72230);
  xor GNAME72196(G72196,G70760,G70605);
  and GNAME72197(G72197,G70760,G72230);
  and GNAME72198(G72198,G70605,G72230);
  and GNAME72199(G72199,G70760,G70605);
  or GNAME72200(G72200,G72199,G72198,G72197);
  xor GNAME72210(G72210,G72211,G72260);
  xor GNAME72211(G72211,G70775,G70620);
  and GNAME72212(G72212,G70775,G72260);
  and GNAME72213(G72213,G70620,G72260);
  and GNAME72214(G72214,G70775,G70620);
  or GNAME72215(G72215,G72214,G72213,G72212);
  xor GNAME72225(G72225,G72226,G72245);
  xor GNAME72226(G72226,G70790,G70755);
  and GNAME72227(G72227,G70790,G72245);
  and GNAME72228(G72228,G70755,G72245);
  and GNAME72229(G72229,G70790,G70755);
  or GNAME72230(G72230,G72229,G72228,G72227);
  xor GNAME72240(G72240,G72241,G72290);
  xor GNAME72241(G72241,G70940,G70785);
  and GNAME72242(G72242,G70940,G72290);
  and GNAME72243(G72243,G70785,G72290);
  and GNAME72244(G72244,G70940,G70785);
  or GNAME72245(G72245,G72244,G72243,G72242);
  xor GNAME72255(G72255,G72256,G72275);
  xor GNAME72256(G72256,G70805,G70770);
  and GNAME72257(G72257,G70805,G72275);
  and GNAME72258(G72258,G70770,G72275);
  and GNAME72259(G72259,G70805,G70770);
  or GNAME72260(G72260,G72259,G72258,G72257);
  xor GNAME72270(G72270,G72271,G72320);
  xor GNAME72271(G72271,G70955,G70800);
  and GNAME72272(G72272,G70955,G72320);
  and GNAME72273(G72273,G70800,G72320);
  and GNAME72274(G72274,G70955,G70800);
  or GNAME72275(G72275,G72274,G72273,G72272);
  xor GNAME72285(G72285,G72286,G72305);
  xor GNAME72286(G72286,G70970,G70935);
  and GNAME72287(G72287,G70970,G72305);
  and GNAME72288(G72288,G70935,G72305);
  and GNAME72289(G72289,G70970,G70935);
  or GNAME72290(G72290,G72289,G72288,G72287);
  xor GNAME72300(G72300,G72301,G72350);
  xor GNAME72301(G72301,G71120,G70965);
  and GNAME72302(G72302,G71120,G72350);
  and GNAME72303(G72303,G70965,G72350);
  and GNAME72304(G72304,G71120,G70965);
  or GNAME72305(G72305,G72304,G72303,G72302);
  xor GNAME72315(G72315,G72316,G72335);
  xor GNAME72316(G72316,G70985,G70950);
  and GNAME72317(G72317,G70985,G72335);
  and GNAME72318(G72318,G70950,G72335);
  and GNAME72319(G72319,G70985,G70950);
  or GNAME72320(G72320,G72319,G72318,G72317);
  xor GNAME72330(G72330,G72331,G72380);
  xor GNAME72331(G72331,G71135,G70980);
  and GNAME72332(G72332,G71135,G72380);
  and GNAME72333(G72333,G70980,G72380);
  and GNAME72334(G72334,G71135,G70980);
  or GNAME72335(G72335,G72334,G72333,G72332);
  xor GNAME72345(G72345,G72346,G72365);
  xor GNAME72346(G72346,G71150,G71115);
  and GNAME72347(G72347,G71150,G72365);
  and GNAME72348(G72348,G71115,G72365);
  and GNAME72349(G72349,G71150,G71115);
  or GNAME72350(G72350,G72349,G72348,G72347);
  xor GNAME72360(G72360,G72361,G72410);
  xor GNAME72361(G72361,G71210,G71145);
  and GNAME72362(G72362,G71210,G72410);
  and GNAME72363(G72363,G71145,G72410);
  and GNAME72364(G72364,G71210,G71145);
  or GNAME72365(G72365,G72364,G72363,G72362);
  xor GNAME72375(G72375,G72376,G72395);
  xor GNAME72376(G72376,G71165,G71130);
  and GNAME72377(G72377,G71165,G72395);
  and GNAME72378(G72378,G71130,G72395);
  and GNAME72379(G72379,G71165,G71130);
  or GNAME72380(G72380,G72379,G72378,G72377);
  xor GNAME72390(G72390,G72391,G72425);
  xor GNAME72391(G72391,G71225,G71160);
  and GNAME72392(G72392,G71225,G72425);
  and GNAME72393(G72393,G71160,G72425);
  and GNAME72394(G72394,G71225,G71160);
  or GNAME72395(G72395,G72394,G72393,G72392);
  xor GNAME72405(G72405,G72406,G71840);
  xor GNAME72406(G72406,G71240,G71205);
  and GNAME72407(G72407,G71240,G71840);
  and GNAME72408(G72408,G71205,G71840);
  and GNAME72409(G72409,G71240,G71205);
  or GNAME72410(G72410,G72409,G72408,G72407);
  xor GNAME72420(G72420,G72421,G71855);
  xor GNAME72421(G72421,G71255,G71220);
  and GNAME72422(G72422,G71255,G71855);
  and GNAME72423(G72423,G71220,G71855);
  and GNAME72424(G72424,G71255,G71220);
  or GNAME72425(G72425,G72424,G72423,G72422);
  xor GNAME72435(G72435,G72436,G72935);
  xor GNAME72436(G72436,G80196,G5237);
  and GNAME72437(G72437,G80196,G72935);
  and GNAME72438(G72438,G5237,G72935);
  and GNAME72439(G72439,G80196,G5237);
  or GNAME72440(G72440,G72439,G72438,G72437);
  xor GNAME72450(G72450,G72451,G73760);
  xor GNAME72451(G72451,G80690,G80716);
  and GNAME72452(G72452,G80690,G73760);
  and GNAME72453(G72453,G80716,G73760);
  and GNAME72454(G72454,G80690,G80716);
  or GNAME72455(G72455,G72454,G72453,G72452);
  xor GNAME72465(G72465,G72466,G73823);
  xor GNAME72466(G72466,G78025,G4487);
  and GNAME72467(G72467,G78025,G73823);
  and GNAME72468(G72468,G4487,G73823);
  and GNAME72469(G72469,G78025,G4487);
  or GNAME72470(G72470,G72469,G72468,G72467);
  xor GNAME72480(G72480,G72481,G73822);
  xor GNAME72481(G72481,G78051,G78064);
  and GNAME72482(G72482,G78051,G73822);
  and GNAME72483(G72483,G78064,G73822);
  and GNAME72484(G72484,G78051,G78064);
  or GNAME72485(G72485,G72484,G72483,G72482);
  xor GNAME72495(G72495,G72496,G73821);
  xor GNAME72496(G72496,G74105,G74108);
  and GNAME72497(G72497,G74105,G73821);
  and GNAME72498(G72498,G74108,G73821);
  and GNAME72499(G72499,G74105,G74108);
  or GNAME72500(G72500,G72499,G72498,G72497);
  xor GNAME72510(G72510,G72511,G72470);
  xor GNAME72511(G72511,G78038,G4508);
  and GNAME72512(G72512,G78038,G72470);
  and GNAME72513(G72513,G4508,G72470);
  and GNAME72514(G72514,G78038,G4508);
  or GNAME72515(G72515,G72514,G72513,G72512);
  xor GNAME72525(G72525,G72526,G72515);
  xor GNAME72526(G72526,G78129,G4529);
  and GNAME72527(G72527,G78129,G72515);
  and GNAME72528(G72528,G4529,G72515);
  and GNAME72529(G72529,G78129,G4529);
  or GNAME72530(G72530,G72529,G72528,G72527);
  xor GNAME72540(G72540,G72541,G72530);
  xor GNAME72541(G72541,G78142,G4550);
  and GNAME72542(G72542,G78142,G72530);
  and GNAME72543(G72543,G4550,G72530);
  and GNAME72544(G72544,G78142,G4550);
  or GNAME72545(G72545,G72544,G72543,G72542);
  xor GNAME72555(G72555,G72556,G72545);
  xor GNAME72556(G72556,G78259,G4571);
  and GNAME72557(G72557,G78259,G72545);
  and GNAME72558(G72558,G4571,G72545);
  and GNAME72559(G72559,G78259,G4571);
  or GNAME72560(G72560,G72559,G72558,G72557);
  xor GNAME72570(G72570,G72571,G72560);
  xor GNAME72571(G72571,G78272,G4592);
  and GNAME72572(G72572,G78272,G72560);
  and GNAME72573(G72573,G4592,G72560);
  and GNAME72574(G72574,G78272,G4592);
  or GNAME72575(G72575,G72574,G72573,G72572);
  xor GNAME72585(G72585,G72586,G72575);
  xor GNAME72586(G72586,G78389,G4613);
  and GNAME72587(G72587,G78389,G72575);
  and GNAME72588(G72588,G4613,G72575);
  and GNAME72589(G72589,G78389,G4613);
  or GNAME72590(G72590,G72589,G72588,G72587);
  xor GNAME72600(G72600,G72601,G72590);
  xor GNAME72601(G72601,G78402,G4674);
  and GNAME72602(G72602,G78402,G72590);
  and GNAME72603(G72603,G4674,G72590);
  and GNAME72604(G72604,G78402,G4674);
  or GNAME72605(G72605,G72604,G72603,G72602);
  xor GNAME72615(G72615,G72616,G72605);
  xor GNAME72616(G72616,G78519,G4695);
  and GNAME72617(G72617,G78519,G72605);
  and GNAME72618(G72618,G4695,G72605);
  and GNAME72619(G72619,G78519,G4695);
  or GNAME72620(G72620,G72619,G72618,G72617);
  xor GNAME72630(G72630,G72631,G72620);
  xor GNAME72631(G72631,G78532,G4716);
  and GNAME72632(G72632,G78532,G72620);
  and GNAME72633(G72633,G4716,G72620);
  and GNAME72634(G72634,G78532,G4716);
  or GNAME72635(G72635,G72634,G72633,G72632);
  xor GNAME72645(G72645,G72646,G72635);
  xor GNAME72646(G72646,G78649,G4737);
  and GNAME72647(G72647,G78649,G72635);
  and GNAME72648(G72648,G4737,G72635);
  and GNAME72649(G72649,G78649,G4737);
  or GNAME72650(G72650,G72649,G72648,G72647);
  xor GNAME72660(G72660,G72661,G72650);
  xor GNAME72661(G72661,G78662,G4758);
  and GNAME72662(G72662,G78662,G72650);
  and GNAME72663(G72663,G4758,G72650);
  and GNAME72664(G72664,G78662,G4758);
  or GNAME72665(G72665,G72664,G72663,G72662);
  xor GNAME72675(G72675,G72676,G72665);
  xor GNAME72676(G72676,G78779,G4779);
  and GNAME72677(G72677,G78779,G72665);
  and GNAME72678(G72678,G4779,G72665);
  and GNAME72679(G72679,G78779,G4779);
  or GNAME72680(G72680,G72679,G72678,G72677);
  xor GNAME72690(G72690,G72691,G72680);
  xor GNAME72691(G72691,G78792,G4800);
  and GNAME72692(G72692,G78792,G72680);
  and GNAME72693(G72693,G4800,G72680);
  and GNAME72694(G72694,G78792,G4800);
  or GNAME72695(G72695,G72694,G72693,G72692);
  xor GNAME72705(G72705,G72706,G72695);
  xor GNAME72706(G72706,G78909,G4821);
  and GNAME72707(G72707,G78909,G72695);
  and GNAME72708(G72708,G4821,G72695);
  and GNAME72709(G72709,G78909,G4821);
  or GNAME72710(G72710,G72709,G72708,G72707);
  xor GNAME72720(G72720,G72721,G72710);
  xor GNAME72721(G72721,G78922,G4882);
  and GNAME72722(G72722,G78922,G72710);
  and GNAME72723(G72723,G4882,G72710);
  and GNAME72724(G72724,G78922,G4882);
  or GNAME72725(G72725,G72724,G72723,G72722);
  xor GNAME72735(G72735,G72736,G72725);
  xor GNAME72736(G72736,G79039,G4903);
  and GNAME72737(G72737,G79039,G72725);
  and GNAME72738(G72738,G4903,G72725);
  and GNAME72739(G72739,G79039,G4903);
  or GNAME72740(G72740,G72739,G72738,G72737);
  xor GNAME72750(G72750,G72751,G72740);
  xor GNAME72751(G72751,G79052,G4924);
  and GNAME72752(G72752,G79052,G72740);
  and GNAME72753(G72753,G4924,G72740);
  and GNAME72754(G72754,G79052,G4924);
  or GNAME72755(G72755,G72754,G72753,G72752);
  xor GNAME72765(G72765,G72766,G72755);
  xor GNAME72766(G72766,G79234,G4945);
  and GNAME72767(G72767,G79234,G72755);
  and GNAME72768(G72768,G4945,G72755);
  and GNAME72769(G72769,G79234,G4945);
  or GNAME72770(G72770,G72769,G72768,G72767);
  xor GNAME72780(G72780,G72781,G72770);
  xor GNAME72781(G72781,G79247,G4966);
  and GNAME72782(G72782,G79247,G72770);
  and GNAME72783(G72783,G4966,G72770);
  and GNAME72784(G72784,G79247,G4966);
  or GNAME72785(G72785,G72784,G72783,G72782);
  xor GNAME72795(G72795,G72796,G72785);
  xor GNAME72796(G72796,G79416,G4987);
  and GNAME72797(G72797,G79416,G72785);
  and GNAME72798(G72798,G4987,G72785);
  and GNAME72799(G72799,G79416,G4987);
  or GNAME72800(G72800,G72799,G72798,G72797);
  xor GNAME72810(G72810,G72811,G72800);
  xor GNAME72811(G72811,G79429,G5008);
  and GNAME72812(G72812,G79429,G72800);
  and GNAME72813(G72813,G5008,G72800);
  and GNAME72814(G72814,G79429,G5008);
  or GNAME72815(G72815,G72814,G72813,G72812);
  xor GNAME72825(G72825,G72826,G72815);
  xor GNAME72826(G72826,G79442,G5029);
  and GNAME72827(G72827,G79442,G72815);
  and GNAME72828(G72828,G5029,G72815);
  and GNAME72829(G72829,G79442,G5029);
  or GNAME72830(G72830,G72829,G72828,G72827);
  xor GNAME72840(G72840,G72841,G72830);
  xor GNAME72841(G72841,G79624,G5090);
  and GNAME72842(G72842,G79624,G72830);
  and GNAME72843(G72843,G5090,G72830);
  and GNAME72844(G72844,G79624,G5090);
  or GNAME72845(G72845,G72844,G72843,G72842);
  xor GNAME72855(G72855,G72856,G72845);
  xor GNAME72856(G72856,G79637,G5111);
  and GNAME72857(G72857,G79637,G72845);
  and GNAME72858(G72858,G5111,G72845);
  and GNAME72859(G72859,G79637,G5111);
  or GNAME72860(G72860,G72859,G72858,G72857);
  xor GNAME72870(G72870,G72871,G72860);
  xor GNAME72871(G72871,G79806,G5132);
  and GNAME72872(G72872,G79806,G72860);
  and GNAME72873(G72873,G5132,G72860);
  and GNAME72874(G72874,G79806,G5132);
  or GNAME72875(G72875,G72874,G72873,G72872);
  xor GNAME72885(G72885,G72886,G72875);
  xor GNAME72886(G72886,G79819,G5153);
  and GNAME72887(G72887,G79819,G72875);
  and GNAME72888(G72888,G5153,G72875);
  and GNAME72889(G72889,G79819,G5153);
  or GNAME72890(G72890,G72889,G72888,G72887);
  xor GNAME72900(G72900,G72901,G72890);
  xor GNAME72901(G72901,G80001,G5174);
  and GNAME72902(G72902,G80001,G72890);
  and GNAME72903(G72903,G5174,G72890);
  and GNAME72904(G72904,G80001,G5174);
  or GNAME72905(G72905,G72904,G72903,G72902);
  xor GNAME72915(G72915,G72916,G72905);
  xor GNAME72916(G72916,G80014,G5195);
  and GNAME72917(G72917,G80014,G72905);
  and GNAME72918(G72918,G5195,G72905);
  and GNAME72919(G72919,G80014,G5195);
  or GNAME72920(G72920,G72919,G72918,G72917);
  xor GNAME72930(G72930,G72931,G72920);
  xor GNAME72931(G72931,G80183,G5216);
  and GNAME72932(G72932,G80183,G72920);
  and GNAME72933(G72933,G5216,G72920);
  and GNAME72934(G72934,G80183,G5216);
  or GNAME72935(G72935,G72934,G72933,G72932);
  xor GNAME72945(G72945,G72946,G72485);
  xor GNAME72946(G72946,G78155,G78181);
  and GNAME72947(G72947,G78155,G72485);
  and GNAME72948(G72948,G78181,G72485);
  and GNAME72949(G72949,G78155,G78181);
  or GNAME72950(G72950,G72949,G72948,G72947);
  xor GNAME72960(G72960,G72961,G72950);
  xor GNAME72961(G72961,G78168,G78194);
  and GNAME72962(G72962,G78168,G72950);
  and GNAME72963(G72963,G78194,G72950);
  and GNAME72964(G72964,G78168,G78194);
  or GNAME72965(G72965,G72964,G72963,G72962);
  xor GNAME72975(G72975,G72976,G72965);
  xor GNAME72976(G72976,G78285,G78311);
  and GNAME72977(G72977,G78285,G72965);
  and GNAME72978(G72978,G78311,G72965);
  and GNAME72979(G72979,G78285,G78311);
  or GNAME72980(G72980,G72979,G72978,G72977);
  xor GNAME72990(G72990,G72991,G72500);
  xor GNAME72991(G72991,G74099,G74102);
  and GNAME72992(G72992,G74099,G72500);
  and GNAME72993(G72993,G74102,G72500);
  and GNAME72994(G72994,G74099,G74102);
  or GNAME72995(G72995,G72994,G72993,G72992);
  xor GNAME73005(G73005,G73006,G72980);
  xor GNAME73006(G73006,G78298,G78324);
  and GNAME73007(G73007,G78298,G72980);
  and GNAME73008(G73008,G78324,G72980);
  and GNAME73009(G73009,G78298,G78324);
  or GNAME73010(G73010,G73009,G73008,G73007);
  xor GNAME73020(G73020,G73021,G73010);
  xor GNAME73021(G73021,G78415,G78441);
  and GNAME73022(G73022,G78415,G73010);
  and GNAME73023(G73023,G78441,G73010);
  and GNAME73024(G73024,G78415,G78441);
  or GNAME73025(G73025,G73024,G73023,G73022);
  xor GNAME73035(G73035,G73036,G72995);
  xor GNAME73036(G73036,G74093,G74096);
  and GNAME73037(G73037,G74093,G72995);
  and GNAME73038(G73038,G74096,G72995);
  and GNAME73039(G73039,G74093,G74096);
  or GNAME73040(G73040,G73039,G73038,G73037);
  xor GNAME73050(G73050,G73051,G73040);
  xor GNAME73051(G73051,G74087,G74090);
  and GNAME73052(G73052,G74087,G73040);
  and GNAME73053(G73053,G74090,G73040);
  and GNAME73054(G73054,G74087,G74090);
  or GNAME73055(G73055,G73054,G73053,G73052);
  xor GNAME73065(G73065,G73066,G73025);
  xor GNAME73066(G73066,G78428,G78454);
  and GNAME73067(G73067,G78428,G73025);
  and GNAME73068(G73068,G78454,G73025);
  and GNAME73069(G73069,G78428,G78454);
  or GNAME73070(G73070,G73069,G73068,G73067);
  xor GNAME73080(G73080,G73081,G73070);
  xor GNAME73081(G73081,G78545,G78571);
  and GNAME73082(G73082,G78545,G73070);
  and GNAME73083(G73083,G78571,G73070);
  and GNAME73084(G73084,G78545,G78571);
  or GNAME73085(G73085,G73084,G73083,G73082);
  xor GNAME73095(G73095,G73096,G73055);
  xor GNAME73096(G73096,G74081,G74084);
  and GNAME73097(G73097,G74081,G73055);
  and GNAME73098(G73098,G74084,G73055);
  and GNAME73099(G73099,G74081,G74084);
  or GNAME73100(G73100,G73099,G73098,G73097);
  xor GNAME73110(G73110,G73111,G73100);
  xor GNAME73111(G73111,G74075,G74078);
  and GNAME73112(G73112,G74075,G73100);
  and GNAME73113(G73113,G74078,G73100);
  and GNAME73114(G73114,G74075,G74078);
  or GNAME73115(G73115,G73114,G73113,G73112);
  xor GNAME73125(G73125,G73126,G73085);
  xor GNAME73126(G73126,G78558,G78584);
  and GNAME73127(G73127,G78558,G73085);
  and GNAME73128(G73128,G78584,G73085);
  and GNAME73129(G73129,G78558,G78584);
  or GNAME73130(G73130,G73129,G73128,G73127);
  xor GNAME73140(G73140,G73141,G73130);
  xor GNAME73141(G73141,G78675,G78701);
  and GNAME73142(G73142,G78675,G73130);
  and GNAME73143(G73143,G78701,G73130);
  and GNAME73144(G73144,G78675,G78701);
  or GNAME73145(G73145,G73144,G73143,G73142);
  xor GNAME73155(G73155,G73156,G73115);
  xor GNAME73156(G73156,G74069,G74072);
  and GNAME73157(G73157,G74069,G73115);
  and GNAME73158(G73158,G74072,G73115);
  and GNAME73159(G73159,G74069,G74072);
  or GNAME73160(G73160,G73159,G73158,G73157);
  xor GNAME73170(G73170,G73171,G73160);
  xor GNAME73171(G73171,G74063,G74066);
  and GNAME73172(G73172,G74063,G73160);
  and GNAME73173(G73173,G74066,G73160);
  and GNAME73174(G73174,G74063,G74066);
  or GNAME73175(G73175,G73174,G73173,G73172);
  xor GNAME73185(G73185,G73186,G73175);
  xor GNAME73186(G73186,G74057,G74060);
  and GNAME73187(G73187,G74057,G73175);
  and GNAME73188(G73188,G74060,G73175);
  and GNAME73189(G73189,G74057,G74060);
  or GNAME73190(G73190,G73189,G73188,G73187);
  xor GNAME73200(G73200,G73201,G73145);
  xor GNAME73201(G73201,G78688,G78714);
  and GNAME73202(G73202,G78688,G73145);
  and GNAME73203(G73203,G78714,G73145);
  and GNAME73204(G73204,G78688,G78714);
  or GNAME73205(G73205,G73204,G73203,G73202);
  xor GNAME73215(G73215,G73216,G73205);
  xor GNAME73216(G73216,G78805,G78831);
  and GNAME73217(G73217,G78805,G73205);
  and GNAME73218(G73218,G78831,G73205);
  and GNAME73219(G73219,G78805,G78831);
  or GNAME73220(G73220,G73219,G73218,G73217);
  xor GNAME73230(G73230,G73231,G73190);
  xor GNAME73231(G73231,G74051,G74054);
  and GNAME73232(G73232,G74051,G73190);
  and GNAME73233(G73233,G74054,G73190);
  and GNAME73234(G73234,G74051,G74054);
  or GNAME73235(G73235,G73234,G73233,G73232);
  xor GNAME73245(G73245,G73246,G73235);
  xor GNAME73246(G73246,G74045,G74048);
  and GNAME73247(G73247,G74045,G73235);
  and GNAME73248(G73248,G74048,G73235);
  and GNAME73249(G73249,G74045,G74048);
  or GNAME73250(G73250,G73249,G73248,G73247);
  xor GNAME73260(G73260,G73261,G73220);
  xor GNAME73261(G73261,G78818,G78844);
  and GNAME73262(G73262,G78818,G73220);
  and GNAME73263(G73263,G78844,G73220);
  and GNAME73264(G73264,G78818,G78844);
  or GNAME73265(G73265,G73264,G73263,G73262);
  xor GNAME73275(G73275,G73276,G73265);
  xor GNAME73276(G73276,G78935,G78961);
  and GNAME73277(G73277,G78935,G73265);
  and GNAME73278(G73278,G78961,G73265);
  and GNAME73279(G73279,G78935,G78961);
  or GNAME73280(G73280,G73279,G73278,G73277);
  xor GNAME73290(G73290,G73291,G73250);
  xor GNAME73291(G73291,G74039,G74042);
  and GNAME73292(G73292,G74039,G73250);
  and GNAME73293(G73293,G74042,G73250);
  and GNAME73294(G73294,G74039,G74042);
  or GNAME73295(G73295,G73294,G73293,G73292);
  xor GNAME73305(G73305,G73306,G73295);
  xor GNAME73306(G73306,G74033,G74036);
  and GNAME73307(G73307,G74033,G73295);
  and GNAME73308(G73308,G74036,G73295);
  and GNAME73309(G73309,G74033,G74036);
  or GNAME73310(G73310,G73309,G73308,G73307);
  xor GNAME73320(G73320,G73321,G73280);
  xor GNAME73321(G73321,G78948,G78974);
  and GNAME73322(G73322,G78948,G73280);
  and GNAME73323(G73323,G78974,G73280);
  and GNAME73324(G73324,G78948,G78974);
  or GNAME73325(G73325,G73324,G73323,G73322);
  xor GNAME73335(G73335,G73336,G73325);
  xor GNAME73336(G73336,G79065,G79091);
  and GNAME73337(G73337,G79065,G73325);
  and GNAME73338(G73338,G79091,G73325);
  and GNAME73339(G73339,G79065,G79091);
  or GNAME73340(G73340,G73339,G73338,G73337);
  xor GNAME73350(G73350,G73351,G73310);
  xor GNAME73351(G73351,G74027,G74030);
  and GNAME73352(G73352,G74027,G73310);
  and GNAME73353(G73353,G74030,G73310);
  and GNAME73354(G73354,G74027,G74030);
  or GNAME73355(G73355,G73354,G73353,G73352);
  xor GNAME73365(G73365,G73366,G73355);
  xor GNAME73366(G73366,G74021,G74024);
  and GNAME73367(G73367,G74021,G73355);
  and GNAME73368(G73368,G74024,G73355);
  and GNAME73369(G73369,G74021,G74024);
  or GNAME73370(G73370,G73369,G73368,G73367);
  xor GNAME73380(G73380,G73381,G73340);
  xor GNAME73381(G73381,G79078,G79104);
  and GNAME73382(G73382,G79078,G73340);
  and GNAME73383(G73383,G79104,G73340);
  and GNAME73384(G73384,G79078,G79104);
  or GNAME73385(G73385,G73384,G73383,G73382);
  xor GNAME73395(G73395,G73396,G73385);
  xor GNAME73396(G73396,G79260,G79286);
  and GNAME73397(G73397,G79260,G73385);
  and GNAME73398(G73398,G79286,G73385);
  and GNAME73399(G73399,G79260,G79286);
  or GNAME73400(G73400,G73399,G73398,G73397);
  xor GNAME73410(G73410,G73411,G73370);
  xor GNAME73411(G73411,G74015,G74018);
  and GNAME73412(G73412,G74015,G73370);
  and GNAME73413(G73413,G74018,G73370);
  and GNAME73414(G73414,G74015,G74018);
  or GNAME73415(G73415,G73414,G73413,G73412);
  xor GNAME73425(G73425,G73426,G73415);
  xor GNAME73426(G73426,G74009,G74012);
  and GNAME73427(G73427,G74009,G73415);
  and GNAME73428(G73428,G74012,G73415);
  and GNAME73429(G73429,G74009,G74012);
  or GNAME73430(G73430,G73429,G73428,G73427);
  xor GNAME73440(G73440,G73441,G73400);
  xor GNAME73441(G73441,G79273,G79299);
  and GNAME73442(G73442,G79273,G73400);
  and GNAME73443(G73443,G79299,G73400);
  and GNAME73444(G73444,G79273,G79299);
  or GNAME73445(G73445,G73444,G73443,G73442);
  xor GNAME73455(G73455,G73456,G73445);
  xor GNAME73456(G73456,G79455,G79481);
  and GNAME73457(G73457,G79455,G73445);
  and GNAME73458(G73458,G79481,G73445);
  and GNAME73459(G73459,G79455,G79481);
  or GNAME73460(G73460,G73459,G73458,G73457);
  xor GNAME73470(G73470,G73471,G73460);
  xor GNAME73471(G73471,G79468,G79494);
  and GNAME73472(G73472,G79468,G73460);
  and GNAME73473(G73473,G79494,G73460);
  and GNAME73474(G73474,G79468,G79494);
  or GNAME73475(G73475,G73474,G73473,G73472);
  xor GNAME73485(G73485,G73486,G73430);
  xor GNAME73486(G73486,G74003,G74006);
  and GNAME73487(G73487,G74003,G73430);
  and GNAME73488(G73488,G74006,G73430);
  and GNAME73489(G73489,G74003,G74006);
  or GNAME73490(G73490,G73489,G73488,G73487);
  xor GNAME73500(G73500,G73501,G73490);
  xor GNAME73501(G73501,G73997,G74000);
  and GNAME73502(G73502,G73997,G73490);
  and GNAME73503(G73503,G74000,G73490);
  and GNAME73504(G73504,G73997,G74000);
  or GNAME73505(G73505,G73504,G73503,G73502);
  xor GNAME73515(G73515,G73516,G73475);
  xor GNAME73516(G73516,G79650,G79676);
  and GNAME73517(G73517,G79650,G73475);
  and GNAME73518(G73518,G79676,G73475);
  and GNAME73519(G73519,G79650,G79676);
  or GNAME73520(G73520,G73519,G73518,G73517);
  xor GNAME73530(G73530,G73531,G73520);
  xor GNAME73531(G73531,G79663,G79689);
  and GNAME73532(G73532,G79663,G73520);
  and GNAME73533(G73533,G79689,G73520);
  and GNAME73534(G73534,G79663,G79689);
  or GNAME73535(G73535,G73534,G73533,G73532);
  xor GNAME73545(G73545,G73546,G73505);
  xor GNAME73546(G73546,G73991,G73994);
  and GNAME73547(G73547,G73991,G73505);
  and GNAME73548(G73548,G73994,G73505);
  and GNAME73549(G73549,G73991,G73994);
  or GNAME73550(G73550,G73549,G73548,G73547);
  xor GNAME73560(G73560,G73561,G73550);
  xor GNAME73561(G73561,G73985,G73988);
  and GNAME73562(G73562,G73985,G73550);
  and GNAME73563(G73563,G73988,G73550);
  and GNAME73564(G73564,G73985,G73988);
  or GNAME73565(G73565,G73564,G73563,G73562);
  xor GNAME73575(G73575,G73576,G73535);
  xor GNAME73576(G73576,G79832,G79858);
  and GNAME73577(G73577,G79832,G73535);
  and GNAME73578(G73578,G79858,G73535);
  and GNAME73579(G73579,G79832,G79858);
  or GNAME73580(G73580,G73579,G73578,G73577);
  xor GNAME73590(G73590,G73591,G73580);
  xor GNAME73591(G73591,G79845,G79871);
  and GNAME73592(G73592,G79845,G73580);
  and GNAME73593(G73593,G79871,G73580);
  and GNAME73594(G73594,G79845,G79871);
  or GNAME73595(G73595,G73594,G73593,G73592);
  xor GNAME73605(G73605,G73606,G73565);
  xor GNAME73606(G73606,G73979,G73982);
  and GNAME73607(G73607,G73979,G73565);
  and GNAME73608(G73608,G73982,G73565);
  and GNAME73609(G73609,G73979,G73982);
  or GNAME73610(G73610,G73609,G73608,G73607);
  xor GNAME73620(G73620,G73621,G73610);
  xor GNAME73621(G73621,G73973,G73976);
  and GNAME73622(G73622,G73973,G73610);
  and GNAME73623(G73623,G73976,G73610);
  and GNAME73624(G73624,G73973,G73976);
  or GNAME73625(G73625,G73624,G73623,G73622);
  xor GNAME73635(G73635,G73636,G73595);
  xor GNAME73636(G73636,G80027,G80053);
  and GNAME73637(G73637,G80027,G73595);
  and GNAME73638(G73638,G80053,G73595);
  and GNAME73639(G73639,G80027,G80053);
  or GNAME73640(G73640,G73639,G73638,G73637);
  xor GNAME73650(G73650,G73651,G73640);
  xor GNAME73651(G73651,G80040,G80066);
  and GNAME73652(G73652,G80040,G73640);
  and GNAME73653(G73653,G80066,G73640);
  and GNAME73654(G73654,G80040,G80066);
  or GNAME73655(G73655,G73654,G73653,G73652);
  xor GNAME73665(G73665,G73666,G73625);
  xor GNAME73666(G73666,G73967,G73970);
  and GNAME73667(G73667,G73967,G73625);
  and GNAME73668(G73668,G73970,G73625);
  and GNAME73669(G73669,G73967,G73970);
  or GNAME73670(G73670,G73669,G73668,G73667);
  xor GNAME73680(G73680,G73681,G73670);
  xor GNAME73681(G73681,G73961,G73964);
  and GNAME73682(G73682,G73961,G73670);
  and GNAME73683(G73683,G73964,G73670);
  and GNAME73684(G73684,G73961,G73964);
  or GNAME73685(G73685,G73684,G73683,G73682);
  xor GNAME73695(G73695,G73696,G73655);
  xor GNAME73696(G73696,G80209,G80235);
  and GNAME73697(G73697,G80209,G73655);
  and GNAME73698(G73698,G80235,G73655);
  and GNAME73699(G73699,G80209,G80235);
  or GNAME73700(G73700,G73699,G73698,G73697);
  xor GNAME73710(G73710,G73711,G73700);
  xor GNAME73711(G73711,G80222,G80248);
  and GNAME73712(G73712,G80222,G73700);
  and GNAME73713(G73713,G80248,G73700);
  and GNAME73714(G73714,G80222,G80248);
  or GNAME73715(G73715,G73714,G73713,G73712);
  xor GNAME73725(G73725,G73726,G73685);
  xor GNAME73726(G73726,G73955,G73958);
  and GNAME73727(G73727,G73955,G73685);
  and GNAME73728(G73728,G73958,G73685);
  and GNAME73729(G73729,G73955,G73958);
  or GNAME73730(G73730,G73729,G73728,G73727);
  xor GNAME73740(G73740,G73741,G73730);
  xor GNAME73741(G73741,G73949,G73952);
  and GNAME73742(G73742,G73949,G73730);
  and GNAME73743(G73743,G73952,G73730);
  and GNAME73744(G73744,G73949,G73952);
  or GNAME73745(G73745,G73744,G73743,G73742);
  xor GNAME73755(G73755,G73756,G73715);
  xor GNAME73756(G73756,G80677,G80703);
  and GNAME73757(G73757,G80677,G73715);
  and GNAME73758(G73758,G80703,G73715);
  and GNAME73759(G73759,G80677,G80703);
  or GNAME73760(G73760,G73759,G73758,G73757);
  xor GNAME73770(G73770,G73771,G73745);
  xor GNAME73771(G73771,G73943,G73946);
  and GNAME73772(G73772,G73943,G73745);
  and GNAME73773(G73773,G73946,G73745);
  and GNAME73774(G73774,G73943,G73946);
  or GNAME73775(G73775,G73774,G73773,G73772);
  xor GNAME73785(G73785,G73786,G73775);
  xor GNAME73786(G73786,G73937,G73940);
  and GNAME73787(G73787,G73937,G73775);
  and GNAME73788(G73788,G73940,G73775);
  and GNAME73789(G73789,G73937,G73940);
  or GNAME73790(G73790,G73789,G73788,G73787);
  xor GNAME73800(G73800,G73801,G73790);
  xor GNAME73801(G73801,G73931,G73934);
  and GNAME73802(G73802,G73931,G73790);
  and GNAME73803(G73803,G73934,G73790);
  and GNAME73804(G73804,G73931,G73934);
  or GNAME73805(G73805,G73804,G73803,G73802);
  xor GNAME73815(G73815,G73816,G73805);
  xor GNAME73816(G73816,G73925,G73928);
  and GNAME73817(G73817,G73925,G73805);
  and GNAME73818(G73818,G73928,G73805);
  and GNAME73819(G73819,G73925,G73928);
  or GNAME73820(G73820,G73819,G73818,G73817);
  and GNAME73821(G73821,G74114,G74111);
  and GNAME73822(G73822,G77934,G77960);
  and GNAME73823(G73823,G4466,G77947);
  and GNAME73824(G73824,G76198,G76207);
  and GNAME73825(G73825,G76201,G76210);
  and GNAME73826(G73826,G76204,G76213);
  and GNAME73827(G73827,G74872,G80850);
  and GNAME73828(G73828,G79195,G77696);
  or GNAME73829(G73829,G73828,G73827);
  and GNAME73830(G73830,G74866,G80850);
  and GNAME73831(G73831,G79182,G77696);
  or GNAME73832(G73832,G73831,G73830);
  and GNAME73833(G73833,G74860,G80850);
  and GNAME73834(G73834,G79169,G77696);
  or GNAME73835(G73835,G73834,G73833);
  and GNAME73836(G73836,G74848,G80850);
  and GNAME73837(G73837,G79156,G77696);
  or GNAME73838(G73838,G73837,G73836);
  and GNAME73839(G73839,G77690,G80850);
  and GNAME73840(G73840,G79117,G77696);
  or GNAME73841(G73841,G73840,G73839);
  and GNAME73842(G73842,G74890,G80850);
  and GNAME73843(G73843,G79364,G77696);
  or GNAME73844(G73844,G73843,G73842);
  and GNAME73845(G73845,G74884,G80850);
  and GNAME73846(G73846,G79351,G77696);
  or GNAME73847(G73847,G73846,G73845);
  and GNAME73848(G73848,G74878,G80850);
  and GNAME73849(G73849,G79338,G77696);
  or GNAME73850(G73850,G73849,G73848);
  and GNAME73851(G73851,G74896,G80851);
  and GNAME73852(G73852,G79377,G77696);
  or GNAME73853(G73853,G73852,G73851);
  and GNAME73854(G73854,G80851,G74902);
  and GNAME73855(G73855,G79533,G77696);
  or GNAME73856(G73856,G73855,G73854);
  and GNAME73857(G73857,G74926,G80850);
  and GNAME73858(G73858,G79585,G77696);
  or GNAME73859(G73859,G73858,G73857);
  and GNAME73860(G73860,G74920,G80850);
  and GNAME73861(G73861,G79572,G77696);
  or GNAME73862(G73862,G73861,G73860);
  and GNAME73863(G73863,G74914,G80850);
  and GNAME73864(G73864,G79559,G77696);
  or GNAME73865(G73865,G73864,G73863);
  and GNAME73866(G73866,G74908,G80850);
  and GNAME73867(G73867,G79546,G77696);
  or GNAME73868(G73868,G73867,G73866);
  and GNAME73869(G73869,G74956,G80850);
  and GNAME73870(G73870,G79910,G77696);
  or GNAME73871(G73871,G73870,G73869);
  and GNAME73872(G73872,G74950,G80850);
  and GNAME73873(G73873,G79767,G77696);
  or GNAME73874(G73874,G73873,G73872);
  and GNAME73875(G73875,G74944,G80850);
  and GNAME73876(G73876,G79754,G77696);
  or GNAME73877(G73877,G73876,G73875);
  and GNAME73878(G73878,G74938,G80850);
  and GNAME73879(G73879,G79741,G77696);
  or GNAME73880(G73880,G73879,G73878);
  and GNAME73881(G73881,G74932,G80850);
  and GNAME73882(G73882,G79728,G77696);
  or GNAME73883(G73883,G73882,G73881);
  and GNAME73884(G73884,G74980,G80850);
  and GNAME73885(G73885,G79962,G77696);
  or GNAME73886(G73886,G73885,G73884);
  and GNAME73887(G73887,G74974,G80850);
  and GNAME73888(G73888,G79949,G77696);
  or GNAME73889(G73889,G73888,G73887);
  and GNAME73890(G73890,G74968,G80850);
  and GNAME73891(G73891,G79936,G77696);
  or GNAME73892(G73892,G73891,G73890);
  and GNAME73893(G73893,G74962,G80850);
  and GNAME73894(G73894,G79923,G77696);
  or GNAME73895(G73895,G73894,G73893);
  and GNAME73896(G73896,G75010,G80850);
  and GNAME73897(G73897,G80625,G77696);
  or GNAME73898(G73898,G73897,G73896);
  and GNAME73899(G73899,G75004,G80850);
  and GNAME73900(G73900,G80144,G77696);
  or GNAME73901(G73901,G73900,G73899);
  and GNAME73902(G73902,G74998,G80850);
  and GNAME73903(G73903,G80131,G77696);
  or GNAME73904(G73904,G73903,G73902);
  and GNAME73905(G73905,G74992,G80850);
  and GNAME73906(G73906,G80118,G77696);
  or GNAME73907(G73907,G73906,G73905);
  and GNAME73908(G73908,G74986,G80850);
  and GNAME73909(G73909,G80105,G77696);
  or GNAME73910(G73910,G73909,G73908);
  and GNAME73911(G73911,G77838,G80850);
  and GNAME73912(G73912,G80599,G77696);
  or GNAME73913(G73913,G73912,G73911);
  and GNAME73914(G73914,G74854,G80850);
  and GNAME73915(G73915,G80664,G77696);
  or GNAME73916(G73916,G73915,G73914);
  and GNAME73917(G73917,G75022,G80850);
  and GNAME73918(G73918,G80651,G77696);
  or GNAME73919(G73919,G73918,G73917);
  and GNAME73920(G73920,G75016,G80850);
  and GNAME73921(G73921,G80638,G77696);
  or GNAME73922(G73922,G73921,G73920);
  and GNAME73923(G73923,G77839,G80907);
  and GNAME73924(G73924,G80586,G77773);
  or GNAME73925(G73925,G73924,G73923);
  and GNAME73926(G73926,G77840,G80906);
  and GNAME73927(G73927,G80612,G77772);
  or GNAME73928(G73928,G73927,G73926);
  and GNAME73929(G73929,G74836,G80907);
  and GNAME73930(G73930,G80092,G77773);
  or GNAME73931(G73931,G73930,G73929);
  and GNAME73932(G73932,G74842,G80906);
  and GNAME73933(G73933,G80170,G77772);
  or GNAME73934(G73934,G73933,G73932);
  and GNAME73935(G73935,G74824,G80907);
  and GNAME73936(G73936,G80079,G77773);
  or GNAME73937(G73937,G73936,G73935);
  and GNAME73938(G73938,G74830,G80906);
  and GNAME73939(G73939,G80157,G77772);
  or GNAME73940(G73940,G73939,G73938);
  and GNAME73941(G73941,G74812,G80907);
  and GNAME73942(G73942,G79897,G77773);
  or GNAME73943(G73943,G73942,G73941);
  and GNAME73944(G73944,G74818,G80906);
  and GNAME73945(G73945,G79988,G77772);
  or GNAME73946(G73946,G73945,G73944);
  and GNAME73947(G73947,G74800,G80907);
  and GNAME73948(G73948,G79884,G77773);
  or GNAME73949(G73949,G73948,G73947);
  and GNAME73950(G73950,G74806,G80906);
  and GNAME73951(G73951,G79975,G77772);
  or GNAME73952(G73952,G73951,G73950);
  and GNAME73953(G73953,G74788,G80907);
  and GNAME73954(G73954,G79715,G77773);
  or GNAME73955(G73955,G73954,G73953);
  and GNAME73956(G73956,G74794,G80906);
  and GNAME73957(G73957,G79793,G77772);
  or GNAME73958(G73958,G73957,G73956);
  and GNAME73959(G73959,G74776,G80907);
  and GNAME73960(G73960,G79702,G77773);
  or GNAME73961(G73961,G73960,G73959);
  and GNAME73962(G73962,G74782,G80906);
  and GNAME73963(G73963,G79780,G77772);
  or GNAME73964(G73964,G73963,G73962);
  and GNAME73965(G73965,G74764,G80907);
  and GNAME73966(G73966,G79520,G77773);
  or GNAME73967(G73967,G73966,G73965);
  and GNAME73968(G73968,G74770,G80906);
  and GNAME73969(G73969,G79611,G77772);
  or GNAME73970(G73970,G73969,G73968);
  and GNAME73971(G73971,G74752,G80907);
  and GNAME73972(G73972,G79507,G77773);
  or GNAME73973(G73973,G73972,G73971);
  and GNAME73974(G73974,G74758,G80906);
  and GNAME73975(G73975,G79598,G77772);
  or GNAME73976(G73976,G73975,G73974);
  and GNAME73977(G73977,G74740,G80907);
  and GNAME73978(G73978,G79325,G77773);
  or GNAME73979(G73979,G73978,G73977);
  and GNAME73980(G73980,G74746,G80906);
  and GNAME73981(G73981,G79403,G77772);
  or GNAME73982(G73982,G73981,G73980);
  and GNAME73983(G73983,G74728,G80907);
  and GNAME73984(G73984,G79312,G77773);
  or GNAME73985(G73985,G73984,G73983);
  and GNAME73986(G73986,G74734,G80906);
  and GNAME73987(G73987,G79390,G77772);
  or GNAME73988(G73988,G73987,G73986);
  and GNAME73989(G73989,G74716,G80907);
  and GNAME73990(G73990,G79143,G77773);
  or GNAME73991(G73991,G73990,G73989);
  and GNAME73992(G73992,G74722,G80906);
  and GNAME73993(G73993,G79221,G77772);
  or GNAME73994(G73994,G73993,G73992);
  and GNAME73995(G73995,G74704,G80907);
  and GNAME73996(G73996,G79130,G77773);
  or GNAME73997(G73997,G73996,G73995);
  and GNAME73998(G73998,G74710,G80906);
  and GNAME73999(G73999,G79208,G77772);
  or GNAME74000(G74000,G73999,G73998);
  and GNAME74001(G74001,G74692,G80907);
  and GNAME74002(G74002,G79000,G77773);
  or GNAME74003(G74003,G74002,G74001);
  and GNAME74004(G74004,G74698,G80906);
  and GNAME74005(G74005,G79026,G77772);
  or GNAME74006(G74006,G74005,G74004);
  and GNAME74007(G74007,G74680,G80907);
  and GNAME74008(G74008,G78987,G77773);
  or GNAME74009(G74009,G74008,G74007);
  and GNAME74010(G74010,G74686,G80906);
  and GNAME74011(G74011,G79013,G77772);
  or GNAME74012(G74012,G74011,G74010);
  and GNAME74013(G74013,G74668,G80907);
  and GNAME74014(G74014,G78870,G77773);
  or GNAME74015(G74015,G74014,G74013);
  and GNAME74016(G74016,G74674,G80906);
  and GNAME74017(G74017,G78896,G77772);
  or GNAME74018(G74018,G74017,G74016);
  and GNAME74019(G74019,G74656,G80907);
  and GNAME74020(G74020,G78857,G77773);
  or GNAME74021(G74021,G74020,G74019);
  and GNAME74022(G74022,G74662,G80906);
  and GNAME74023(G74023,G78883,G77772);
  or GNAME74024(G74024,G74023,G74022);
  and GNAME74025(G74025,G74644,G80907);
  and GNAME74026(G74026,G78740,G77773);
  or GNAME74027(G74027,G74026,G74025);
  and GNAME74028(G74028,G74650,G80906);
  and GNAME74029(G74029,G78766,G77772);
  or GNAME74030(G74030,G74029,G74028);
  and GNAME74031(G74031,G74632,G80907);
  and GNAME74032(G74032,G78727,G77773);
  or GNAME74033(G74033,G74032,G74031);
  and GNAME74034(G74034,G74638,G80906);
  and GNAME74035(G74035,G78753,G77772);
  or GNAME74036(G74036,G74035,G74034);
  and GNAME74037(G74037,G74620,G80907);
  and GNAME74038(G74038,G78610,G77773);
  or GNAME74039(G74039,G74038,G74037);
  and GNAME74040(G74040,G74626,G80906);
  and GNAME74041(G74041,G78636,G77772);
  or GNAME74042(G74042,G74041,G74040);
  and GNAME74043(G74043,G74596,G80907);
  and GNAME74044(G74044,G78597,G77773);
  or GNAME74045(G74045,G74044,G74043);
  and GNAME74046(G74046,G74602,G80906);
  and GNAME74047(G74047,G78623,G77772);
  or GNAME74048(G74048,G74047,G74046);
  and GNAME74049(G74049,G74584,G80907);
  and GNAME74050(G74050,G78480,G77773);
  or GNAME74051(G74051,G74050,G74049);
  and GNAME74052(G74052,G74590,G80906);
  and GNAME74053(G74053,G78506,G77772);
  or GNAME74054(G74054,G74053,G74052);
  and GNAME74055(G74055,G80915,G74608);
  and GNAME74056(G74056,G78467,G77773);
  or GNAME74057(G74057,G74056,G74055);
  and GNAME74058(G74058,G80914,G74614);
  and GNAME74059(G74059,G78493,G77772);
  or GNAME74060(G74060,G74059,G74058);
  and GNAME74061(G74061,G74572,G80915);
  and GNAME74062(G74062,G78350,G77773);
  or GNAME74063(G74063,G74062,G74061);
  and GNAME74064(G74064,G74578,G80914);
  and GNAME74065(G74065,G78376,G77772);
  or GNAME74066(G74066,G74065,G74064);
  and GNAME74067(G74067,G74560,G80907);
  and GNAME74068(G74068,G78337,G77773);
  or GNAME74069(G74069,G74068,G74067);
  and GNAME74070(G74070,G74566,G80906);
  and GNAME74071(G74071,G78363,G77772);
  or GNAME74072(G74072,G74071,G74070);
  and GNAME74073(G74073,G74548,G80907);
  and GNAME74074(G74074,G78220,G77773);
  or GNAME74075(G74075,G74074,G74073);
  and GNAME74076(G74076,G74554,G80906);
  and GNAME74077(G74077,G78246,G77772);
  or GNAME74078(G74078,G74077,G74076);
  and GNAME74079(G74079,G74536,G80907);
  and GNAME74080(G74080,G78207,G77773);
  or GNAME74081(G74081,G74080,G74079);
  and GNAME74082(G74082,G74542,G80906);
  and GNAME74083(G74083,G78233,G77772);
  or GNAME74084(G74084,G74083,G74082);
  and GNAME74085(G74085,G74524,G80907);
  and GNAME74086(G74086,G78090,G77773);
  or GNAME74087(G74087,G74086,G74085);
  and GNAME74088(G74088,G74530,G80906);
  and GNAME74089(G74089,G78116,G77772);
  or GNAME74090(G74090,G74089,G74088);
  and GNAME74091(G74091,G74512,G80907);
  and GNAME74092(G74092,G78077,G77773);
  or GNAME74093(G74093,G74092,G74091);
  and GNAME74094(G74094,G74518,G80906);
  and GNAME74095(G74095,G78103,G77772);
  or GNAME74096(G74096,G74095,G74094);
  and GNAME74097(G74097,G74500,G80907);
  and GNAME74098(G74098,G77986,G77773);
  or GNAME74099(G74099,G74098,G74097);
  and GNAME74100(G74100,G74506,G80906);
  and GNAME74101(G74101,G78012,G77772);
  or GNAME74102(G74102,G74101,G74100);
  and GNAME74103(G74103,G74488,G80907);
  and GNAME74104(G74104,G77973,G77773);
  or GNAME74105(G74105,G74104,G74103);
  and GNAME74106(G74106,G74494,G80906);
  and GNAME74107(G74107,G77999,G77772);
  or GNAME74108(G74108,G74107,G74106);
  and GNAME74109(G74109,G77691,G80907);
  and GNAME74110(G74110,G77882,G77773);
  or GNAME74111(G74111,G74110,G74109);
  and GNAME74112(G74112,G77692,G80906);
  and GNAME74113(G74113,G77895,G77772);
  or GNAME74114(G74114,G74113,G74112);
  not GNAME74115(G74115,G74117);
  not GNAME74116(G74116,G80931);
  and GNAME74117(G74117,G80908,G74116);
  not GNAME74118(G74118,G74120);
  not GNAME74119(G74119,G80932);
  and GNAME74120(G74120,G80909,G74119);
  not GNAME74121(G74121,G74123);
  not GNAME74122(G74122,G80933);
  and GNAME74123(G74123,G80910,G74122);
  not GNAME74124(G74124,G74126);
  not GNAME74125(G74125,G80931);
  and GNAME74126(G74126,G80911,G74125);
  not GNAME74127(G74127,G74129);
  not GNAME74128(G74128,G80932);
  and GNAME74129(G74129,G80912,G74128);
  not GNAME74130(G74130,G74132);
  not GNAME74131(G74131,G80933);
  and GNAME74132(G74132,G80913,G74131);
  not GNAME74133(G74133,G74135);
  not GNAME74134(G74134,G80931);
  and GNAME74135(G74135,G80928,G74134);
  not GNAME74136(G74136,G74138);
  not GNAME74137(G74137,G80932);
  and GNAME74138(G74138,G80929,G74137);
  not GNAME74139(G74139,G74141);
  not GNAME74140(G74140,G80933);
  and GNAME74141(G74141,G80930,G74140);
  not GNAME74142(G74142,G74144);
  not GNAME74143(G74143,G80964);
  and GNAME74144(G74144,G80943,G74143);
  not GNAME74145(G74145,G74147);
  not GNAME74146(G74146,G80965);
  and GNAME74147(G74147,G80944,G74146);
  not GNAME74148(G74148,G74150);
  not GNAME74149(G74149,G80966);
  and GNAME74150(G74150,G80945,G74149);
  not GNAME74151(G74151,G74153);
  not GNAME74152(G74152,G80964);
  and GNAME74153(G74153,G80958,G74152);
  not GNAME74154(G74154,G74156);
  not GNAME74155(G74155,G80965);
  and GNAME74156(G74156,G80959,G74155);
  not GNAME74157(G74157,G74159);
  not GNAME74158(G74158,G80966);
  and GNAME74159(G74159,G80960,G74158);
  not GNAME74160(G74160,G74162);
  not GNAME74161(G74161,G80964);
  and GNAME74162(G74162,G80973,G74161);
  not GNAME74163(G74163,G74165);
  not GNAME74164(G74164,G80965);
  and GNAME74165(G74165,G80974,G74164);
  not GNAME74166(G74166,G74168);
  not GNAME74167(G74167,G80966);
  and GNAME74168(G74168,G80975,G74167);
  not GNAME74169(G74169,G74171);
  not GNAME74170(G74170,G80964);
  and GNAME74171(G74171,G80961,G74170);
  not GNAME74172(G74172,G74174);
  not GNAME74173(G74173,G80965);
  and GNAME74174(G74174,G80962,G74173);
  not GNAME74175(G74175,G74177);
  not GNAME74176(G74176,G80966);
  and GNAME74177(G74177,G80963,G74176);
  not GNAME74178(G74178,G74180);
  not GNAME74179(G74179,G80964);
  and GNAME74180(G74180,G80976,G74179);
  not GNAME74181(G74181,G74183);
  not GNAME74182(G74182,G80965);
  and GNAME74183(G74183,G80977,G74182);
  not GNAME74184(G74184,G74186);
  not GNAME74185(G74185,G80966);
  and GNAME74186(G74186,G80978,G74185);
  xor GNAME74187(G74187,G74188,G75175);
  xor GNAME74188(G74188,G75843,G75241);
  xor GNAME74189(G74189,G74190,G75176);
  xor GNAME74190(G74190,G75845,G75242);
  xor GNAME74191(G74191,G74192,G75177);
  xor GNAME74192(G74192,G75847,G75243);
  xor GNAME74193(G74193,G74194,G72440);
  xor GNAME74194(G74194,G80729,G5258);
  not GNAME74195(G74195,G74197);
  not GNAME74196(G74196,G80931);
  or GNAME74197(G74197,G81039,G74196);
  not GNAME74198(G74198,G74200);
  not GNAME74199(G74199,G80932);
  or GNAME74200(G74200,G81040,G74199);
  not GNAME74201(G74201,G74203);
  not GNAME74202(G74202,G80933);
  or GNAME74203(G74203,G81041,G74202);
  not GNAME74204(G74204,G74206);
  not GNAME74205(G74205,G80931);
  or GNAME74206(G74206,G80985,G74205);
  not GNAME74207(G74207,G74209);
  not GNAME74208(G74208,G80932);
  or GNAME74209(G74209,G80986,G74208);
  not GNAME74210(G74210,G74212);
  not GNAME74211(G74211,G80933);
  or GNAME74212(G74212,G80987,G74211);
  not GNAME74213(G74213,G74215);
  not GNAME74214(G74214,G72705);
  or GNAME74215(G74215,G80979,G74214);
  not GNAME74216(G74216,G74218);
  not GNAME74217(G74217,G72690);
  or GNAME74218(G74218,G80979,G74217);
  not GNAME74219(G74219,G74221);
  not GNAME74220(G74220,G72675);
  or GNAME74221(G74221,G80979,G74220);
  not GNAME74222(G74222,G74224);
  not GNAME74223(G74223,G72660);
  or GNAME74224(G74224,G80979,G74223);
  not GNAME74225(G74225,G74227);
  not GNAME74226(G74226,G72645);
  or GNAME74227(G74227,G80979,G74226);
  not GNAME74228(G74228,G74230);
  not GNAME74229(G74229,G72630);
  or GNAME74230(G74230,G80979,G74229);
  not GNAME74231(G74231,G74233);
  not GNAME74232(G74232,G72615);
  or GNAME74233(G74233,G80983,G74232);
  not GNAME74234(G74234,G74236);
  not GNAME74235(G74235,G72600);
  or GNAME74236(G74236,G80983,G74235);
  not GNAME74237(G74237,G74239);
  not GNAME74238(G74238,G72825);
  or GNAME74239(G74239,G80984,G74238);
  not GNAME74240(G74240,G74242);
  not GNAME74241(G74241,G72810);
  or GNAME74242(G74242,G80984,G74241);
  not GNAME74243(G74243,G74245);
  not GNAME74244(G74244,G72795);
  or GNAME74245(G74245,G80984,G74244);
  not GNAME74246(G74246,G74248);
  not GNAME74247(G74247,G72780);
  or GNAME74248(G74248,G80984,G74247);
  not GNAME74249(G74249,G74251);
  not GNAME74250(G74250,G72765);
  or GNAME74251(G74251,G80984,G74250);
  not GNAME74252(G74252,G74254);
  not GNAME74253(G74253,G72750);
  or GNAME74254(G74254,G80984,G74253);
  not GNAME74255(G74255,G74257);
  not GNAME74256(G74256,G72735);
  or GNAME74257(G74257,G80984,G74256);
  not GNAME74258(G74258,G74260);
  not GNAME74259(G74259,G72720);
  or GNAME74260(G74260,G80984,G74259);
  not GNAME74261(G74261,G74263);
  not GNAME74262(G74262,G72930);
  or GNAME74263(G74263,G80983,G74262);
  not GNAME74264(G74264,G74266);
  not GNAME74265(G74265,G72915);
  or GNAME74266(G74266,G80983,G74265);
  not GNAME74267(G74267,G74269);
  not GNAME74268(G74268,G72900);
  or GNAME74269(G74269,G80983,G74268);
  not GNAME74270(G74270,G74272);
  not GNAME74271(G74271,G72885);
  or GNAME74272(G74272,G80983,G74271);
  not GNAME74273(G74273,G74275);
  not GNAME74274(G74274,G72870);
  or GNAME74275(G74275,G80984,G74274);
  not GNAME74276(G74276,G74278);
  not GNAME74277(G74277,G72855);
  or GNAME74278(G74278,G80984,G74277);
  not GNAME74279(G74279,G74281);
  not GNAME74280(G74280,G72840);
  or GNAME74281(G74281,G80984,G74280);
  not GNAME74282(G74282,G74284);
  not GNAME74283(G74283,G72585);
  or GNAME74284(G74284,G80983,G74283);
  not GNAME74285(G74285,G74287);
  not GNAME74286(G74286,G72570);
  or GNAME74287(G74287,G80983,G74286);
  not GNAME74288(G74288,G74290);
  not GNAME74289(G74289,G72555);
  or GNAME74290(G74290,G80983,G74289);
  not GNAME74291(G74291,G74293);
  not GNAME74292(G74292,G72540);
  or GNAME74293(G74293,G80983,G74292);
  not GNAME74294(G74294,G74296);
  not GNAME74295(G74295,G72525);
  or GNAME74296(G74296,G80983,G74295);
  not GNAME74297(G74297,G74299);
  not GNAME74298(G74298,G72510);
  or GNAME74299(G74299,G80983,G74298);
  not GNAME74300(G74300,G74302);
  not GNAME74301(G74301,G72465);
  or GNAME74302(G74302,G80984,G74301);
  not GNAME74303(G74303,G74305);
  not GNAME74304(G74304,G80931);
  or GNAME74305(G74305,G80991,G74304);
  not GNAME74306(G74306,G74308);
  not GNAME74307(G74307,G80932);
  or GNAME74308(G74308,G80992,G74307);
  not GNAME74309(G74309,G74311);
  not GNAME74310(G74310,G80933);
  or GNAME74311(G74311,G80993,G74310);
  not GNAME74312(G74312,G74314);
  not GNAME74313(G74313,G80931);
  or GNAME74314(G74314,G81000,G74313);
  not GNAME74315(G74315,G74317);
  not GNAME74316(G74316,G80932);
  or GNAME74317(G74317,G81001,G74316);
  not GNAME74318(G74318,G74320);
  not GNAME74319(G74319,G80933);
  or GNAME74320(G74320,G81002,G74319);
  not GNAME74321(G74321,G74323);
  not GNAME74322(G74322,G80931);
  or GNAME74323(G74323,G81063,G74322);
  not GNAME74324(G74324,G74326);
  not GNAME74325(G74325,G80932);
  or GNAME74326(G74326,G81064,G74325);
  not GNAME74327(G74327,G74329);
  not GNAME74328(G74328,G80933);
  or GNAME74329(G74329,G81065,G74328);
  not GNAME74330(G74330,G74332);
  not GNAME74331(G74331,G80964);
  or GNAME74332(G74332,G81066,G74331);
  not GNAME74333(G74333,G74335);
  not GNAME74334(G74334,G80965);
  or GNAME74335(G74335,G81067,G74334);
  not GNAME74336(G74336,G74338);
  not GNAME74337(G74337,G80966);
  or GNAME74338(G74338,G81068,G74337);
  not GNAME74339(G74339,G74341);
  not GNAME74340(G74340,G80964);
  or GNAME74341(G74341,G81027,G74340);
  not GNAME74342(G74342,G74344);
  not GNAME74343(G74343,G80965);
  or GNAME74344(G74344,G81029,G74343);
  not GNAME74345(G74345,G74347);
  not GNAME74346(G74346,G80966);
  or GNAME74347(G74347,G81031,G74346);
  not GNAME74348(G74348,G74350);
  not GNAME74349(G74349,G80964);
  or GNAME74350(G74350,G81028,G74349);
  not GNAME74351(G74351,G74353);
  not GNAME74352(G74352,G80965);
  or GNAME74353(G74353,G81030,G74352);
  not GNAME74354(G74354,G74356);
  not GNAME74355(G74355,G80966);
  or GNAME74356(G74356,G81032,G74355);
  or GNAME74357(G74357,G72435,G74193);
  xor GNAME74362(G74362,G75991,G75994);
  and GNAME74363(G74363,G75991,G75994);
  xor GNAME74368(G74368,G75997,G76000);
  and GNAME74369(G74369,G75997,G76000);
  xor GNAME74374(G74374,G76003,G76006);
  and GNAME74375(G74375,G76003,G76006);
  xor GNAME74380(G74380,G76009,G76012);
  and GNAME74381(G74381,G76009,G76012);
  xor GNAME74386(G74386,G76015,G76018);
  and GNAME74387(G74387,G76015,G76018);
  xor GNAME74392(G74392,G76021,G76024);
  and GNAME74393(G74393,G76021,G76024);
  xor GNAME74398(G74398,G76045,G76048);
  and GNAME74399(G74399,G76045,G76048);
  xor GNAME74404(G74404,G76051,G76054);
  and GNAME74405(G74405,G76051,G76054);
  xor GNAME74410(G74410,G76057,G76060);
  and GNAME74411(G74411,G76057,G76060);
  xor GNAME74416(G74416,G76081,G76084);
  and GNAME74417(G74417,G76081,G76084);
  xor GNAME74422(G74422,G76087,G76090);
  and GNAME74423(G74423,G76087,G76090);
  xor GNAME74428(G74428,G76093,G76096);
  and GNAME74429(G74429,G76093,G76096);
  xor GNAME74434(G74434,G76117,G76120);
  and GNAME74435(G74435,G76117,G76120);
  xor GNAME74440(G74440,G76123,G76126);
  and GNAME74441(G74441,G76123,G76126);
  xor GNAME74446(G74446,G76129,G76132);
  and GNAME74447(G74447,G76129,G76132);
  xor GNAME74452(G74452,G76216,G77683);
  and GNAME74453(G74453,G76216,G77683);
  xor GNAME74458(G74458,G76219,G77686);
  and GNAME74459(G74459,G76219,G77686);
  xor GNAME74464(G74464,G76222,G77689);
  and GNAME74465(G74465,G76222,G77689);
  xor GNAME74470(G74470,G77665,G77668);
  and GNAME74471(G74471,G77665,G77668);
  xor GNAME74476(G74476,G77671,G77674);
  and GNAME74477(G74477,G77671,G77674);
  xor GNAME74482(G74482,G77677,G77680);
  and GNAME74483(G74483,G77677,G77680);
  xor GNAME74488(G74488,G77973,G77882);
  and GNAME74489(G74489,G77973,G77882);
  xor GNAME74494(G74494,G77999,G77895);
  and GNAME74495(G74495,G77999,G77895);
  xor GNAME74500(G74500,G77986,G74489);
  and GNAME74501(G74501,G77986,G74489);
  xor GNAME74506(G74506,G78012,G74495);
  and GNAME74507(G74507,G78012,G74495);
  xor GNAME74512(G74512,G78077,G74501);
  and GNAME74513(G74513,G78077,G74501);
  xor GNAME74518(G74518,G78103,G74507);
  and GNAME74519(G74519,G78103,G74507);
  xor GNAME74524(G74524,G78090,G74513);
  and GNAME74525(G74525,G78090,G74513);
  xor GNAME74530(G74530,G78116,G74519);
  and GNAME74531(G74531,G78116,G74519);
  xor GNAME74536(G74536,G78207,G74525);
  and GNAME74537(G74537,G78207,G74525);
  xor GNAME74542(G74542,G78233,G74531);
  and GNAME74543(G74543,G78233,G74531);
  xor GNAME74548(G74548,G78220,G74537);
  and GNAME74549(G74549,G78220,G74537);
  xor GNAME74554(G74554,G78246,G74543);
  and GNAME74555(G74555,G78246,G74543);
  xor GNAME74560(G74560,G78337,G74549);
  and GNAME74561(G74561,G78337,G74549);
  xor GNAME74566(G74566,G78363,G74555);
  and GNAME74567(G74567,G78363,G74555);
  xor GNAME74572(G74572,G78350,G74561);
  and GNAME74573(G74573,G78350,G74561);
  xor GNAME74578(G74578,G78376,G74567);
  and GNAME74579(G74579,G78376,G74567);
  xor GNAME74584(G74584,G78480,G74609);
  and GNAME74585(G74585,G78480,G74609);
  xor GNAME74590(G74590,G78506,G74615);
  and GNAME74591(G74591,G78506,G74615);
  xor GNAME74596(G74596,G78597,G74585);
  and GNAME74597(G74597,G78597,G74585);
  xor GNAME74602(G74602,G78623,G74591);
  and GNAME74603(G74603,G78623,G74591);
  xor GNAME74608(G74608,G78467,G74573);
  and GNAME74609(G74609,G78467,G74573);
  xor GNAME74614(G74614,G78493,G74579);
  and GNAME74615(G74615,G78493,G74579);
  xor GNAME74620(G74620,G78610,G74597);
  and GNAME74621(G74621,G78610,G74597);
  xor GNAME74626(G74626,G78636,G74603);
  and GNAME74627(G74627,G78636,G74603);
  xor GNAME74632(G74632,G78727,G74621);
  and GNAME74633(G74633,G78727,G74621);
  xor GNAME74638(G74638,G78753,G74627);
  and GNAME74639(G74639,G78753,G74627);
  xor GNAME74644(G74644,G78740,G74633);
  and GNAME74645(G74645,G78740,G74633);
  xor GNAME74650(G74650,G78766,G74639);
  and GNAME74651(G74651,G78766,G74639);
  xor GNAME74656(G74656,G78857,G74645);
  and GNAME74657(G74657,G78857,G74645);
  xor GNAME74662(G74662,G78883,G74651);
  and GNAME74663(G74663,G78883,G74651);
  xor GNAME74668(G74668,G78870,G74657);
  and GNAME74669(G74669,G78870,G74657);
  xor GNAME74674(G74674,G78896,G74663);
  and GNAME74675(G74675,G78896,G74663);
  xor GNAME74680(G74680,G78987,G74669);
  and GNAME74681(G74681,G78987,G74669);
  xor GNAME74686(G74686,G79013,G74675);
  and GNAME74687(G74687,G79013,G74675);
  xor GNAME74692(G74692,G79000,G74681);
  and GNAME74693(G74693,G79000,G74681);
  xor GNAME74698(G74698,G79026,G74687);
  and GNAME74699(G74699,G79026,G74687);
  xor GNAME74704(G74704,G79130,G74693);
  and GNAME74705(G74705,G79130,G74693);
  xor GNAME74710(G74710,G79208,G74699);
  and GNAME74711(G74711,G79208,G74699);
  xor GNAME74716(G74716,G79143,G74705);
  and GNAME74717(G74717,G79143,G74705);
  xor GNAME74722(G74722,G79221,G74711);
  and GNAME74723(G74723,G79221,G74711);
  xor GNAME74728(G74728,G79312,G74717);
  and GNAME74729(G74729,G79312,G74717);
  xor GNAME74734(G74734,G79390,G74723);
  and GNAME74735(G74735,G79390,G74723);
  xor GNAME74740(G74740,G79325,G74729);
  and GNAME74741(G74741,G79325,G74729);
  xor GNAME74746(G74746,G79403,G74735);
  and GNAME74747(G74747,G79403,G74735);
  xor GNAME74752(G74752,G79507,G74741);
  and GNAME74753(G74753,G79507,G74741);
  xor GNAME74758(G74758,G79598,G74747);
  and GNAME74759(G74759,G79598,G74747);
  xor GNAME74764(G74764,G79520,G74753);
  and GNAME74765(G74765,G79520,G74753);
  xor GNAME74770(G74770,G79611,G74759);
  and GNAME74771(G74771,G79611,G74759);
  xor GNAME74776(G74776,G79702,G74765);
  and GNAME74777(G74777,G79702,G74765);
  xor GNAME74782(G74782,G79780,G74771);
  and GNAME74783(G74783,G79780,G74771);
  xor GNAME74788(G74788,G79715,G74777);
  and GNAME74789(G74789,G79715,G74777);
  xor GNAME74794(G74794,G79793,G74783);
  and GNAME74795(G74795,G79793,G74783);
  xor GNAME74800(G74800,G79884,G74789);
  and GNAME74801(G74801,G79884,G74789);
  xor GNAME74806(G74806,G79975,G74795);
  and GNAME74807(G74807,G79975,G74795);
  xor GNAME74812(G74812,G79897,G74801);
  and GNAME74813(G74813,G79897,G74801);
  xor GNAME74818(G74818,G79988,G74807);
  and GNAME74819(G74819,G79988,G74807);
  xor GNAME74824(G74824,G80079,G74813);
  and GNAME74825(G74825,G80079,G74813);
  xor GNAME74830(G74830,G80157,G74819);
  and GNAME74831(G74831,G80157,G74819);
  xor GNAME74836(G74836,G80092,G74825);
  and GNAME74837(G74837,G80092,G74825);
  xor GNAME74842(G74842,G80170,G74831);
  and GNAME74843(G74843,G80170,G74831);
  xor GNAME74848(G74848,G79156,G79117);
  and GNAME74849(G74849,G79156,G79117);
  xor GNAME74854(G74854,G80664,G75023);
  and GNAME74855(G74855,G80664,G75023);
  xor GNAME74860(G74860,G79169,G74849);
  and GNAME74861(G74861,G79169,G74849);
  xor GNAME74866(G74866,G79182,G74861);
  and GNAME74867(G74867,G79182,G74861);
  xor GNAME74872(G74872,G79195,G74867);
  and GNAME74873(G74873,G79195,G74867);
  xor GNAME74878(G74878,G79338,G74873);
  and GNAME74879(G74879,G79338,G74873);
  xor GNAME74884(G74884,G79351,G74879);
  and GNAME74885(G74885,G79351,G74879);
  xor GNAME74890(G74890,G79364,G74885);
  and GNAME74891(G74891,G79364,G74885);
  xor GNAME74896(G74896,G79377,G74891);
  and GNAME74897(G74897,G79377,G74891);
  xor GNAME74902(G74902,G79533,G74897);
  and GNAME74903(G74903,G79533,G74897);
  xor GNAME74908(G74908,G79546,G74903);
  and GNAME74909(G74909,G79546,G74903);
  xor GNAME74914(G74914,G79559,G74909);
  and GNAME74915(G74915,G79559,G74909);
  xor GNAME74920(G74920,G79572,G74915);
  and GNAME74921(G74921,G79572,G74915);
  xor GNAME74926(G74926,G79585,G74921);
  and GNAME74927(G74927,G79585,G74921);
  xor GNAME74932(G74932,G79728,G74927);
  and GNAME74933(G74933,G79728,G74927);
  xor GNAME74938(G74938,G79741,G74933);
  and GNAME74939(G74939,G79741,G74933);
  xor GNAME74944(G74944,G79754,G74939);
  and GNAME74945(G74945,G79754,G74939);
  xor GNAME74950(G74950,G79767,G74945);
  and GNAME74951(G74951,G79767,G74945);
  xor GNAME74956(G74956,G79910,G74951);
  and GNAME74957(G74957,G79910,G74951);
  xor GNAME74962(G74962,G79923,G74957);
  and GNAME74963(G74963,G79923,G74957);
  xor GNAME74968(G74968,G79936,G74963);
  and GNAME74969(G74969,G79936,G74963);
  xor GNAME74974(G74974,G79949,G74969);
  and GNAME74975(G74975,G79949,G74969);
  xor GNAME74980(G74980,G79962,G74975);
  and GNAME74981(G74981,G79962,G74975);
  xor GNAME74986(G74986,G80105,G74981);
  and GNAME74987(G74987,G80105,G74981);
  xor GNAME74992(G74992,G80118,G74987);
  and GNAME74993(G74993,G80118,G74987);
  xor GNAME74998(G74998,G80131,G74993);
  and GNAME74999(G74999,G80131,G74993);
  xor GNAME75004(G75004,G80144,G74999);
  and GNAME75005(G75005,G80144,G74999);
  xor GNAME75010(G75010,G80625,G75005);
  and GNAME75011(G75011,G80625,G75005);
  xor GNAME75016(G75016,G80638,G75011);
  and GNAME75017(G75017,G80638,G75011);
  xor GNAME75022(G75022,G80651,G75017);
  and GNAME75023(G75023,G80651,G75017);
  and GNAME75030(G75030,G73824,G74348);
  and GNAME75031(G75031,G76189,G73824);
  and GNAME75032(G75032,G74348,G76189);
  or GNAME75033(G75033,G75032,G75031,G75030);
  and GNAME75040(G75040,G73825,G74351);
  and GNAME75041(G75041,G76192,G73825);
  and GNAME75042(G75042,G74351,G76192);
  or GNAME75043(G75043,G75042,G75041,G75040);
  and GNAME75050(G75050,G73826,G74354);
  and GNAME75051(G75051,G76195,G73826);
  and GNAME75052(G75052,G74354,G76195);
  or GNAME75053(G75053,G75052,G75051,G75050);
  and GNAME75060(G75060,G75033,G77656);
  and GNAME75061(G75061,G74452,G75033);
  and GNAME75062(G75062,G77656,G74452);
  or GNAME75063(G75063,G75062,G75061,G75060);
  and GNAME75070(G75070,G75063,G74453);
  and GNAME75071(G75071,G64110,G75063);
  and GNAME75072(G75072,G74453,G64110);
  or GNAME75073(G75073,G75072,G75071,G75070);
  and GNAME75080(G75080,G75043,G77659);
  and GNAME75081(G75081,G74458,G75043);
  and GNAME75082(G75082,G77659,G74458);
  or GNAME75083(G75083,G75082,G75081,G75080);
  and GNAME75090(G75090,G75083,G74459);
  and GNAME75091(G75091,G64125,G75083);
  and GNAME75092(G75092,G74459,G64125);
  or GNAME75093(G75093,G75092,G75091,G75090);
  and GNAME75100(G75100,G75053,G77662);
  and GNAME75101(G75101,G74464,G75053);
  and GNAME75102(G75102,G77662,G74464);
  or GNAME75103(G75103,G75102,G75101,G75100);
  and GNAME75110(G75110,G75103,G74465);
  and GNAME75111(G75111,G64140,G75103);
  and GNAME75112(G75112,G74465,G64140);
  or GNAME75113(G75113,G75112,G75111,G75110);
  and GNAME75120(G75120,G75073,G64115);
  and GNAME75121(G75121,G64065,G75073);
  and GNAME75122(G75122,G64115,G64065);
  or GNAME75123(G75123,G75122,G75121,G75120);
  and GNAME75130(G75130,G75123,G64070);
  and GNAME75131(G75131,G68025,G75123);
  and GNAME75132(G75132,G64070,G68025);
  or GNAME75133(G75133,G75132,G75131,G75130);
  and GNAME75140(G75140,G75093,G64130);
  and GNAME75141(G75141,G64080,G75093);
  and GNAME75142(G75142,G64130,G64080);
  or GNAME75143(G75143,G75142,G75141,G75140);
  and GNAME75150(G75150,G75143,G64085);
  and GNAME75151(G75151,G68055,G75143);
  and GNAME75152(G75152,G64085,G68055);
  or GNAME75153(G75153,G75152,G75151,G75150);
  and GNAME75160(G75160,G75113,G64145);
  and GNAME75161(G75161,G64095,G75113);
  and GNAME75162(G75162,G64145,G64095);
  or GNAME75163(G75163,G75162,G75161,G75160);
  and GNAME75170(G75170,G75163,G64100);
  and GNAME75171(G75171,G68085,G75163);
  and GNAME75172(G75172,G64100,G68085);
  or GNAME75173(G75173,G75172,G75171,G75170);
  nor GNAME75174(G75174,G75244,G80979);
  nor GNAME75175(G75175,G81036,G77700);
  nor GNAME75176(G75176,G81037,G77701);
  nor GNAME75177(G75177,G81038,G77702);
  nor GNAME75178(G75178,G81037,G77703);
  nor GNAME75179(G75179,G81036,G77704);
  nor GNAME75180(G75180,G81038,G77705);
  nor GNAME75181(G75181,G81037,G77706);
  nor GNAME75182(G75182,G81036,G77707);
  nor GNAME75183(G75183,G81038,G77708);
  nor GNAME75184(G75184,G81037,G77709);
  nor GNAME75185(G75185,G81036,G77710);
  nor GNAME75186(G75186,G81038,G77711);
  nor GNAME75187(G75187,G81037,G77712);
  nor GNAME75188(G75188,G81036,G77713);
  nor GNAME75189(G75189,G81038,G77714);
  nor GNAME75190(G75190,G81037,G77715);
  nor GNAME75191(G75191,G81036,G77716);
  nor GNAME75192(G75192,G81038,G77717);
  nor GNAME75193(G75193,G81037,G77718);
  nor GNAME75194(G75194,G81036,G77719);
  nor GNAME75195(G75195,G81038,G77720);
  nor GNAME75196(G75196,G81037,G77721);
  nor GNAME75197(G75197,G81036,G77722);
  nor GNAME75198(G75198,G81038,G77723);
  nor GNAME75199(G75199,G81037,G77724);
  nor GNAME75200(G75200,G81036,G77725);
  nor GNAME75201(G75201,G81038,G77726);
  nor GNAME75202(G75202,G81037,G77727);
  nor GNAME75203(G75203,G81036,G77728);
  nor GNAME75204(G75204,G81038,G77729);
  nor GNAME75205(G75205,G81037,G77730);
  nor GNAME75206(G75206,G81036,G77731);
  nor GNAME75207(G75207,G81038,G77732);
  nor GNAME75208(G75208,G81039,G77736);
  nor GNAME75209(G75209,G81040,G77737);
  nor GNAME75210(G75210,G81041,G77738);
  nor GNAME75211(G75211,G81039,G77739);
  nor GNAME75212(G75212,G81040,G77740);
  nor GNAME75213(G75213,G81041,G77741);
  nor GNAME75214(G75214,G81039,G77742);
  nor GNAME75215(G75215,G81040,G77743);
  nor GNAME75216(G75216,G81041,G77744);
  nor GNAME75217(G75217,G81039,G77733);
  nor GNAME75218(G75218,G81040,G77734);
  nor GNAME75219(G75219,G81041,G77735);
  nor GNAME75220(G75220,G81039,G77745);
  nor GNAME75221(G75221,G81039,G77746);
  nor GNAME75222(G75222,G81040,G77747);
  nor GNAME75223(G75223,G81041,G77748);
  nor GNAME75224(G75224,G81040,G77749);
  nor GNAME75225(G75225,G81041,G77750);
  nor GNAME75226(G75226,G81039,G77751);
  nor GNAME75227(G75227,G81039,G77752);
  nor GNAME75228(G75228,G81040,G77753);
  nor GNAME75229(G75229,G81041,G77754);
  nor GNAME75230(G75230,G81040,G77755);
  nor GNAME75231(G75231,G81041,G77756);
  nor GNAME75232(G75232,G81039,G77757);
  nor GNAME75233(G75233,G81039,G77758);
  nor GNAME75234(G75234,G81040,G77759);
  nor GNAME75235(G75235,G81041,G77760);
  nor GNAME75236(G75236,G81040,G77761);
  nor GNAME75237(G75237,G81041,G77762);
  nor GNAME75238(G75238,G81039,G77763);
  nor GNAME75239(G75239,G81040,G77764);
  nor GNAME75240(G75240,G81041,G77765);
  nor GNAME75241(G75241,G81036,G77697);
  nor GNAME75242(G75242,G81037,G77698);
  nor GNAME75243(G75243,G81038,G77699);
  xnor GNAME75244(G75244,G77947,G4466);
  xnor GNAME75245(G75245,G2678,G2657);
  xnor GNAME75246(G75246,G2262,G2241);
  xnor GNAME75247(G75247,G1846,G1825);
  xnor GNAME75248(G75248,G2636,G2615);
  xnor GNAME75249(G75249,G2220,G2199);
  xnor GNAME75250(G75250,G1804,G1783);
  xnor GNAME75251(G75251,G2552,G2491);
  xnor GNAME75252(G75252,G2136,G2075);
  xnor GNAME75253(G75253,G1720,G1659);
  xnor GNAME75254(G75254,G2594,G2573);
  xnor GNAME75255(G75255,G2178,G2157);
  xnor GNAME75256(G75256,G1762,G1741);
  xnor GNAME75257(G75257,G2470,G2449);
  xnor GNAME75258(G75258,G2054,G2033);
  xnor GNAME75259(G75259,G1638,G1617);
  xnor GNAME75260(G75260,G2428,G2407);
  xnor GNAME75261(G75261,G2012,G1991);
  xnor GNAME75262(G75262,G1596,G1575);
  xnor GNAME75263(G75263,G2386,G2365);
  xnor GNAME75264(G75264,G1970,G1949);
  xnor GNAME75265(G75265,G1554,G1533);
  xnor GNAME75266(G75266,G80852,G80855);
  xnor GNAME75267(G75267,G80852,G80864);
  xnor GNAME75268(G75268,G80853,G80856);
  xnor GNAME75269(G75269,G80853,G80865);
  xnor GNAME75270(G75270,G80854,G80857);
  xnor GNAME75271(G75271,G80854,G80866);
  xnor GNAME75272(G75272,G80852,G80861);
  xnor GNAME75273(G75273,G80858,G80855);
  xnor GNAME75274(G75274,G80858,G80864);
  xnor GNAME75275(G75275,G80852,G80873);
  xnor GNAME75276(G75276,G80853,G80862);
  xnor GNAME75277(G75277,G80859,G80856);
  xnor GNAME75278(G75278,G80859,G80865);
  xnor GNAME75279(G75279,G80853,G80874);
  xnor GNAME75280(G75280,G80854,G80863);
  xnor GNAME75281(G75281,G80860,G80857);
  xnor GNAME75282(G75282,G80860,G80866);
  xnor GNAME75283(G75283,G80854,G80875);
  xnor GNAME75284(G75284,G80852,G80882);
  xnor GNAME75285(G75285,G80858,G80873);
  xnor GNAME75286(G75286,G80853,G80883);
  xnor GNAME75287(G75287,G80859,G80874);
  xnor GNAME75288(G75288,G80854,G80884);
  xnor GNAME75289(G75289,G80860,G80875);
  xnor GNAME75290(G75290,G80858,G80861);
  xnor GNAME75291(G75291,G80867,G80855);
  xnor GNAME75292(G75292,G80852,G80870);
  xnor GNAME75293(G75293,G80859,G80862);
  xnor GNAME75294(G75294,G80868,G80856);
  xnor GNAME75295(G75295,G80860,G80863);
  xnor GNAME75296(G75296,G80869,G80857);
  xnor GNAME75297(G75297,G80853,G80871);
  xnor GNAME75298(G75298,G80854,G80872);
  xnor GNAME75299(G75299,G80867,G80864);
  xnor GNAME75300(G75300,G80867,G80861);
  xnor GNAME75301(G75301,G80876,G80855);
  xnor GNAME75302(G75302,G80852,G80879);
  xnor GNAME75303(G75303,G80858,G80870);
  xnor GNAME75304(G75304,G80868,G80865);
  xnor GNAME75305(G75305,G80868,G80862);
  xnor GNAME75306(G75306,G80877,G80856);
  xnor GNAME75307(G75307,G80869,G80866);
  xnor GNAME75308(G75308,G80869,G80863);
  xnor GNAME75309(G75309,G80878,G80857);
  xnor GNAME75310(G75310,G80853,G80880);
  xnor GNAME75311(G75311,G80859,G80871);
  xnor GNAME75312(G75312,G80854,G80881);
  xnor GNAME75313(G75313,G80860,G80872);
  xnor GNAME75314(G75314,G80867,G80873);
  xnor GNAME75315(G75315,G80852,G80891);
  xnor GNAME75316(G75316,G80858,G80882);
  xnor GNAME75317(G75317,G80858,G80879);
  xnor GNAME75318(G75318,G80885,G80855);
  xnor GNAME75319(G75319,G80868,G80874);
  xnor GNAME75320(G75320,G80853,G80892);
  xnor GNAME75321(G75321,G80859,G80883);
  xnor GNAME75322(G75322,G80869,G80875);
  xnor GNAME75323(G75323,G80854,G80893);
  xnor GNAME75324(G75324,G80860,G80884);
  xnor GNAME75325(G75325,G80859,G80880);
  xnor GNAME75326(G75326,G80886,G80856);
  xnor GNAME75327(G75327,G80860,G80881);
  xnor GNAME75328(G75328,G80887,G80857);
  xnor GNAME75329(G75329,G80867,G80870);
  xnor GNAME75330(G75330,G80852,G80888);
  xnor GNAME75331(G75331,G80876,G80864);
  xnor GNAME75332(G75332,G80876,G80861);
  xnor GNAME75333(G75333,G80868,G80871);
  xnor GNAME75334(G75334,G80853,G80889);
  xnor GNAME75335(G75335,G80877,G80865);
  xnor GNAME75336(G75336,G80877,G80862);
  xnor GNAME75337(G75337,G80869,G80872);
  xnor GNAME75338(G75338,G80854,G80890);
  xnor GNAME75339(G75339,G80878,G80866);
  xnor GNAME75340(G75340,G80878,G80863);
  xnor GNAME75341(G75341,G80858,G80891);
  xnor GNAME75342(G75342,G80859,G80892);
  xnor GNAME75343(G75343,G80860,G80893);
  xnor GNAME75344(G75344,G80876,G80873);
  xnor GNAME75345(G75345,G80852,G80898);
  xnor GNAME75346(G75346,G80867,G80882);
  xnor GNAME75347(G75347,G80885,G80864);
  xnor GNAME75348(G75348,G80885,G80861);
  xnor GNAME75349(G75349,G80894,G80855);
  xnor GNAME75350(G75350,G80867,G80879);
  xnor GNAME75351(G75351,G80852,G80897);
  xnor GNAME75352(G75352,G80876,G80870);
  xnor GNAME75353(G75353,G80858,G80888);
  xnor GNAME75354(G75354,G80877,G80874);
  xnor GNAME75355(G75355,G80853,G80900);
  xnor GNAME75356(G75356,G80868,G80883);
  xnor GNAME75357(G75357,G80878,G80875);
  xnor GNAME75358(G75358,G80854,G80902);
  xnor GNAME75359(G75359,G80869,G80884);
  xnor GNAME75360(G75360,G80886,G80865);
  xnor GNAME75361(G75361,G80886,G80862);
  xnor GNAME75362(G75362,G80895,G80856);
  xnor GNAME75363(G75363,G80868,G80880);
  xnor GNAME75364(G75364,G80853,G80899);
  xnor GNAME75365(G75365,G80877,G80871);
  xnor GNAME75366(G75366,G80859,G80889);
  xnor GNAME75367(G75367,G80887,G80866);
  xnor GNAME75368(G75368,G80887,G80863);
  xnor GNAME75369(G75369,G80896,G80857);
  xnor GNAME75370(G75370,G80869,G80881);
  xnor GNAME75371(G75371,G80854,G80901);
  xnor GNAME75372(G75372,G80878,G80872);
  xnor GNAME75373(G75373,G80860,G80890);
  xnor GNAME75374(G75374,G80885,G80873);
  xnor GNAME75375(G75375,G80852,G80916);
  xnor GNAME75376(G75376,G80894,G80864);
  xnor GNAME75377(G75377,G80876,G80882);
  xnor GNAME75378(G75378,G80858,G80898);
  xnor GNAME75379(G75379,G80867,G80891);
  xnor GNAME75380(G75380,G80876,G80879);
  xnor GNAME75381(G75381,G80867,G80888);
  xnor GNAME75382(G75382,G80885,G80870);
  xnor GNAME75383(G75383,G80858,G80897);
  xnor GNAME75384(G75384,G80852,G80917);
  xnor GNAME75385(G75385,G80894,G80861);
  xnor GNAME75386(G75386,G80903,G80855);
  xnor GNAME75387(G75387,G80886,G80874);
  xnor GNAME75388(G75388,G80853,G80919);
  xnor GNAME75389(G75389,G80895,G80865);
  xnor GNAME75390(G75390,G80877,G80883);
  xnor GNAME75391(G75391,G80859,G80900);
  xnor GNAME75392(G75392,G80868,G80892);
  xnor GNAME75393(G75393,G80887,G80875);
  xnor GNAME75394(G75394,G80854,G80921);
  xnor GNAME75395(G75395,G80896,G80866);
  xnor GNAME75396(G75396,G80878,G80884);
  xnor GNAME75397(G75397,G80860,G80902);
  xnor GNAME75398(G75398,G80869,G80893);
  xnor GNAME75399(G75399,G80877,G80880);
  xnor GNAME75400(G75400,G80868,G80889);
  xnor GNAME75401(G75401,G80886,G80871);
  xnor GNAME75402(G75402,G80859,G80899);
  xnor GNAME75403(G75403,G80853,G80920);
  xnor GNAME75404(G75404,G80895,G80862);
  xnor GNAME75405(G75405,G80904,G80856);
  xnor GNAME75406(G75406,G80878,G80881);
  xnor GNAME75407(G75407,G80869,G80890);
  xnor GNAME75408(G75408,G80887,G80872);
  xnor GNAME75409(G75409,G80860,G80901);
  xnor GNAME75410(G75410,G80854,G80922);
  xnor GNAME75411(G75411,G80896,G80863);
  xnor GNAME75412(G75412,G80905,G80857);
  xnor GNAME75413(G75413,G80908,G80918);
  xnor GNAME75414(G75414,G80876,G80891);
  xnor GNAME75415(G75415,G80894,G80873);
  xnor GNAME75416(G75416,G80867,G80898);
  xnor GNAME75417(G75417,G80903,G80864);
  xnor GNAME75418(G75418,G80885,G80882);
  xnor GNAME75419(G75419,G80858,G80916);
  xnor GNAME75420(G75420,G80876,G80888);
  xnor GNAME75421(G75421,G80867,G80897);
  xnor GNAME75422(G75422,G80885,G80879);
  xnor GNAME75423(G75423,G80858,G80917);
  xnor GNAME75424(G75424,G80908,G80940);
  xnor GNAME75425(G75425,G80894,G80870);
  xnor GNAME75426(G75426,G80903,G80861);
  xnor GNAME75427(G75427,G80909,G80923);
  xnor GNAME75428(G75428,G80877,G80892);
  xnor GNAME75429(G75429,G80895,G80874);
  xnor GNAME75430(G75430,G80868,G80900);
  xnor GNAME75431(G75431,G80904,G80865);
  xnor GNAME75432(G75432,G80886,G80883);
  xnor GNAME75433(G75433,G80859,G80919);
  xnor GNAME75434(G75434,G80910,G80924);
  xnor GNAME75435(G75435,G80878,G80893);
  xnor GNAME75436(G75436,G80896,G80875);
  xnor GNAME75437(G75437,G80869,G80902);
  xnor GNAME75438(G75438,G80905,G80866);
  xnor GNAME75439(G75439,G80887,G80884);
  xnor GNAME75440(G75440,G80860,G80921);
  xnor GNAME75441(G75441,G80877,G80889);
  xnor GNAME75442(G75442,G80868,G80899);
  xnor GNAME75443(G75443,G80886,G80880);
  xnor GNAME75444(G75444,G80859,G80920);
  xnor GNAME75445(G75445,G80909,G80941);
  xnor GNAME75446(G75446,G80895,G80871);
  xnor GNAME75447(G75447,G80904,G80862);
  xnor GNAME75448(G75448,G80878,G80890);
  xnor GNAME75449(G75449,G80869,G80901);
  xnor GNAME75450(G75450,G80887,G80881);
  xnor GNAME75451(G75451,G80860,G80922);
  xnor GNAME75452(G75452,G80910,G80942);
  xnor GNAME75453(G75453,G80896,G80872);
  xnor GNAME75454(G75454,G80905,G80863);
  xnor GNAME75455(G75455,G80925,G80855);
  xnor GNAME75456(G75456,G80926,G80856);
  xnor GNAME75457(G75457,G80927,G80857);
  xnor GNAME75458(G75458,G80876,G80898);
  xnor GNAME75459(G75459,G80867,G80916);
  xnor GNAME75460(G75460,G80885,G80891);
  xnor GNAME75461(G75461,G80911,G80918);
  xnor GNAME75462(G75462,G80908,G80935);
  xnor GNAME75463(G75463,G80894,G80882);
  xnor GNAME75464(G75464,G80903,G80873);
  xnor GNAME75465(G75465,G80876,G80897);
  xnor GNAME75466(G75466,G80867,G80917);
  xnor GNAME75467(G75467,G80885,G80888);
  xnor GNAME75468(G75468,G80911,G80940);
  xnor GNAME75469(G75469,G80908,G80934);
  xnor GNAME75470(G75470,G80894,G80879);
  xnor GNAME75471(G75471,G80903,G80870);
  xnor GNAME75472(G75472,G80877,G80900);
  xnor GNAME75473(G75473,G80868,G80919);
  xnor GNAME75474(G75474,G80886,G80892);
  xnor GNAME75475(G75475,G80912,G80923);
  xnor GNAME75476(G75476,G80909,G80937);
  xnor GNAME75477(G75477,G80895,G80883);
  xnor GNAME75478(G75478,G80904,G80874);
  xnor GNAME75479(G75479,G80878,G80902);
  xnor GNAME75480(G75480,G80869,G80921);
  xnor GNAME75481(G75481,G80887,G80893);
  xnor GNAME75482(G75482,G80913,G80924);
  xnor GNAME75483(G75483,G80910,G80939);
  xnor GNAME75484(G75484,G80896,G80884);
  xnor GNAME75485(G75485,G80905,G80875);
  xnor GNAME75486(G75486,G80877,G80899);
  xnor GNAME75487(G75487,G80868,G80920);
  xnor GNAME75488(G75488,G80886,G80889);
  xnor GNAME75489(G75489,G80912,G80941);
  xnor GNAME75490(G75490,G80909,G80936);
  xnor GNAME75491(G75491,G80895,G80880);
  xnor GNAME75492(G75492,G80904,G80871);
  xnor GNAME75493(G75493,G80878,G80901);
  xnor GNAME75494(G75494,G80869,G80922);
  xnor GNAME75495(G75495,G80887,G80890);
  xnor GNAME75496(G75496,G80913,G80942);
  xnor GNAME75497(G75497,G80910,G80938);
  xnor GNAME75498(G75498,G80896,G80881);
  xnor GNAME75499(G75499,G80905,G80872);
  xnor GNAME75500(G75500,G80925,G80864);
  xnor GNAME75501(G75501,G80925,G80861);
  xnor GNAME75502(G75502,G80926,G80865);
  xnor GNAME75503(G75503,G80927,G80866);
  xnor GNAME75504(G75504,G80926,G80862);
  xnor GNAME75505(G75505,G80927,G80863);
  xnor GNAME75506(G75506,G80876,G80916);
  xnor GNAME75507(G75507,G80928,G80918);
  xnor GNAME75508(G75508,G80885,G80898);
  xnor GNAME75509(G75509,G80911,G80935);
  xnor GNAME75510(G75510,G80908,G80949);
  xnor GNAME75511(G75511,G80894,G80891);
  xnor GNAME75512(G75512,G80903,G80882);
  xnor GNAME75513(G75513,G80876,G80917);
  xnor GNAME75514(G75514,G80928,G80940);
  xnor GNAME75515(G75515,G80885,G80897);
  xnor GNAME75516(G75516,G80911,G80934);
  xnor GNAME75517(G75517,G80908,G80946);
  xnor GNAME75518(G75518,G80894,G80888);
  xnor GNAME75519(G75519,G80903,G80879);
  xnor GNAME75520(G75520,G80877,G80919);
  xnor GNAME75521(G75521,G80929,G80923);
  xnor GNAME75522(G75522,G80886,G80900);
  xnor GNAME75523(G75523,G80912,G80937);
  xnor GNAME75524(G75524,G80909,G80950);
  xnor GNAME75525(G75525,G80895,G80892);
  xnor GNAME75526(G75526,G80904,G80883);
  xnor GNAME75527(G75527,G80878,G80921);
  xnor GNAME75528(G75528,G80930,G80924);
  xnor GNAME75529(G75529,G80887,G80902);
  xnor GNAME75530(G75530,G80913,G80939);
  xnor GNAME75531(G75531,G80910,G80951);
  xnor GNAME75532(G75532,G80896,G80893);
  xnor GNAME75533(G75533,G80905,G80884);
  xnor GNAME75534(G75534,G80877,G80920);
  xnor GNAME75535(G75535,G80929,G80941);
  xnor GNAME75536(G75536,G80886,G80899);
  xnor GNAME75537(G75537,G80912,G80936);
  xnor GNAME75538(G75538,G80909,G80954);
  xnor GNAME75539(G75539,G80895,G80889);
  xnor GNAME75540(G75540,G80904,G80880);
  xnor GNAME75541(G75541,G80878,G80922);
  xnor GNAME75542(G75542,G80930,G80942);
  xnor GNAME75543(G75543,G80887,G80901);
  xnor GNAME75544(G75544,G80913,G80938);
  xnor GNAME75545(G75545,G80910,G80957);
  xnor GNAME75546(G75546,G80896,G80890);
  xnor GNAME75547(G75547,G80905,G80881);
  xnor GNAME75548(G75548,G80925,G80873);
  xnor GNAME75549(G75549,G80925,G80870);
  xnor GNAME75550(G75550,G80926,G80874);
  xnor GNAME75551(G75551,G80927,G80875);
  xnor GNAME75552(G75552,G80926,G80871);
  xnor GNAME75553(G75553,G80927,G80872);
  xnor GNAME75554(G75554,G80943,G80918);
  xnor GNAME75555(G75555,G80928,G80935);
  xnor GNAME75556(G75556,G80885,G80916);
  xnor GNAME75557(G75557,G80911,G80949);
  xnor GNAME75558(G75558,G80908,G80947);
  xnor GNAME75559(G75559,G80894,G80898);
  xnor GNAME75560(G75560,G80903,G80891);
  xnor GNAME75561(G75561,G80943,G80940);
  xnor GNAME75562(G75562,G80928,G80934);
  xnor GNAME75563(G75563,G80885,G80917);
  xnor GNAME75564(G75564,G80911,G80946);
  xnor GNAME75565(G75565,G80908,G80948);
  xnor GNAME75566(G75566,G80894,G80897);
  xnor GNAME75567(G75567,G80903,G80888);
  xnor GNAME75568(G75568,G80944,G80923);
  xnor GNAME75569(G75569,G80929,G80937);
  xnor GNAME75570(G75570,G80886,G80919);
  xnor GNAME75571(G75571,G80912,G80950);
  xnor GNAME75572(G75572,G80909,G80953);
  xnor GNAME75573(G75573,G80895,G80900);
  xnor GNAME75574(G75574,G80904,G80892);
  xnor GNAME75575(G75575,G80945,G80924);
  xnor GNAME75576(G75576,G80930,G80939);
  xnor GNAME75577(G75577,G80887,G80921);
  xnor GNAME75578(G75578,G80913,G80951);
  xnor GNAME75579(G75579,G80910,G80956);
  xnor GNAME75580(G75580,G80896,G80902);
  xnor GNAME75581(G75581,G80905,G80893);
  xnor GNAME75582(G75582,G80944,G80941);
  xnor GNAME75583(G75583,G80929,G80936);
  xnor GNAME75584(G75584,G80886,G80920);
  xnor GNAME75585(G75585,G80912,G80954);
  xnor GNAME75586(G75586,G80909,G80952);
  xnor GNAME75587(G75587,G80895,G80899);
  xnor GNAME75588(G75588,G80904,G80889);
  xnor GNAME75589(G75589,G80945,G80942);
  xnor GNAME75590(G75590,G80930,G80938);
  xnor GNAME75591(G75591,G80887,G80922);
  xnor GNAME75592(G75592,G80913,G80957);
  xnor GNAME75593(G75593,G80910,G80955);
  xnor GNAME75594(G75594,G80896,G80901);
  xnor GNAME75595(G75595,G80905,G80890);
  xnor GNAME75596(G75596,G80925,G80882);
  xnor GNAME75597(G75597,G80925,G80879);
  xnor GNAME75598(G75598,G80926,G80883);
  xnor GNAME75599(G75599,G80927,G80884);
  xnor GNAME75600(G75600,G80926,G80880);
  xnor GNAME75601(G75601,G80927,G80881);
  xnor GNAME75602(G75602,G80894,G80917);
  xnor GNAME75603(G75603,G80895,G80920);
  xnor GNAME75604(G75604,G80896,G80922);
  xnor GNAME75605(G75605,G80943,G80935);
  xnor GNAME75606(G75606,G80928,G80949);
  xnor GNAME75607(G75607,G80958,G80918);
  xnor GNAME75608(G75608,G80911,G80947);
  xnor GNAME75609(G75609,G80908,G80967);
  xnor GNAME75610(G75610,G80894,G80916);
  xnor GNAME75611(G75611,G80903,G80898);
  xnor GNAME75612(G75612,G80943,G80934);
  xnor GNAME75613(G75613,G80928,G80946);
  xnor GNAME75614(G75614,G80958,G80940);
  xnor GNAME75615(G75615,G80911,G80948);
  xnor GNAME75616(G75616,G80903,G80897);
  xnor GNAME75617(G75617,G80944,G80937);
  xnor GNAME75618(G75618,G80929,G80950);
  xnor GNAME75619(G75619,G80959,G80923);
  xnor GNAME75620(G75620,G80912,G80953);
  xnor GNAME75621(G75621,G80909,G80969);
  xnor GNAME75622(G75622,G80895,G80919);
  xnor GNAME75623(G75623,G80904,G80900);
  xnor GNAME75624(G75624,G80945,G80939);
  xnor GNAME75625(G75625,G80930,G80951);
  xnor GNAME75626(G75626,G80960,G80924);
  xnor GNAME75627(G75627,G80913,G80956);
  xnor GNAME75628(G75628,G80910,G80971);
  xnor GNAME75629(G75629,G80896,G80921);
  xnor GNAME75630(G75630,G80905,G80902);
  xnor GNAME75631(G75631,G80944,G80936);
  xnor GNAME75632(G75632,G80929,G80954);
  xnor GNAME75633(G75633,G80959,G80941);
  xnor GNAME75634(G75634,G80912,G80952);
  xnor GNAME75635(G75635,G80904,G80899);
  xnor GNAME75636(G75636,G80945,G80938);
  xnor GNAME75637(G75637,G80930,G80957);
  xnor GNAME75638(G75638,G80960,G80942);
  xnor GNAME75639(G75639,G80913,G80955);
  xnor GNAME75640(G75640,G80905,G80901);
  xnor GNAME75641(G75641,G80925,G80891);
  xnor GNAME75642(G75642,G80926,G80892);
  xnor GNAME75643(G75643,G80927,G80893);
  xnor GNAME75644(G75644,G80911,G80931);
  xnor GNAME75645(G75645,G80912,G80932);
  xnor GNAME75646(G75646,G80913,G80933);
  xnor GNAME75647(G75647,G80908,G80931);
  xnor GNAME75648(G75648,G80909,G80932);
  xnor GNAME75649(G75649,G80910,G80933);
  xnor GNAME75650(G75650,G80958,G80949);
  xnor GNAME75651(G75651,G80959,G80950);
  xnor GNAME75652(G75652,G80960,G80951);
  xnor GNAME75653(G75653,G80908,G80968);
  xnor GNAME75654(G75654,G80958,G80935);
  xnor GNAME75655(G75655,G80903,G80916);
  xnor GNAME75656(G75656,G80928,G80947);
  xnor GNAME75657(G75657,G80911,G80967);
  xnor GNAME75658(G75658,G80943,G80949);
  xnor GNAME75659(G75659,G80903,G80917);
  xnor GNAME75660(G75660,G80928,G80948);
  xnor GNAME75661(G75661,G80911,G80968);
  xnor GNAME75662(G75662,G80961,G80918);
  xnor GNAME75663(G75663,G80961,G80940);
  xnor GNAME75664(G75664,G80943,G80946);
  xnor GNAME75665(G75665,G80958,G80934);
  xnor GNAME75666(G75666,G80909,G80970);
  xnor GNAME75667(G75667,G80959,G80937);
  xnor GNAME75668(G75668,G80904,G80919);
  xnor GNAME75669(G75669,G80929,G80953);
  xnor GNAME75670(G75670,G80912,G80969);
  xnor GNAME75671(G75671,G80944,G80950);
  xnor GNAME75672(G75672,G80910,G80972);
  xnor GNAME75673(G75673,G80960,G80939);
  xnor GNAME75674(G75674,G80905,G80921);
  xnor GNAME75675(G75675,G80930,G80956);
  xnor GNAME75676(G75676,G80913,G80971);
  xnor GNAME75677(G75677,G80945,G80951);
  xnor GNAME75678(G75678,G80904,G80920);
  xnor GNAME75679(G75679,G80929,G80952);
  xnor GNAME75680(G75680,G80912,G80970);
  xnor GNAME75681(G75681,G80962,G80923);
  xnor GNAME75682(G75682,G80962,G80941);
  xnor GNAME75683(G75683,G80944,G80954);
  xnor GNAME75684(G75684,G80959,G80936);
  xnor GNAME75685(G75685,G80905,G80922);
  xnor GNAME75686(G75686,G80930,G80955);
  xnor GNAME75687(G75687,G80913,G80972);
  xnor GNAME75688(G75688,G80963,G80924);
  xnor GNAME75689(G75689,G80963,G80942);
  xnor GNAME75690(G75690,G80945,G80957);
  xnor GNAME75691(G75691,G80960,G80938);
  xnor GNAME75692(G75692,G80925,G80888);
  xnor GNAME75693(G75693,G80925,G80898);
  xnor GNAME75694(G75694,G80925,G80897);
  xnor GNAME75695(G75695,G80926,G80889);
  xnor GNAME75696(G75696,G80926,G80900);
  xnor GNAME75697(G75697,G80927,G80890);
  xnor GNAME75698(G75698,G80927,G80902);
  xnor GNAME75699(G75699,G80926,G80899);
  xnor GNAME75700(G75700,G80927,G80901);
  xnor GNAME75701(G75701,G80943,G80948);
  xnor GNAME75702(G75702,G80943,G80967);
  xnor GNAME75703(G75703,G80961,G80934);
  xnor GNAME75704(G75704,G80961,G80949);
  xnor GNAME75705(G75705,G80958,G80947);
  xnor GNAME75706(G75706,G80944,G80952);
  xnor GNAME75707(G75707,G80944,G80969);
  xnor GNAME75708(G75708,G80962,G80936);
  xnor GNAME75709(G75709,G80962,G80950);
  xnor GNAME75710(G75710,G80959,G80953);
  xnor GNAME75711(G75711,G80945,G80955);
  xnor GNAME75712(G75712,G80945,G80971);
  xnor GNAME75713(G75713,G80963,G80938);
  xnor GNAME75714(G75714,G80963,G80951);
  xnor GNAME75715(G75715,G80960,G80956);
  xnor GNAME75716(G75716,G80928,G80967);
  xnor GNAME75717(G75717,G80961,G80935);
  xnor GNAME75718(G75718,G80973,G80918);
  xnor GNAME75719(G75719,G80943,G80947);
  xnor GNAME75720(G75720,G80928,G80968);
  xnor GNAME75721(G75721,G80973,G80940);
  xnor GNAME75722(G75722,G80958,G80946);
  xnor GNAME75723(G75723,G80929,G80969);
  xnor GNAME75724(G75724,G80962,G80937);
  xnor GNAME75725(G75725,G80974,G80923);
  xnor GNAME75726(G75726,G80944,G80953);
  xnor GNAME75727(G75727,G80930,G80971);
  xnor GNAME75728(G75728,G80963,G80939);
  xnor GNAME75729(G75729,G80975,G80924);
  xnor GNAME75730(G75730,G80945,G80956);
  xnor GNAME75731(G75731,G80929,G80970);
  xnor GNAME75732(G75732,G80974,G80941);
  xnor GNAME75733(G75733,G80959,G80954);
  xnor GNAME75734(G75734,G80930,G80972);
  xnor GNAME75735(G75735,G80975,G80942);
  xnor GNAME75736(G75736,G80960,G80957);
  xnor GNAME75737(G75737,G80925,G80916);
  xnor GNAME75738(G75738,G80925,G80917);
  xnor GNAME75739(G75739,G80926,G80919);
  xnor GNAME75740(G75740,G80926,G80920);
  xnor GNAME75741(G75741,G80927,G80921);
  xnor GNAME75742(G75742,G80927,G80922);
  xnor GNAME75743(G75743,G80928,G80931);
  xnor GNAME75744(G75744,G80929,G80932);
  xnor GNAME75745(G75745,G80930,G80933);
  xnor GNAME75746(G75746,G80943,G80931);
  xnor GNAME75747(G75747,G80944,G80932);
  xnor GNAME75748(G75748,G80945,G80933);
  xnor GNAME75749(G75749,G80973,G80934);
  xnor GNAME75750(G75750,G80958,G80967);
  xnor GNAME75751(G75751,G80961,G80947);
  xnor GNAME75752(G75752,G80974,G80936);
  xnor GNAME75753(G75753,G80975,G80938);
  xnor GNAME75754(G75754,G80959,G80969);
  xnor GNAME75755(G75755,G80962,G80953);
  xnor GNAME75756(G75756,G80960,G80971);
  xnor GNAME75757(G75757,G80963,G80956);
  xnor GNAME75758(G75758,G80958,G80948);
  xnor GNAME75759(G75759,G80943,G80968);
  xnor GNAME75760(G75760,G80961,G80946);
  xnor GNAME75761(G75761,G80973,G80935);
  xnor GNAME75762(G75762,G80973,G80949);
  xnor GNAME75763(G75763,G80958,G80968);
  xnor GNAME75764(G75764,G80959,G80952);
  xnor GNAME75765(G75765,G80944,G80970);
  xnor GNAME75766(G75766,G80962,G80954);
  xnor GNAME75767(G75767,G80974,G80937);
  xnor GNAME75768(G75768,G80960,G80955);
  xnor GNAME75769(G75769,G80945,G80972);
  xnor GNAME75770(G75770,G80963,G80957);
  xnor GNAME75771(G75771,G80975,G80939);
  xnor GNAME75772(G75772,G80974,G80950);
  xnor GNAME75773(G75773,G80975,G80951);
  xnor GNAME75774(G75774,G80959,G80970);
  xnor GNAME75775(G75775,G80960,G80972);
  xnor GNAME75776(G75776,G80976,G80918);
  xnor GNAME75777(G75777,G80976,G80940);
  xnor GNAME75778(G75778,G80976,G80935);
  xnor GNAME75779(G75779,G80976,G80934);
  xnor GNAME75780(G75780,G80977,G80923);
  xnor GNAME75781(G75781,G80977,G80941);
  xnor GNAME75782(G75782,G80978,G80924);
  xnor GNAME75783(G75783,G80978,G80942);
  xnor GNAME75784(G75784,G80977,G80937);
  xnor GNAME75785(G75785,G80977,G80936);
  xnor GNAME75786(G75786,G80978,G80939);
  xnor GNAME75787(G75787,G80978,G80938);
  xnor GNAME75788(G75788,G80958,G80964);
  xnor GNAME75789(G75789,G80959,G80965);
  xnor GNAME75790(G75790,G80960,G80966);
  xnor GNAME75791(G75791,G80961,G80964);
  xnor GNAME75792(G75792,G80962,G80965);
  xnor GNAME75793(G75793,G80963,G80966);
  xnor GNAME75794(G75794,G80961,G80967);
  xnor GNAME75795(G75795,G80961,G80948);
  xnor GNAME75796(G75796,G80973,G80946);
  xnor GNAME75797(G75797,G80973,G80947);
  xnor GNAME75798(G75798,G80962,G80952);
  xnor GNAME75799(G75799,G80962,G80969);
  xnor GNAME75800(G75800,G80974,G80954);
  xnor GNAME75801(G75801,G80974,G80953);
  xnor GNAME75802(G75802,G80963,G80955);
  xnor GNAME75803(G75803,G80963,G80971);
  xnor GNAME75804(G75804,G80975,G80957);
  xnor GNAME75805(G75805,G80975,G80956);
  xnor GNAME75806(G75806,G80973,G80948);
  xnor GNAME75807(G75807,G80961,G80968);
  xnor GNAME75808(G75808,G80974,G80952);
  xnor GNAME75809(G75809,G80962,G80970);
  xnor GNAME75810(G75810,G80975,G80955);
  xnor GNAME75811(G75811,G80963,G80972);
  xnor GNAME75812(G75812,G80976,G80946);
  xnor GNAME75813(G75813,G80976,G80949);
  xnor GNAME75814(G75814,G80977,G80950);
  xnor GNAME75815(G75815,G80978,G80951);
  xnor GNAME75816(G75816,G80977,G80954);
  xnor GNAME75817(G75817,G80978,G80957);
  xnor GNAME75818(G75818,G80973,G80967);
  xnor GNAME75819(G75819,G80973,G80968);
  xnor GNAME75820(G75820,G80974,G80969);
  xnor GNAME75821(G75821,G80974,G80970);
  xnor GNAME75822(G75822,G80975,G80971);
  xnor GNAME75823(G75823,G80975,G80972);
  xnor GNAME75824(G75824,G80976,G80947);
  xnor GNAME75825(G75825,G80976,G80948);
  xnor GNAME75826(G75826,G80977,G80953);
  xnor GNAME75827(G75827,G80977,G80952);
  xnor GNAME75828(G75828,G80978,G80956);
  xnor GNAME75829(G75829,G80978,G80955);
  xnor GNAME75830(G75830,G80976,G80967);
  xnor GNAME75831(G75831,G80976,G80968);
  xnor GNAME75832(G75832,G80977,G80969);
  xnor GNAME75833(G75833,G80977,G80970);
  xnor GNAME75834(G75834,G80978,G80971);
  xnor GNAME75835(G75835,G80978,G80972);
  xnor GNAME75836(G75836,G80976,G80964);
  xnor GNAME75837(G75837,G80977,G80965);
  xnor GNAME75838(G75838,G80978,G80966);
  xnor GNAME75839(G75839,G80973,G80964);
  xnor GNAME75840(G75840,G80974,G80965);
  xnor GNAME75841(G75841,G80975,G80966);
  and GNAME75842(G75842,G81049,G80981);
  or GNAME75843(G75843,G77766,G75842);
  and GNAME75844(G75844,G81048,G80980);
  or GNAME75845(G75845,G77767,G75844);
  and GNAME75846(G75846,G81050,G80982);
  or GNAME75847(G75847,G77768,G75846);
  and GNAME75848(G75848,G81054,G80988);
  or GNAME75849(G75849,G77769,G75848);
  and GNAME75850(G75850,G81055,G80989);
  or GNAME75851(G75851,G77770,G75850);
  and GNAME75852(G75852,G81056,G80990);
  or GNAME75853(G75853,G77771,G75852);
  and GNAME75854(G75854,G81003,G80994);
  or GNAME75855(G75855,G77774,G75854);
  and GNAME75856(G75856,G81005,G80996);
  or GNAME75857(G75857,G77776,G75856);
  and GNAME75858(G75858,G81006,G80997);
  or GNAME75859(G75859,G77777,G75858);
  and GNAME75860(G75860,G81004,G80995);
  or GNAME75861(G75861,G77775,G75860);
  and GNAME75862(G75862,G81007,G80998);
  or GNAME75863(G75863,G77778,G75862);
  and GNAME75864(G75864,G81008,G80999);
  or GNAME75865(G75865,G77779,G75864);
  and GNAME75866(G75866,G81081,G81057);
  or GNAME75867(G75867,G77780,G75866);
  and GNAME75868(G75868,G81082,G81058);
  or GNAME75869(G75869,G77781,G75868);
  and GNAME75870(G75870,G81083,G81059);
  or GNAME75871(G75871,G77782,G75870);
  and GNAME75872(G75872,G81078,G81060);
  or GNAME75873(G75873,G77786,G75872);
  and GNAME75874(G75874,G81079,G81061);
  or GNAME75875(G75875,G77783,G75874);
  and GNAME75876(G75876,G81080,G81062);
  or GNAME75877(G75877,G77784,G75876);
  and GNAME75878(G75878,G81033,G81015);
  or GNAME75879(G75879,G77785,G75878);
  and GNAME75880(G75880,G81034,G81016);
  or GNAME75881(G75881,G77787,G75880);
  and GNAME75882(G75882,G81035,G81017);
  or GNAME75883(G75883,G77788,G75882);
  and GNAME75884(G75884,G81018,G81012);
  or GNAME75885(G75885,G77789,G75884);
  and GNAME75886(G75886,G81019,G81013);
  or GNAME75887(G75887,G77790,G75886);
  and GNAME75888(G75888,G81020,G81014);
  or GNAME75889(G75889,G77791,G75888);
  or GNAME75890(G75890,G81048,G75266);
  or GNAME75891(G75891,G80980,G75267);
  nand GNAME75892(G75892,G75891,G75890);
  or GNAME75893(G75893,G81049,G75268);
  or GNAME75894(G75894,G80981,G75269);
  nand GNAME75895(G75895,G75894,G75893);
  or GNAME75896(G75896,G81050,G75270);
  or GNAME75897(G75897,G80982,G75271);
  nand GNAME75898(G75898,G75897,G75896);
  or GNAME75899(G75899,G81054,G75273);
  or GNAME75900(G75900,G80988,G75274);
  nand GNAME75901(G75901,G75900,G75899);
  or GNAME75902(G75902,G81055,G75277);
  or GNAME75903(G75903,G80989,G75278);
  nand GNAME75904(G75904,G75903,G75902);
  or GNAME75905(G75905,G81056,G75281);
  or GNAME75906(G75906,G80990,G75282);
  nand GNAME75907(G75907,G75906,G75905);
  or GNAME75908(G75908,G81003,G75291);
  or GNAME75909(G75909,G80994,G75299);
  nand GNAME75910(G75910,G75909,G75908);
  or GNAME75911(G75911,G81005,G75294);
  or GNAME75912(G75912,G80996,G75304);
  nand GNAME75913(G75913,G75912,G75911);
  or GNAME75914(G75914,G81006,G75296);
  or GNAME75915(G75915,G80997,G75307);
  nand GNAME75916(G75916,G75915,G75914);
  or GNAME75917(G75917,G81003,G75300);
  or GNAME75918(G75918,G80994,G75314);
  nand GNAME75919(G75919,G75918,G75917);
  or GNAME75920(G75920,G81005,G75305);
  or GNAME75921(G75921,G80996,G75319);
  nand GNAME75922(G75922,G75921,G75920);
  or GNAME75923(G75923,G81006,G75308);
  or GNAME75924(G75924,G80997,G75322);
  nand GNAME75925(G75925,G75924,G75923);
  or GNAME75926(G75926,G81004,G75332);
  or GNAME75927(G75927,G80995,G75344);
  nand GNAME75928(G75928,G75927,G75926);
  or GNAME75929(G75929,G81007,G75336);
  or GNAME75930(G75930,G80998,G75354);
  nand GNAME75931(G75931,G75930,G75929);
  or GNAME75932(G75932,G81008,G75340);
  or GNAME75933(G75933,G80999,G75357);
  nand GNAME75934(G75934,G75933,G75932);
  or GNAME75935(G75935,G81004,G75352);
  or GNAME75936(G75936,G80995,G75377);
  nand GNAME75937(G75937,G75936,G75935);
  or GNAME75938(G75938,G81007,G75365);
  or GNAME75939(G75939,G80998,G75390);
  nand GNAME75940(G75940,G75939,G75938);
  or GNAME75941(G75941,G81008,G75372);
  or GNAME75942(G75942,G80999,G75396);
  nand GNAME75943(G75943,G75942,G75941);
  or GNAME75944(G75944,G81033,G77785);
  or GNAME75945(G75945,G81015,G75386);
  nand GNAME75946(G75946,G75945,G75944);
  or GNAME75947(G75947,G81034,G77787);
  or GNAME75948(G75948,G81016,G75405);
  nand GNAME75949(G75949,G75948,G75947);
  or GNAME75950(G75950,G81035,G77788);
  or GNAME75951(G75951,G81017,G75412);
  nand GNAME75952(G75952,G75951,G75950);
  or GNAME75953(G75953,G81033,G75611);
  or GNAME75954(G75954,G81015,G75616);
  nand GNAME75955(G75955,G75954,G75953);
  or GNAME75956(G75956,G75641,G81018);
  or GNAME75957(G75957,G81012,G75692);
  nand GNAME75958(G75958,G75957,G75956);
  or GNAME75959(G75959,G81034,G75623);
  or GNAME75960(G75960,G81016,G75635);
  nand GNAME75961(G75961,G75960,G75959);
  or GNAME75962(G75962,G75642,G81019);
  or GNAME75963(G75963,G81013,G75695);
  nand GNAME75964(G75964,G75963,G75962);
  or GNAME75965(G75965,G81035,G75630);
  or GNAME75966(G75966,G81017,G75640);
  nand GNAME75967(G75967,G75966,G75965);
  or GNAME75968(G75968,G75643,G81020);
  or GNAME75969(G75969,G81014,G75697);
  nand GNAME75970(G75970,G75969,G75968);
  or GNAME75971(G75971,G81028,G75655);
  or GNAME75972(G75972,G81024,G75659);
  nand GNAME75973(G75973,G75972,G75971);
  or GNAME75974(G75974,G75693,G81018);
  or GNAME75975(G75975,G81012,G75694);
  nand GNAME75976(G75976,G75975,G75974);
  or GNAME75977(G75977,G81030,G75668);
  or GNAME75978(G75978,G81025,G75678);
  nand GNAME75979(G75979,G75978,G75977);
  or GNAME75980(G75980,G75696,G81019);
  or GNAME75981(G75981,G81013,G75699);
  nand GNAME75982(G75982,G75981,G75980);
  or GNAME75983(G75983,G81032,G75674);
  or GNAME75984(G75984,G81026,G75685);
  nand GNAME75985(G75985,G75984,G75983);
  or GNAME75986(G75986,G75698,G81020);
  or GNAME75987(G75987,G81014,G75700);
  nand GNAME75988(G75988,G75987,G75986);
  or GNAME75989(G75989,G80991,G75661);
  or GNAME75990(G75990,G81043,G75644);
  nand GNAME75991(G75991,G75990,G75989);
  or GNAME75992(G75992,G75694,G81018);
  or GNAME75993(G75993,G81021,G75737);
  nand GNAME75994(G75994,G75993,G75992);
  or GNAME75995(G75995,G80992,G75680);
  or GNAME75996(G75996,G81046,G75645);
  nand GNAME75997(G75997,G75996,G75995);
  or GNAME75998(G75998,G75699,G81019);
  or GNAME75999(G75999,G81022,G75739);
  nand GNAME76000(G76000,G75999,G75998);
  or GNAME76001(G76001,G80993,G75687);
  or GNAME76002(G76002,G81047,G75646);
  nand GNAME76003(G76003,G76002,G76001);
  or GNAME76004(G76004,G75700,G81020);
  or GNAME76005(G76005,G81023,G75741);
  nand GNAME76006(G76006,G76005,G76004);
  or GNAME76007(G76007,G80985,G75653);
  or GNAME76008(G76008,G81042,G75647);
  nand GNAME76009(G76009,G76008,G76007);
  or GNAME76010(G76010,G75692,G81018);
  or GNAME76011(G76011,G81012,G75693);
  nand GNAME76012(G76012,G76011,G76010);
  or GNAME76013(G76013,G80986,G75666);
  or GNAME76014(G76014,G81044,G75648);
  nand GNAME76015(G76015,G76014,G76013);
  or GNAME76016(G76016,G75695,G81019);
  or GNAME76017(G76017,G81013,G75696);
  nand GNAME76018(G76018,G76017,G76016);
  or GNAME76019(G76019,G80987,G75672);
  or GNAME76020(G76020,G81045,G75649);
  nand GNAME76021(G76021,G76020,G76019);
  or GNAME76022(G76022,G75697,G81020);
  or GNAME76023(G76023,G81014,G75698);
  nand GNAME76024(G76024,G76023,G76022);
  or GNAME76025(G76025,G81028,G75718);
  or GNAME76026(G76026,G81024,G75721);
  nand GNAME76027(G76027,G76026,G76025);
  or GNAME76028(G76028,G75737,G81009);
  or GNAME76029(G76029,G81021,G75738);
  nand GNAME76030(G76030,G76029,G76028);
  or GNAME76031(G76031,G81030,G75725);
  or GNAME76032(G76032,G81025,G75732);
  nand GNAME76033(G76033,G76032,G76031);
  or GNAME76034(G76034,G75739,G81010);
  or GNAME76035(G76035,G81022,G75740);
  nand GNAME76036(G76036,G76035,G76034);
  or GNAME76037(G76037,G81032,G75729);
  or GNAME76038(G76038,G81026,G75735);
  nand GNAME76039(G76039,G76038,G76037);
  or GNAME76040(G76040,G75741,G81011);
  or GNAME76041(G76041,G81023,G75742);
  nand GNAME76042(G76042,G76041,G76040);
  or GNAME76043(G76043,G81000,G75720);
  or GNAME76044(G76044,G81051,G75743);
  nand GNAME76045(G76045,G76044,G76043);
  or GNAME76046(G76046,G75738,G81009);
  or GNAME76047(G76047,G81021,G75776);
  nand GNAME76048(G76048,G76047,G76046);
  or GNAME76049(G76049,G81001,G75731);
  or GNAME76050(G76050,G81052,G75744);
  nand GNAME76051(G76051,G76050,G76049);
  or GNAME76052(G76052,G75740,G81010);
  or GNAME76053(G76053,G81022,G75780);
  nand GNAME76054(G76054,G76053,G76052);
  or GNAME76055(G76055,G81002,G75734);
  or GNAME76056(G76056,G81053,G75745);
  nand GNAME76057(G76057,G76056,G76055);
  or GNAME76058(G76058,G75742,G81011);
  or GNAME76059(G76059,G81023,G75782);
  nand GNAME76060(G76060,G76059,G76058);
  or GNAME76061(G76061,G81028,G75761);
  or GNAME76062(G76062,G81024,G75749);
  nand GNAME76063(G76063,G76062,G76061);
  or GNAME76064(G76064,G75776,G81009);
  or GNAME76065(G76065,G81021,G75777);
  nand GNAME76066(G76066,G76065,G76064);
  or GNAME76067(G76067,G81030,G75767);
  or GNAME76068(G76068,G81025,G75752);
  nand GNAME76069(G76069,G76068,G76067);
  or GNAME76070(G76070,G75780,G81010);
  or GNAME76071(G76071,G81022,G75781);
  nand GNAME76072(G76072,G76071,G76070);
  or GNAME76073(G76073,G81032,G75771);
  or GNAME76074(G76074,G81026,G75753);
  nand GNAME76075(G76075,G76074,G76073);
  or GNAME76076(G76076,G75782,G81011);
  or GNAME76077(G76077,G81023,G75783);
  nand GNAME76078(G76078,G76077,G76076);
  or GNAME76079(G76079,G81063,G75759);
  or GNAME76080(G76080,G81069,G75746);
  nand GNAME76081(G76081,G76080,G76079);
  or GNAME76082(G76082,G75777,G81009);
  or GNAME76083(G76083,G81021,G75778);
  nand GNAME76084(G76084,G76083,G76082);
  or GNAME76085(G76085,G81064,G75765);
  or GNAME76086(G76086,G81070,G75747);
  nand GNAME76087(G76087,G76086,G76085);
  or GNAME76088(G76088,G75781,G81010);
  or GNAME76089(G76089,G81022,G75784);
  nand GNAME76090(G76090,G76089,G76088);
  or GNAME76091(G76091,G81065,G75769);
  or GNAME76092(G76092,G81071,G75748);
  nand GNAME76093(G76093,G76092,G76091);
  or GNAME76094(G76094,G75783,G81011);
  or GNAME76095(G76095,G81023,G75786);
  nand GNAME76096(G76096,G76095,G76094);
  or GNAME76097(G76097,G81028,G75762);
  or GNAME76098(G76098,G81024,G75796);
  nand GNAME76099(G76099,G76098,G76097);
  or GNAME76100(G76100,G75778,G81009);
  or GNAME76101(G76101,G81021,G75779);
  nand GNAME76102(G76102,G76101,G76100);
  or GNAME76103(G76103,G81030,G75772);
  or GNAME76104(G76104,G81025,G75800);
  nand GNAME76105(G76105,G76104,G76103);
  or GNAME76106(G76106,G75784,G81010);
  or GNAME76107(G76107,G81022,G75785);
  nand GNAME76108(G76108,G76107,G76106);
  or GNAME76109(G76109,G81032,G75773);
  or GNAME76110(G76110,G81026,G75804);
  nand GNAME76111(G76111,G76110,G76109);
  or GNAME76112(G76112,G75786,G81011);
  or GNAME76113(G76113,G81023,G75787);
  nand GNAME76114(G76114,G76113,G76112);
  or GNAME76115(G76115,G81066,G75763);
  or GNAME76116(G76116,G81075,G75788);
  nand GNAME76117(G76117,G76116,G76115);
  or GNAME76118(G76118,G75779,G81009);
  or GNAME76119(G76119,G81021,G75813);
  nand GNAME76120(G76120,G76119,G76118);
  or GNAME76121(G76121,G81067,G75774);
  or GNAME76122(G76122,G81076,G75789);
  nand GNAME76123(G76123,G76122,G76121);
  or GNAME76124(G76124,G75785,G81010);
  or GNAME76125(G76125,G81022,G75814);
  nand GNAME76126(G76126,G76125,G76124);
  or GNAME76127(G76127,G81068,G75775);
  or GNAME76128(G76128,G81077,G75790);
  nand GNAME76129(G76129,G76128,G76127);
  or GNAME76130(G76130,G75787,G81011);
  or GNAME76131(G76131,G81023,G75815);
  nand GNAME76132(G76132,G76131,G76130);
  or GNAME76133(G76133,G81028,G75797);
  or GNAME76134(G76134,G81024,G75806);
  nand GNAME76135(G76135,G76134,G76133);
  or GNAME76136(G76136,G75813,G81009);
  or GNAME76137(G76137,G81021,G75812);
  nand GNAME76138(G76138,G76137,G76136);
  or GNAME76139(G76139,G81030,G75801);
  or GNAME76140(G76140,G81025,G75808);
  nand GNAME76141(G76141,G76140,G76139);
  or GNAME76142(G76142,G75814,G81010);
  or GNAME76143(G76143,G81022,G75816);
  nand GNAME76144(G76144,G76143,G76142);
  or GNAME76145(G76145,G81032,G75805);
  or GNAME76146(G76146,G81026,G75810);
  nand GNAME76147(G76147,G76146,G76145);
  or GNAME76148(G76148,G75815,G81011);
  or GNAME76149(G76149,G81023,G75817);
  nand GNAME76150(G76150,G76149,G76148);
  or GNAME76151(G76151,G81027,G75807);
  or GNAME76152(G76152,G81072,G75791);
  nand GNAME76153(G76153,G76152,G76151);
  or GNAME76154(G76154,G81078,G74169);
  or GNAME76155(G76155,G81060,G77786);
  nand GNAME76156(G76156,G76155,G76154);
  or GNAME76157(G76157,G81029,G75809);
  or GNAME76158(G76158,G81073,G75792);
  nand GNAME76159(G76159,G76158,G76157);
  or GNAME76160(G76160,G81079,G74172);
  or GNAME76161(G76161,G81061,G77783);
  nand GNAME76162(G76162,G76161,G76160);
  or GNAME76163(G76163,G81031,G75811);
  or GNAME76164(G76164,G81074,G75793);
  nand GNAME76165(G76165,G76164,G76163);
  or GNAME76166(G76166,G81080,G74175);
  or GNAME76167(G76167,G81062,G77784);
  nand GNAME76168(G76168,G76167,G76166);
  or GNAME76169(G76169,G81028,G75818);
  or GNAME76170(G76170,G81024,G75819);
  nand GNAME76171(G76171,G76170,G76169);
  or GNAME76172(G76172,G75824,G81009);
  or GNAME76173(G76173,G81021,G75825);
  nand GNAME76174(G76174,G76173,G76172);
  or GNAME76175(G76175,G81030,G75820);
  or GNAME76176(G76176,G81025,G75821);
  nand GNAME76177(G76177,G76176,G76175);
  or GNAME76178(G76178,G75826,G81010);
  or GNAME76179(G76179,G81022,G75827);
  nand GNAME76180(G76180,G76179,G76178);
  or GNAME76181(G76181,G81032,G75822);
  or GNAME76182(G76182,G81026,G75823);
  nand GNAME76183(G76183,G76182,G76181);
  or GNAME76184(G76184,G75828,G81011);
  or GNAME76185(G76185,G81023,G75829);
  nand GNAME76186(G76186,G76185,G76184);
  or GNAME76187(G76187,G75830,G81009);
  or GNAME76188(G76188,G81021,G75831);
  nand GNAME76189(G76189,G76188,G76187);
  or GNAME76190(G76190,G75832,G81010);
  or GNAME76191(G76191,G81022,G75833);
  nand GNAME76192(G76192,G76191,G76190);
  or GNAME76193(G76193,G75834,G81011);
  or GNAME76194(G76194,G81023,G75835);
  nand GNAME76195(G76195,G76194,G76193);
  or GNAME76196(G76196,G75831,G81009);
  or GNAME76197(G76197,G81021,G75836);
  nand GNAME76198(G76198,G76197,G76196);
  or GNAME76199(G76199,G75833,G81010);
  or GNAME76200(G76200,G81022,G75837);
  nand GNAME76201(G76201,G76200,G76199);
  or GNAME76202(G76202,G75835,G81011);
  or GNAME76203(G76203,G81023,G75838);
  nand GNAME76204(G76204,G76203,G76202);
  or GNAME76205(G76205,G74178,G81018);
  or GNAME76206(G76206,G81012,G77789);
  nand GNAME76207(G76207,G76206,G76205);
  or GNAME76208(G76208,G74181,G81019);
  or GNAME76209(G76209,G81013,G77790);
  nand GNAME76210(G76210,G76209,G76208);
  or GNAME76211(G76211,G74184,G81020);
  or GNAME76212(G76212,G81014,G77791);
  nand GNAME76213(G76213,G76212,G76211);
  or GNAME76214(G76214,G81028,G75819);
  or GNAME76215(G76215,G81024,G75839);
  nand GNAME76216(G76216,G76215,G76214);
  or GNAME76217(G76217,G81030,G75821);
  or GNAME76218(G76218,G81025,G75840);
  nand GNAME76219(G76219,G76218,G76217);
  or GNAME76220(G76220,G81032,G75823);
  or GNAME76221(G76221,G81026,G75841);
  nand GNAME76222(G76222,G76221,G76220);
  or GNAME76223(G76223,G81048,G77767);
  or GNAME76224(G76224,G80980,G75266);
  nand GNAME76225(G76225,G76224,G76223);
  or GNAME76226(G76226,G81049,G77766);
  or GNAME76227(G76227,G80981,G75268);
  nand GNAME76228(G76228,G76227,G76226);
  or GNAME76229(G76229,G81050,G77768);
  or GNAME76230(G76230,G80982,G75270);
  nand GNAME76231(G76231,G76230,G76229);
  or GNAME76232(G76232,G81054,G77769);
  or GNAME76233(G76233,G80988,G75273);
  nand GNAME76234(G76234,G76233,G76232);
  or GNAME76235(G76235,G81048,G75267);
  or GNAME76236(G76236,G80980,G75272);
  nand GNAME76237(G76237,G76236,G76235);
  or GNAME76238(G76238,G81055,G77770);
  or GNAME76239(G76239,G80989,G75277);
  nand GNAME76240(G76240,G76239,G76238);
  or GNAME76241(G76241,G81049,G75269);
  or GNAME76242(G76242,G80981,G75276);
  nand GNAME76243(G76243,G76242,G76241);
  or GNAME76244(G76244,G81056,G77771);
  or GNAME76245(G76245,G80990,G75281);
  nand GNAME76246(G76246,G76245,G76244);
  or GNAME76247(G76247,G81050,G75271);
  or GNAME76248(G76248,G80982,G75280);
  nand GNAME76249(G76249,G76248,G76247);
  or GNAME76250(G76250,G81048,G75272);
  or GNAME76251(G76251,G80980,G75275);
  nand GNAME76252(G76252,G76251,G76250);
  or GNAME76253(G76253,G81049,G75276);
  or GNAME76254(G76254,G80981,G75279);
  nand GNAME76255(G76255,G76254,G76253);
  or GNAME76256(G76256,G81050,G75280);
  or GNAME76257(G76257,G80982,G75283);
  nand GNAME76258(G76258,G76257,G76256);
  or GNAME76259(G76259,G81048,G75275);
  or GNAME76260(G76260,G80980,G75292);
  nand GNAME76261(G76261,G76260,G76259);
  or GNAME76262(G76262,G81049,G75279);
  or GNAME76263(G76263,G80981,G75297);
  nand GNAME76264(G76264,G76263,G76262);
  or GNAME76265(G76265,G81050,G75283);
  or GNAME76266(G76266,G80982,G75298);
  nand GNAME76267(G76267,G76266,G76265);
  or GNAME76268(G76268,G81003,G77774);
  or GNAME76269(G76269,G80994,G75291);
  nand GNAME76270(G76270,G76269,G76268);
  or GNAME76271(G76271,G81054,G75274);
  or GNAME76272(G76272,G80988,G75290);
  nand GNAME76273(G76273,G76272,G76271);
  or GNAME76274(G76274,G81005,G77776);
  or GNAME76275(G76275,G80996,G75294);
  nand GNAME76276(G76276,G76275,G76274);
  or GNAME76277(G76277,G81055,G75278);
  or GNAME76278(G76278,G80989,G75293);
  nand GNAME76279(G76279,G76278,G76277);
  or GNAME76280(G76280,G81006,G77777);
  or GNAME76281(G76281,G80997,G75296);
  nand GNAME76282(G76282,G76281,G76280);
  or GNAME76283(G76283,G81056,G75282);
  or GNAME76284(G76284,G80990,G75295);
  nand GNAME76285(G76285,G76284,G76283);
  or GNAME76286(G76286,G81048,G75292);
  or GNAME76287(G76287,G80980,G75284);
  nand GNAME76288(G76288,G76287,G76286);
  or GNAME76289(G76289,G81054,G75290);
  or GNAME76290(G76290,G80988,G75285);
  nand GNAME76291(G76291,G76290,G76289);
  or GNAME76292(G76292,G81049,G75297);
  or GNAME76293(G76293,G80981,G75286);
  nand GNAME76294(G76294,G76293,G76292);
  or GNAME76295(G76295,G81055,G75293);
  or GNAME76296(G76296,G80989,G75287);
  nand GNAME76297(G76297,G76296,G76295);
  or GNAME76298(G76298,G81050,G75298);
  or GNAME76299(G76299,G80982,G75288);
  nand GNAME76300(G76300,G76299,G76298);
  or GNAME76301(G76301,G81056,G75295);
  or GNAME76302(G76302,G80990,G75289);
  nand GNAME76303(G76303,G76302,G76301);
  or GNAME76304(G76304,G81004,G77775);
  or GNAME76305(G76305,G80995,G75301);
  nand GNAME76306(G76306,G76305,G76304);
  or GNAME76307(G76307,G81003,G75299);
  or GNAME76308(G76308,G80994,G75300);
  nand GNAME76309(G76309,G76308,G76307);
  or GNAME76310(G76310,G81007,G77778);
  or GNAME76311(G76311,G80998,G75306);
  nand GNAME76312(G76312,G76311,G76310);
  or GNAME76313(G76313,G81005,G75304);
  or GNAME76314(G76314,G80996,G75305);
  nand GNAME76315(G76315,G76314,G76313);
  or GNAME76316(G76316,G81008,G77779);
  or GNAME76317(G76317,G80999,G75309);
  nand GNAME76318(G76318,G76317,G76316);
  or GNAME76319(G76319,G81006,G75307);
  or GNAME76320(G76320,G80997,G75308);
  nand GNAME76321(G76321,G76320,G76319);
  or GNAME76322(G76322,G81054,G75285);
  or GNAME76323(G76323,G80988,G75303);
  nand GNAME76324(G76324,G76323,G76322);
  or GNAME76325(G76325,G81048,G75284);
  or GNAME76326(G76326,G80980,G75302);
  nand GNAME76327(G76327,G76326,G76325);
  or GNAME76328(G76328,G81055,G75287);
  or GNAME76329(G76329,G80989,G75311);
  nand GNAME76330(G76330,G76329,G76328);
  or GNAME76331(G76331,G81049,G75286);
  or GNAME76332(G76332,G80981,G75310);
  nand GNAME76333(G76333,G76332,G76331);
  or GNAME76334(G76334,G81056,G75289);
  or GNAME76335(G76335,G80990,G75313);
  nand GNAME76336(G76336,G76335,G76334);
  or GNAME76337(G76337,G81050,G75288);
  or GNAME76338(G76338,G80982,G75312);
  nand GNAME76339(G76339,G76338,G76337);
  or GNAME76340(G76340,G81081,G77780);
  or GNAME76341(G76341,G81057,G75318);
  nand GNAME76342(G76342,G76341,G76340);
  or GNAME76343(G76343,G81004,G75331);
  or GNAME76344(G76344,G80995,G75332);
  nand GNAME76345(G76345,G76344,G76343);
  or GNAME76346(G76346,G81082,G77781);
  or GNAME76347(G76347,G81058,G75326);
  nand GNAME76348(G76348,G76347,G76346);
  or GNAME76349(G76349,G81007,G75335);
  or GNAME76350(G76350,G80998,G75336);
  nand GNAME76351(G76351,G76350,G76349);
  or GNAME76352(G76352,G81083,G77782);
  or GNAME76353(G76353,G81059,G75328);
  nand GNAME76354(G76354,G76353,G76352);
  or GNAME76355(G76355,G81008,G75339);
  or GNAME76356(G76356,G80999,G75340);
  nand GNAME76357(G76357,G76356,G76355);
  or GNAME76358(G76358,G81004,G75301);
  or GNAME76359(G76359,G80995,G75331);
  nand GNAME76360(G76360,G76359,G76358);
  or GNAME76361(G76361,G81007,G75306);
  or GNAME76362(G76362,G80998,G75335);
  nand GNAME76363(G76363,G76362,G76361);
  or GNAME76364(G76364,G81008,G75309);
  or GNAME76365(G76365,G80999,G75339);
  nand GNAME76366(G76366,G76365,G76364);
  or GNAME76367(G76367,G81048,G75315);
  or GNAME76368(G76368,G80980,G75330);
  nand GNAME76369(G76369,G76368,G76367);
  or GNAME76370(G76370,G81054,G75316);
  or GNAME76371(G76371,G80988,G75317);
  nand GNAME76372(G76372,G76371,G76370);
  or GNAME76373(G76373,G81003,G75314);
  or GNAME76374(G76374,G80994,G75329);
  nand GNAME76375(G76375,G76374,G76373);
  or GNAME76376(G76376,G81049,G75320);
  or GNAME76377(G76377,G80981,G75334);
  nand GNAME76378(G76378,G76377,G76376);
  or GNAME76379(G76379,G81055,G75321);
  or GNAME76380(G76380,G80989,G75325);
  nand GNAME76381(G76381,G76380,G76379);
  or GNAME76382(G76382,G81005,G75319);
  or GNAME76383(G76383,G80996,G75333);
  nand GNAME76384(G76384,G76383,G76382);
  or GNAME76385(G76385,G81050,G75323);
  or GNAME76386(G76386,G80982,G75338);
  nand GNAME76387(G76387,G76386,G76385);
  or GNAME76388(G76388,G81056,G75324);
  or GNAME76389(G76389,G80990,G75327);
  nand GNAME76390(G76390,G76389,G76388);
  or GNAME76391(G76391,G81006,G75322);
  or GNAME76392(G76392,G80997,G75337);
  nand GNAME76393(G76393,G76392,G76391);
  or GNAME76394(G76394,G81054,G75303);
  or GNAME76395(G76395,G80988,G75316);
  nand GNAME76396(G76396,G76395,G76394);
  or GNAME76397(G76397,G81048,G75302);
  or GNAME76398(G76398,G80980,G75315);
  nand GNAME76399(G76399,G76398,G76397);
  or GNAME76400(G76400,G81055,G75311);
  or GNAME76401(G76401,G80989,G75321);
  nand GNAME76402(G76402,G76401,G76400);
  or GNAME76403(G76403,G81049,G75310);
  or GNAME76404(G76404,G80981,G75320);
  nand GNAME76405(G76405,G76404,G76403);
  or GNAME76406(G76406,G81056,G75313);
  or GNAME76407(G76407,G80990,G75324);
  nand GNAME76408(G76408,G76407,G76406);
  or GNAME76409(G76409,G81050,G75312);
  or GNAME76410(G76410,G80982,G75323);
  nand GNAME76411(G76411,G76410,G76409);
  or GNAME76412(G76412,G81003,G75329);
  or GNAME76413(G76413,G80994,G75346);
  nand GNAME76414(G76414,G76413,G76412);
  or GNAME76415(G76415,G81048,G75330);
  or GNAME76416(G76416,G80980,G75345);
  nand GNAME76417(G76417,G76416,G76415);
  or GNAME76418(G76418,G81005,G75333);
  or GNAME76419(G76419,G80996,G75356);
  nand GNAME76420(G76420,G76419,G76418);
  or GNAME76421(G76421,G81049,G75334);
  or GNAME76422(G76422,G80981,G75355);
  nand GNAME76423(G76423,G76422,G76421);
  or GNAME76424(G76424,G81006,G75337);
  or GNAME76425(G76425,G80997,G75359);
  nand GNAME76426(G76426,G76425,G76424);
  or GNAME76427(G76427,G81050,G75338);
  or GNAME76428(G76428,G80982,G75358);
  nand GNAME76429(G76429,G76428,G76427);
  or GNAME76430(G76430,G81081,G75318);
  or GNAME76431(G76431,G81057,G75347);
  nand GNAME76432(G76432,G76431,G76430);
  or GNAME76433(G76433,G81054,G75317);
  or GNAME76434(G76434,G80988,G75341);
  nand GNAME76435(G76435,G76434,G76433);
  or GNAME76436(G76436,G81082,G75326);
  or GNAME76437(G76437,G81058,G75360);
  nand GNAME76438(G76438,G76437,G76436);
  or GNAME76439(G76439,G81055,G75325);
  or GNAME76440(G76440,G80989,G75342);
  nand GNAME76441(G76441,G76440,G76439);
  or GNAME76442(G76442,G81083,G75328);
  or GNAME76443(G76443,G81059,G75367);
  nand GNAME76444(G76444,G76443,G76442);
  or GNAME76445(G76445,G81056,G75327);
  or GNAME76446(G76446,G80990,G75343);
  nand GNAME76447(G76447,G76446,G76445);
  or GNAME76448(G76448,G81078,G77786);
  or GNAME76449(G76449,G81060,G75349);
  nand GNAME76450(G76450,G76449,G76448);
  or GNAME76451(G76451,G81081,G75347);
  or GNAME76452(G76452,G81057,G75348);
  nand GNAME76453(G76453,G76452,G76451);
  or GNAME76454(G76454,G81079,G77783);
  or GNAME76455(G76455,G81061,G75362);
  nand GNAME76456(G76456,G76455,G76454);
  or GNAME76457(G76457,G81082,G75360);
  or GNAME76458(G76458,G81058,G75361);
  nand GNAME76459(G76459,G76458,G76457);
  or GNAME76460(G76460,G81080,G77784);
  or GNAME76461(G76461,G81062,G75369);
  nand GNAME76462(G76462,G76461,G76460);
  or GNAME76463(G76463,G81083,G75367);
  or GNAME76464(G76464,G81059,G75368);
  nand GNAME76465(G76465,G76464,G76463);
  or GNAME76466(G76466,G81004,G75344);
  or GNAME76467(G76467,G80995,G75352);
  nand GNAME76468(G76468,G76467,G76466);
  or GNAME76469(G76469,G81048,G75345);
  or GNAME76470(G76470,G80980,G75351);
  nand GNAME76471(G76471,G76470,G76469);
  or GNAME76472(G76472,G81003,G75346);
  or GNAME76473(G76473,G80994,G75350);
  nand GNAME76474(G76474,G76473,G76472);
  or GNAME76475(G76475,G81007,G75354);
  or GNAME76476(G76476,G80998,G75365);
  nand GNAME76477(G76477,G76476,G76475);
  or GNAME76478(G76478,G81049,G75355);
  or GNAME76479(G76479,G80981,G75364);
  nand GNAME76480(G76480,G76479,G76478);
  or GNAME76481(G76481,G81005,G75356);
  or GNAME76482(G76482,G80996,G75363);
  nand GNAME76483(G76483,G76482,G76481);
  or GNAME76484(G76484,G81008,G75357);
  or GNAME76485(G76485,G80999,G75372);
  nand GNAME76486(G76486,G76485,G76484);
  or GNAME76487(G76487,G81050,G75358);
  or GNAME76488(G76488,G80982,G75371);
  nand GNAME76489(G76489,G76488,G76487);
  or GNAME76490(G76490,G81006,G75359);
  or GNAME76491(G76491,G80997,G75370);
  nand GNAME76492(G76492,G76491,G76490);
  or GNAME76493(G76493,G81003,G75350);
  or GNAME76494(G76494,G80994,G75379);
  nand GNAME76495(G76495,G76494,G76493);
  or GNAME76496(G76496,G81054,G75353);
  or GNAME76497(G76497,G80988,G75378);
  nand GNAME76498(G76498,G76497,G76496);
  or GNAME76499(G76499,G81005,G75363);
  or GNAME76500(G76500,G80996,G75392);
  nand GNAME76501(G76501,G76500,G76499);
  or GNAME76502(G76502,G81055,G75366);
  or GNAME76503(G76503,G80989,G75391);
  nand GNAME76504(G76504,G76503,G76502);
  or GNAME76505(G76505,G81006,G75370);
  or GNAME76506(G76506,G80997,G75398);
  nand GNAME76507(G76507,G76506,G76505);
  or GNAME76508(G76508,G81056,G75373);
  or GNAME76509(G76509,G80990,G75397);
  nand GNAME76510(G76510,G76509,G76508);
  or GNAME76511(G76511,G81054,G75341);
  or GNAME76512(G76512,G80988,G75353);
  nand GNAME76513(G76513,G76512,G76511);
  or GNAME76514(G76514,G81055,G75342);
  or GNAME76515(G76515,G80989,G75366);
  nand GNAME76516(G76516,G76515,G76514);
  or GNAME76517(G76517,G81056,G75343);
  or GNAME76518(G76518,G80990,G75373);
  nand GNAME76519(G76519,G76518,G76517);
  or GNAME76520(G76520,G81078,G75349);
  or GNAME76521(G76521,G81060,G75376);
  nand GNAME76522(G76522,G76521,G76520);
  or GNAME76523(G76523,G81048,G75351);
  or GNAME76524(G76524,G81042,G75375);
  nand GNAME76525(G76525,G76524,G76523);
  or GNAME76526(G76526,G81081,G75348);
  or GNAME76527(G76527,G81057,G75374);
  nand GNAME76528(G76528,G76527,G76526);
  or GNAME76529(G76529,G81081,G75374);
  or GNAME76530(G76530,G81057,G75382);
  nand GNAME76531(G76531,G76530,G76529);
  or GNAME76532(G76532,G81003,G75379);
  or GNAME76533(G76533,G80994,G75381);
  nand GNAME76534(G76534,G76533,G76532);
  or GNAME76535(G76535,G81004,G75377);
  or GNAME76536(G76536,G80995,G75380);
  nand GNAME76537(G76537,G76536,G76535);
  or GNAME76538(G76538,G81079,G75362);
  or GNAME76539(G76539,G81061,G75389);
  nand GNAME76540(G76540,G76539,G76538);
  or GNAME76541(G76541,G81049,G75364);
  or GNAME76542(G76542,G81044,G75388);
  nand GNAME76543(G76543,G76542,G76541);
  or GNAME76544(G76544,G81082,G75361);
  or GNAME76545(G76545,G81058,G75387);
  nand GNAME76546(G76546,G76545,G76544);
  or GNAME76547(G76547,G81080,G75369);
  or GNAME76548(G76548,G81062,G75395);
  nand GNAME76549(G76549,G76548,G76547);
  or GNAME76550(G76550,G81050,G75371);
  or GNAME76551(G76551,G81045,G75394);
  nand GNAME76552(G76552,G76551,G76550);
  or GNAME76553(G76553,G81083,G75368);
  or GNAME76554(G76554,G81059,G75393);
  nand GNAME76555(G76555,G76554,G76553);
  or GNAME76556(G76556,G81082,G75387);
  or GNAME76557(G76557,G81058,G75401);
  nand GNAME76558(G76558,G76557,G76556);
  or GNAME76559(G76559,G81005,G75392);
  or GNAME76560(G76560,G80996,G75400);
  nand GNAME76561(G76561,G76560,G76559);
  or GNAME76562(G76562,G81007,G75390);
  or GNAME76563(G76563,G80998,G75399);
  nand GNAME76564(G76564,G76563,G76562);
  or GNAME76565(G76565,G81083,G75393);
  or GNAME76566(G76566,G81059,G75408);
  nand GNAME76567(G76567,G76566,G76565);
  or GNAME76568(G76568,G81006,G75398);
  or GNAME76569(G76569,G80997,G75407);
  nand GNAME76570(G76570,G76569,G76568);
  or GNAME76571(G76571,G81008,G75396);
  or GNAME76572(G76572,G80999,G75406);
  nand GNAME76573(G76573,G76572,G76571);
  or GNAME76574(G76574,G81078,G75376);
  or GNAME76575(G76575,G81060,G75385);
  nand GNAME76576(G76576,G76575,G76574);
  or GNAME76577(G76577,G80985,G75375);
  or GNAME76578(G76578,G81042,G75384);
  nand GNAME76579(G76579,G76578,G76577);
  or GNAME76580(G76580,G81054,G75378);
  or GNAME76581(G76581,G80988,G75383);
  nand GNAME76582(G76582,G76581,G76580);
  or GNAME76583(G76583,G81079,G75389);
  or GNAME76584(G76584,G81061,G75404);
  nand GNAME76585(G76585,G76584,G76583);
  or GNAME76586(G76586,G80986,G75388);
  or GNAME76587(G76587,G81044,G75403);
  nand GNAME76588(G76588,G76587,G76586);
  or GNAME76589(G76589,G81055,G75391);
  or GNAME76590(G76590,G80989,G75402);
  nand GNAME76591(G76591,G76590,G76589);
  or GNAME76592(G76592,G81080,G75395);
  or GNAME76593(G76593,G81062,G75411);
  nand GNAME76594(G76594,G76593,G76592);
  or GNAME76595(G76595,G80987,G75394);
  or GNAME76596(G76596,G81045,G75410);
  nand GNAME76597(G76597,G76596,G76595);
  or GNAME76598(G76598,G81056,G75397);
  or GNAME76599(G76599,G80990,G75409);
  nand GNAME76600(G76600,G76599,G76598);
  or GNAME76601(G76601,G81004,G75380);
  or GNAME76602(G76602,G80995,G75414);
  nand GNAME76603(G76603,G76602,G76601);
  or GNAME76604(G76604,G80985,G75384);
  or GNAME76605(G76605,G81042,G75413);
  nand GNAME76606(G76606,G76605,G76604);
  or GNAME76607(G76607,G81007,G75399);
  or GNAME76608(G76608,G80998,G75428);
  nand GNAME76609(G76609,G76608,G76607);
  or GNAME76610(G76610,G80986,G75403);
  or GNAME76611(G76611,G81044,G75427);
  nand GNAME76612(G76612,G76611,G76610);
  or GNAME76613(G76613,G81008,G75406);
  or GNAME76614(G76614,G80999,G75435);
  nand GNAME76615(G76615,G76614,G76613);
  or GNAME76616(G76616,G80987,G75410);
  or GNAME76617(G76617,G81045,G75434);
  nand GNAME76618(G76618,G76617,G76616);
  or GNAME76619(G76619,G81081,G75418);
  or GNAME76620(G76620,G81057,G75422);
  nand GNAME76621(G76621,G76620,G76619);
  or GNAME76622(G76622,G81003,G75416);
  or GNAME76623(G76623,G80994,G75421);
  nand GNAME76624(G76624,G76623,G76622);
  or GNAME76625(G76625,G81004,G75414);
  or GNAME76626(G76626,G80995,G75420);
  nand GNAME76627(G76627,G76626,G76625);
  or GNAME76628(G76628,G81082,G75432);
  or GNAME76629(G76629,G81058,G75443);
  nand GNAME76630(G76630,G76629,G76628);
  or GNAME76631(G76631,G81005,G75430);
  or GNAME76632(G76632,G80996,G75442);
  nand GNAME76633(G76633,G76632,G76631);
  or GNAME76634(G76634,G81007,G75428);
  or GNAME76635(G76635,G80998,G75441);
  nand GNAME76636(G76636,G76635,G76634);
  or GNAME76637(G76637,G81083,G75439);
  or GNAME76638(G76638,G81059,G75450);
  nand GNAME76639(G76639,G76638,G76637);
  or GNAME76640(G76640,G81006,G75437);
  or GNAME76641(G76641,G80997,G75449);
  nand GNAME76642(G76642,G76641,G76640);
  or GNAME76643(G76643,G81008,G75435);
  or GNAME76644(G76644,G80999,G75448);
  nand GNAME76645(G76645,G76644,G76643);
  or GNAME76646(G76646,G81033,G75417);
  or GNAME76647(G76647,G81015,G75426);
  nand GNAME76648(G76648,G76647,G76646);
  or GNAME76649(G76649,G77789,G81018);
  or GNAME76650(G76650,G81012,G75455);
  nand GNAME76651(G76651,G76650,G76649);
  or GNAME76652(G76652,G81034,G75431);
  or GNAME76653(G76653,G81016,G75447);
  nand GNAME76654(G76654,G76653,G76652);
  or GNAME76655(G76655,G77790,G81019);
  or GNAME76656(G76656,G81013,G75456);
  nand GNAME76657(G76657,G76656,G76655);
  or GNAME76658(G76658,G81035,G75438);
  or GNAME76659(G76659,G81017,G75454);
  nand GNAME76660(G76660,G76659,G76658);
  or GNAME76661(G76661,G77791,G81020);
  or GNAME76662(G76662,G81014,G75457);
  nand GNAME76663(G76663,G76662,G76661);
  or GNAME76664(G76664,G81054,G75383);
  or GNAME76665(G76665,G81043,G75419);
  nand GNAME76666(G76666,G76665,G76664);
  or GNAME76667(G76667,G81081,G75382);
  or GNAME76668(G76668,G81057,G75418);
  nand GNAME76669(G76669,G76668,G76667);
  or GNAME76670(G76670,G81055,G75402);
  or GNAME76671(G76671,G81046,G75433);
  nand GNAME76672(G76672,G76671,G76670);
  or GNAME76673(G76673,G81082,G75401);
  or GNAME76674(G76674,G81058,G75432);
  nand GNAME76675(G76675,G76674,G76673);
  or GNAME76676(G76676,G81056,G75409);
  or GNAME76677(G76677,G81047,G75440);
  nand GNAME76678(G76678,G76677,G76676);
  or GNAME76679(G76679,G81083,G75408);
  or GNAME76680(G76680,G81059,G75439);
  nand GNAME76681(G76681,G76680,G76679);
  or GNAME76682(G76682,G81033,G75386);
  or GNAME76683(G76683,G81015,G75417);
  nand GNAME76684(G76684,G76683,G76682);
  or GNAME76685(G76685,G81003,G75381);
  or GNAME76686(G76686,G80994,G75416);
  nand GNAME76687(G76687,G76686,G76685);
  or GNAME76688(G76688,G81078,G75385);
  or GNAME76689(G76689,G81060,G75415);
  nand GNAME76690(G76690,G76689,G76688);
  or GNAME76691(G76691,G81078,G75415);
  or GNAME76692(G76692,G81060,G75425);
  nand GNAME76693(G76693,G76692,G76691);
  or GNAME76694(G76694,G80985,G75413);
  or GNAME76695(G76695,G81042,G75424);
  nand GNAME76696(G76696,G76695,G76694);
  or GNAME76697(G76697,G80991,G75419);
  or GNAME76698(G76698,G81043,G75423);
  nand GNAME76699(G76699,G76698,G76697);
  or GNAME76700(G76700,G81034,G75405);
  or GNAME76701(G76701,G81016,G75431);
  nand GNAME76702(G76702,G76701,G76700);
  or GNAME76703(G76703,G81005,G75400);
  or GNAME76704(G76704,G80996,G75430);
  nand GNAME76705(G76705,G76704,G76703);
  or GNAME76706(G76706,G81079,G75404);
  or GNAME76707(G76707,G81061,G75429);
  nand GNAME76708(G76708,G76707,G76706);
  or GNAME76709(G76709,G81035,G75412);
  or GNAME76710(G76710,G81017,G75438);
  nand GNAME76711(G76711,G76710,G76709);
  or GNAME76712(G76712,G81006,G75407);
  or GNAME76713(G76713,G80997,G75437);
  nand GNAME76714(G76714,G76713,G76712);
  or GNAME76715(G76715,G81080,G75411);
  or GNAME76716(G76716,G81062,G75436);
  nand GNAME76717(G76717,G76716,G76715);
  or GNAME76718(G76718,G81079,G75429);
  or GNAME76719(G76719,G81061,G75446);
  nand GNAME76720(G76720,G76719,G76718);
  or GNAME76721(G76721,G80986,G75427);
  or GNAME76722(G76722,G81044,G75445);
  nand GNAME76723(G76723,G76722,G76721);
  or GNAME76724(G76724,G80992,G75433);
  or GNAME76725(G76725,G81046,G75444);
  nand GNAME76726(G76726,G76725,G76724);
  or GNAME76727(G76727,G81080,G75436);
  or GNAME76728(G76728,G81062,G75453);
  nand GNAME76729(G76729,G76728,G76727);
  or GNAME76730(G76730,G80987,G75434);
  or GNAME76731(G76731,G81045,G75452);
  nand GNAME76732(G76732,G76731,G76730);
  or GNAME76733(G76733,G80993,G75440);
  or GNAME76734(G76734,G81047,G75451);
  nand GNAME76735(G76735,G76734,G76733);
  or GNAME76736(G76736,G81081,G75422);
  or GNAME76737(G76737,G81057,G75460);
  nand GNAME76738(G76738,G76737,G76736);
  or GNAME76739(G76739,G81003,G75421);
  or GNAME76740(G76740,G81051,G75459);
  nand GNAME76741(G76741,G76740,G76739);
  or GNAME76742(G76742,G81004,G75420);
  or GNAME76743(G76743,G80995,G75458);
  nand GNAME76744(G76744,G76743,G76742);
  or GNAME76745(G76745,G81081,G75460);
  or GNAME76746(G76746,G81057,G75467);
  nand GNAME76747(G76747,G76746,G76745);
  or GNAME76748(G76748,G81000,G75459);
  or GNAME76749(G76749,G81051,G75466);
  nand GNAME76750(G76750,G76749,G76748);
  or GNAME76751(G76751,G81004,G75458);
  or GNAME76752(G76752,G80995,G75465);
  nand GNAME76753(G76753,G76752,G76751);
  or GNAME76754(G76754,G81082,G75443);
  or GNAME76755(G76755,G81058,G75474);
  nand GNAME76756(G76756,G76755,G76754);
  or GNAME76757(G76757,G81005,G75442);
  or GNAME76758(G76758,G81052,G75473);
  nand GNAME76759(G76759,G76758,G76757);
  or GNAME76760(G76760,G81007,G75441);
  or GNAME76761(G76761,G80998,G75472);
  nand GNAME76762(G76762,G76761,G76760);
  or GNAME76763(G76763,G81083,G75450);
  or GNAME76764(G76764,G81059,G75481);
  nand GNAME76765(G76765,G76764,G76763);
  or GNAME76766(G76766,G81006,G75449);
  or GNAME76767(G76767,G81053,G75480);
  nand GNAME76768(G76768,G76767,G76766);
  or GNAME76769(G76769,G81008,G75448);
  or GNAME76770(G76770,G80999,G75479);
  nand GNAME76771(G76771,G76770,G76769);
  or GNAME76772(G76772,G81082,G75474);
  or GNAME76773(G76773,G81058,G75488);
  nand GNAME76774(G76774,G76773,G76772);
  or GNAME76775(G76775,G81001,G75473);
  or GNAME76776(G76776,G81052,G75487);
  nand GNAME76777(G76777,G76776,G76775);
  or GNAME76778(G76778,G81007,G75472);
  or GNAME76779(G76779,G80998,G75486);
  nand GNAME76780(G76780,G76779,G76778);
  or GNAME76781(G76781,G81083,G75481);
  or GNAME76782(G76782,G81059,G75495);
  nand GNAME76783(G76783,G76782,G76781);
  or GNAME76784(G76784,G81002,G75480);
  or GNAME76785(G76785,G81053,G75494);
  nand GNAME76786(G76786,G76785,G76784);
  or GNAME76787(G76787,G81008,G75479);
  or GNAME76788(G76788,G80999,G75493);
  nand GNAME76789(G76789,G76788,G76787);
  or GNAME76790(G76790,G81033,G75426);
  or GNAME76791(G76791,G81015,G75464);
  nand GNAME76792(G76792,G76791,G76790);
  or GNAME76793(G76793,G75455,G81018);
  or GNAME76794(G76794,G81012,G75500);
  nand GNAME76795(G76795,G76794,G76793);
  or GNAME76796(G76796,G81033,G75464);
  or GNAME76797(G76797,G81015,G75471);
  nand GNAME76798(G76798,G76797,G76796);
  or GNAME76799(G76799,G75500,G81018);
  or GNAME76800(G76800,G81012,G75501);
  nand GNAME76801(G76801,G76800,G76799);
  or GNAME76802(G76802,G81034,G75447);
  or GNAME76803(G76803,G81016,G75478);
  nand GNAME76804(G76804,G76803,G76802);
  or GNAME76805(G76805,G75456,G81019);
  or GNAME76806(G76806,G81013,G75502);
  nand GNAME76807(G76807,G76806,G76805);
  or GNAME76808(G76808,G81035,G75454);
  or GNAME76809(G76809,G81017,G75485);
  nand GNAME76810(G76810,G76809,G76808);
  or GNAME76811(G76811,G75457,G81020);
  or GNAME76812(G76812,G81014,G75503);
  nand GNAME76813(G76813,G76812,G76811);
  or GNAME76814(G76814,G81034,G75478);
  or GNAME76815(G76815,G81016,G75492);
  nand GNAME76816(G76816,G76815,G76814);
  or GNAME76817(G76817,G75502,G81019);
  or GNAME76818(G76818,G81013,G75504);
  nand GNAME76819(G76819,G76818,G76817);
  or GNAME76820(G76820,G81035,G75485);
  or GNAME76821(G76821,G81017,G75499);
  nand GNAME76822(G76822,G76821,G76820);
  or GNAME76823(G76823,G75503,G81020);
  or GNAME76824(G76824,G81014,G75505);
  nand GNAME76825(G76825,G76824,G76823);
  or GNAME76826(G76826,G81078,G75425);
  or GNAME76827(G76827,G81060,G75463);
  nand GNAME76828(G76828,G76827,G76826);
  or GNAME76829(G76829,G80985,G75424);
  or GNAME76830(G76830,G81042,G75462);
  nand GNAME76831(G76831,G76830,G76829);
  or GNAME76832(G76832,G80991,G75423);
  or GNAME76833(G76833,G81043,G75461);
  nand GNAME76834(G76834,G76833,G76832);
  or GNAME76835(G76835,G81078,G75463);
  or GNAME76836(G76836,G81060,G75470);
  nand GNAME76837(G76837,G76836,G76835);
  or GNAME76838(G76838,G80985,G75462);
  or GNAME76839(G76839,G81042,G75469);
  nand GNAME76840(G76840,G76839,G76838);
  or GNAME76841(G76841,G80991,G75461);
  or GNAME76842(G76842,G81043,G75468);
  nand GNAME76843(G76843,G76842,G76841);
  or GNAME76844(G76844,G81079,G75446);
  or GNAME76845(G76845,G81061,G75477);
  nand GNAME76846(G76846,G76845,G76844);
  or GNAME76847(G76847,G80986,G75445);
  or GNAME76848(G76848,G81044,G75476);
  nand GNAME76849(G76849,G76848,G76847);
  or GNAME76850(G76850,G80992,G75444);
  or GNAME76851(G76851,G81046,G75475);
  nand GNAME76852(G76852,G76851,G76850);
  or GNAME76853(G76853,G81080,G75453);
  or GNAME76854(G76854,G81062,G75484);
  nand GNAME76855(G76855,G76854,G76853);
  or GNAME76856(G76856,G80987,G75452);
  or GNAME76857(G76857,G81045,G75483);
  nand GNAME76858(G76858,G76857,G76856);
  or GNAME76859(G76859,G80993,G75451);
  or GNAME76860(G76860,G81047,G75482);
  nand GNAME76861(G76861,G76860,G76859);
  or GNAME76862(G76862,G81079,G75477);
  or GNAME76863(G76863,G81061,G75491);
  nand GNAME76864(G76864,G76863,G76862);
  or GNAME76865(G76865,G80986,G75476);
  or GNAME76866(G76866,G81044,G75490);
  nand GNAME76867(G76867,G76866,G76865);
  or GNAME76868(G76868,G80992,G75475);
  or GNAME76869(G76869,G81046,G75489);
  nand GNAME76870(G76870,G76869,G76868);
  or GNAME76871(G76871,G81080,G75484);
  or GNAME76872(G76872,G81062,G75498);
  nand GNAME76873(G76873,G76872,G76871);
  or GNAME76874(G76874,G80987,G75483);
  or GNAME76875(G76875,G81045,G75497);
  nand GNAME76876(G76876,G76875,G76874);
  or GNAME76877(G76877,G80993,G75482);
  or GNAME76878(G76878,G81047,G75496);
  nand GNAME76879(G76879,G76878,G76877);
  or GNAME76880(G76880,G81081,G75467);
  or GNAME76881(G76881,G81057,G75508);
  nand GNAME76882(G76882,G76881,G76880);
  or GNAME76883(G76883,G81000,G75466);
  or GNAME76884(G76884,G81051,G75507);
  nand GNAME76885(G76885,G76884,G76883);
  or GNAME76886(G76886,G81004,G75465);
  or GNAME76887(G76887,G81069,G75506);
  nand GNAME76888(G76888,G76887,G76886);
  or GNAME76889(G76889,G81081,G75508);
  or GNAME76890(G76890,G81057,G75515);
  nand GNAME76891(G76891,G76890,G76889);
  or GNAME76892(G76892,G81000,G75507);
  or GNAME76893(G76893,G81051,G75514);
  nand GNAME76894(G76894,G76893,G76892);
  or GNAME76895(G76895,G81063,G75506);
  or GNAME76896(G76896,G81069,G75513);
  nand GNAME76897(G76897,G76896,G76895);
  or GNAME76898(G76898,G81082,G75488);
  or GNAME76899(G76899,G81058,G75522);
  nand GNAME76900(G76900,G76899,G76898);
  or GNAME76901(G76901,G81001,G75487);
  or GNAME76902(G76902,G81052,G75521);
  nand GNAME76903(G76903,G76902,G76901);
  or GNAME76904(G76904,G81007,G75486);
  or GNAME76905(G76905,G81070,G75520);
  nand GNAME76906(G76906,G76905,G76904);
  or GNAME76907(G76907,G81083,G75495);
  or GNAME76908(G76908,G81059,G75529);
  nand GNAME76909(G76909,G76908,G76907);
  or GNAME76910(G76910,G81002,G75494);
  or GNAME76911(G76911,G81053,G75528);
  nand GNAME76912(G76912,G76911,G76910);
  or GNAME76913(G76913,G81008,G75493);
  or GNAME76914(G76914,G81071,G75527);
  nand GNAME76915(G76915,G76914,G76913);
  or GNAME76916(G76916,G81082,G75522);
  or GNAME76917(G76917,G81058,G75536);
  nand GNAME76918(G76918,G76917,G76916);
  or GNAME76919(G76919,G81001,G75521);
  or GNAME76920(G76920,G81052,G75535);
  nand GNAME76921(G76921,G76920,G76919);
  or GNAME76922(G76922,G81064,G75520);
  or GNAME76923(G76923,G81070,G75534);
  nand GNAME76924(G76924,G76923,G76922);
  or GNAME76925(G76925,G81083,G75529);
  or GNAME76926(G76926,G81059,G75543);
  nand GNAME76927(G76927,G76926,G76925);
  or GNAME76928(G76928,G81002,G75528);
  or GNAME76929(G76929,G81053,G75542);
  nand GNAME76930(G76930,G76929,G76928);
  or GNAME76931(G76931,G81065,G75527);
  or GNAME76932(G76932,G81071,G75541);
  nand GNAME76933(G76933,G76932,G76931);
  or GNAME76934(G76934,G81033,G75471);
  or GNAME76935(G76935,G81015,G75512);
  nand GNAME76936(G76936,G76935,G76934);
  or GNAME76937(G76937,G75501,G81018);
  or GNAME76938(G76938,G81012,G75548);
  nand GNAME76939(G76939,G76938,G76937);
  or GNAME76940(G76940,G81033,G75512);
  or GNAME76941(G76941,G81015,G75519);
  nand GNAME76942(G76942,G76941,G76940);
  or GNAME76943(G76943,G75548,G81018);
  or GNAME76944(G76944,G81012,G75549);
  nand GNAME76945(G76945,G76944,G76943);
  or GNAME76946(G76946,G81034,G75492);
  or GNAME76947(G76947,G81016,G75526);
  nand GNAME76948(G76948,G76947,G76946);
  or GNAME76949(G76949,G75504,G81019);
  or GNAME76950(G76950,G81013,G75550);
  nand GNAME76951(G76951,G76950,G76949);
  or GNAME76952(G76952,G81035,G75499);
  or GNAME76953(G76953,G81017,G75533);
  nand GNAME76954(G76954,G76953,G76952);
  or GNAME76955(G76955,G75505,G81020);
  or GNAME76956(G76956,G81014,G75551);
  nand GNAME76957(G76957,G76956,G76955);
  or GNAME76958(G76958,G81034,G75526);
  or GNAME76959(G76959,G81016,G75540);
  nand GNAME76960(G76960,G76959,G76958);
  or GNAME76961(G76961,G75550,G81019);
  or GNAME76962(G76962,G81013,G75552);
  nand GNAME76963(G76963,G76962,G76961);
  or GNAME76964(G76964,G81035,G75533);
  or GNAME76965(G76965,G81017,G75547);
  nand GNAME76966(G76966,G76965,G76964);
  or GNAME76967(G76967,G75551,G81020);
  or GNAME76968(G76968,G81014,G75553);
  nand GNAME76969(G76969,G76968,G76967);
  or GNAME76970(G76970,G81078,G75470);
  or GNAME76971(G76971,G81060,G75511);
  nand GNAME76972(G76972,G76971,G76970);
  or GNAME76973(G76973,G80985,G75469);
  or GNAME76974(G76974,G81042,G75510);
  nand GNAME76975(G76975,G76974,G76973);
  or GNAME76976(G76976,G80991,G75468);
  or GNAME76977(G76977,G81043,G75509);
  nand GNAME76978(G76978,G76977,G76976);
  or GNAME76979(G76979,G81078,G75511);
  or GNAME76980(G76980,G81060,G75518);
  nand GNAME76981(G76981,G76980,G76979);
  or GNAME76982(G76982,G80985,G75510);
  or GNAME76983(G76983,G81042,G75517);
  nand GNAME76984(G76984,G76983,G76982);
  or GNAME76985(G76985,G80991,G75509);
  or GNAME76986(G76986,G81043,G75516);
  nand GNAME76987(G76987,G76986,G76985);
  or GNAME76988(G76988,G81079,G75491);
  or GNAME76989(G76989,G81061,G75525);
  nand GNAME76990(G76990,G76989,G76988);
  or GNAME76991(G76991,G80986,G75490);
  or GNAME76992(G76992,G81044,G75524);
  nand GNAME76993(G76993,G76992,G76991);
  or GNAME76994(G76994,G80992,G75489);
  or GNAME76995(G76995,G81046,G75523);
  nand GNAME76996(G76996,G76995,G76994);
  or GNAME76997(G76997,G81080,G75498);
  or GNAME76998(G76998,G81062,G75532);
  nand GNAME76999(G76999,G76998,G76997);
  or GNAME77000(G77000,G80987,G75497);
  or GNAME77001(G77001,G81045,G75531);
  nand GNAME77002(G77002,G77001,G77000);
  or GNAME77003(G77003,G80993,G75496);
  or GNAME77004(G77004,G81047,G75530);
  nand GNAME77005(G77005,G77004,G77003);
  or GNAME77006(G77006,G81079,G75525);
  or GNAME77007(G77007,G81061,G75539);
  nand GNAME77008(G77008,G77007,G77006);
  or GNAME77009(G77009,G80986,G75524);
  or GNAME77010(G77010,G81044,G75538);
  nand GNAME77011(G77011,G77010,G77009);
  or GNAME77012(G77012,G80992,G75523);
  or GNAME77013(G77013,G81046,G75537);
  nand GNAME77014(G77014,G77013,G77012);
  or GNAME77015(G77015,G81080,G75532);
  or GNAME77016(G77016,G81062,G75546);
  nand GNAME77017(G77017,G77016,G77015);
  or GNAME77018(G77018,G80987,G75531);
  or GNAME77019(G77019,G81045,G75545);
  nand GNAME77020(G77020,G77019,G77018);
  or GNAME77021(G77021,G80993,G75530);
  or GNAME77022(G77022,G81047,G75544);
  nand GNAME77023(G77023,G77022,G77021);
  or GNAME77024(G77024,G81081,G75515);
  or GNAME77025(G77025,G81075,G75556);
  nand GNAME77026(G77026,G77025,G77024);
  or GNAME77027(G77027,G81000,G75514);
  or GNAME77028(G77028,G81051,G75555);
  nand GNAME77029(G77029,G77028,G77027);
  or GNAME77030(G77030,G81063,G75513);
  or GNAME77031(G77031,G81069,G75554);
  nand GNAME77032(G77032,G77031,G77030);
  or GNAME77033(G77033,G81066,G75556);
  or GNAME77034(G77034,G81075,G75563);
  nand GNAME77035(G77035,G77034,G77033);
  or GNAME77036(G77036,G81000,G75555);
  or GNAME77037(G77037,G81051,G75562);
  nand GNAME77038(G77038,G77037,G77036);
  or GNAME77039(G77039,G81063,G75554);
  or GNAME77040(G77040,G81069,G75561);
  nand GNAME77041(G77041,G77040,G77039);
  or GNAME77042(G77042,G81082,G75536);
  or GNAME77043(G77043,G81076,G75570);
  nand GNAME77044(G77044,G77043,G77042);
  or GNAME77045(G77045,G81001,G75535);
  or GNAME77046(G77046,G81052,G75569);
  nand GNAME77047(G77047,G77046,G77045);
  or GNAME77048(G77048,G81064,G75534);
  or GNAME77049(G77049,G81070,G75568);
  nand GNAME77050(G77050,G77049,G77048);
  or GNAME77051(G77051,G81083,G75543);
  or GNAME77052(G77052,G81077,G75577);
  nand GNAME77053(G77053,G77052,G77051);
  or GNAME77054(G77054,G81002,G75542);
  or GNAME77055(G77055,G81053,G75576);
  nand GNAME77056(G77056,G77055,G77054);
  or GNAME77057(G77057,G81065,G75541);
  or GNAME77058(G77058,G81071,G75575);
  nand GNAME77059(G77059,G77058,G77057);
  or GNAME77060(G77060,G81067,G75570);
  or GNAME77061(G77061,G81076,G75584);
  nand GNAME77062(G77062,G77061,G77060);
  or GNAME77063(G77063,G81001,G75569);
  or GNAME77064(G77064,G81052,G75583);
  nand GNAME77065(G77065,G77064,G77063);
  or GNAME77066(G77066,G81064,G75568);
  or GNAME77067(G77067,G81070,G75582);
  nand GNAME77068(G77068,G77067,G77066);
  or GNAME77069(G77069,G81068,G75577);
  or GNAME77070(G77070,G81077,G75591);
  nand GNAME77071(G77071,G77070,G77069);
  or GNAME77072(G77072,G81002,G75576);
  or GNAME77073(G77073,G81053,G75590);
  nand GNAME77074(G77074,G77073,G77072);
  or GNAME77075(G77075,G81065,G75575);
  or GNAME77076(G77076,G81071,G75589);
  nand GNAME77077(G77077,G77076,G77075);
  or GNAME77078(G77078,G81033,G75519);
  or GNAME77079(G77079,G81015,G75560);
  nand GNAME77080(G77080,G77079,G77078);
  or GNAME77081(G77081,G75549,G81018);
  or GNAME77082(G77082,G81012,G75596);
  nand GNAME77083(G77083,G77082,G77081);
  or GNAME77084(G77084,G81033,G75560);
  or GNAME77085(G77085,G81015,G75567);
  nand GNAME77086(G77086,G77085,G77084);
  or GNAME77087(G77087,G75596,G81018);
  or GNAME77088(G77088,G81012,G75597);
  nand GNAME77089(G77089,G77088,G77087);
  or GNAME77090(G77090,G81034,G75540);
  or GNAME77091(G77091,G81016,G75574);
  nand GNAME77092(G77092,G77091,G77090);
  or GNAME77093(G77093,G75552,G81019);
  or GNAME77094(G77094,G81013,G75598);
  nand GNAME77095(G77095,G77094,G77093);
  or GNAME77096(G77096,G81035,G75547);
  or GNAME77097(G77097,G81017,G75581);
  nand GNAME77098(G77098,G77097,G77096);
  or GNAME77099(G77099,G75553,G81020);
  or GNAME77100(G77100,G81014,G75599);
  nand GNAME77101(G77101,G77100,G77099);
  or GNAME77102(G77102,G81034,G75574);
  or GNAME77103(G77103,G81016,G75588);
  nand GNAME77104(G77104,G77103,G77102);
  or GNAME77105(G77105,G75598,G81019);
  or GNAME77106(G77106,G81013,G75600);
  nand GNAME77107(G77107,G77106,G77105);
  or GNAME77108(G77108,G81035,G75581);
  or GNAME77109(G77109,G81017,G75595);
  nand GNAME77110(G77110,G77109,G77108);
  or GNAME77111(G77111,G75599,G81020);
  or GNAME77112(G77112,G81014,G75601);
  nand GNAME77113(G77113,G77112,G77111);
  or GNAME77114(G77114,G81078,G75518);
  or GNAME77115(G77115,G81060,G75559);
  nand GNAME77116(G77116,G77115,G77114);
  or GNAME77117(G77117,G80985,G75517);
  or GNAME77118(G77118,G81042,G75558);
  nand GNAME77119(G77119,G77118,G77117);
  or GNAME77120(G77120,G80991,G75516);
  or GNAME77121(G77121,G81043,G75557);
  nand GNAME77122(G77122,G77121,G77120);
  or GNAME77123(G77123,G81078,G75559);
  or GNAME77124(G77124,G81060,G75566);
  nand GNAME77125(G77125,G77124,G77123);
  or GNAME77126(G77126,G80985,G75558);
  or GNAME77127(G77127,G81042,G75565);
  nand GNAME77128(G77128,G77127,G77126);
  or GNAME77129(G77129,G80991,G75557);
  or GNAME77130(G77130,G81043,G75564);
  nand GNAME77131(G77131,G77130,G77129);
  or GNAME77132(G77132,G81079,G75539);
  or GNAME77133(G77133,G81061,G75573);
  nand GNAME77134(G77134,G77133,G77132);
  or GNAME77135(G77135,G80986,G75538);
  or GNAME77136(G77136,G81044,G75572);
  nand GNAME77137(G77137,G77136,G77135);
  or GNAME77138(G77138,G80992,G75537);
  or GNAME77139(G77139,G81046,G75571);
  nand GNAME77140(G77140,G77139,G77138);
  or GNAME77141(G77141,G81080,G75546);
  or GNAME77142(G77142,G81062,G75580);
  nand GNAME77143(G77143,G77142,G77141);
  or GNAME77144(G77144,G80987,G75545);
  or GNAME77145(G77145,G81045,G75579);
  nand GNAME77146(G77146,G77145,G77144);
  or GNAME77147(G77147,G80993,G75544);
  or GNAME77148(G77148,G81047,G75578);
  nand GNAME77149(G77149,G77148,G77147);
  or GNAME77150(G77150,G81079,G75573);
  or GNAME77151(G77151,G81061,G75587);
  nand GNAME77152(G77152,G77151,G77150);
  or GNAME77153(G77153,G80986,G75572);
  or GNAME77154(G77154,G81044,G75586);
  nand GNAME77155(G77155,G77154,G77153);
  or GNAME77156(G77156,G80992,G75571);
  or GNAME77157(G77157,G81046,G75585);
  nand GNAME77158(G77158,G77157,G77156);
  or GNAME77159(G77159,G81080,G75580);
  or GNAME77160(G77160,G81062,G75594);
  nand GNAME77161(G77161,G77160,G77159);
  or GNAME77162(G77162,G80987,G75579);
  or GNAME77163(G77163,G81045,G75593);
  nand GNAME77164(G77164,G77163,G77162);
  or GNAME77165(G77165,G80993,G75578);
  or GNAME77166(G77166,G81047,G75592);
  nand GNAME77167(G77167,G77166,G77165);
  or GNAME77168(G77168,G81066,G75563);
  or GNAME77169(G77169,G81075,G75607);
  nand GNAME77170(G77170,G77169,G77168);
  or GNAME77171(G77171,G81000,G75562);
  or GNAME77172(G77172,G81051,G75606);
  nand GNAME77173(G77173,G77172,G77171);
  or GNAME77174(G77174,G81063,G75561);
  or GNAME77175(G77175,G81069,G75605);
  nand GNAME77176(G77176,G77175,G77174);
  or GNAME77177(G77177,G81066,G75607);
  or GNAME77178(G77178,G81075,G75614);
  nand GNAME77179(G77179,G77178,G77177);
  or GNAME77180(G77180,G81000,G75606);
  or GNAME77181(G77181,G81051,G75613);
  nand GNAME77182(G77182,G77181,G77180);
  or GNAME77183(G77183,G81063,G75605);
  or GNAME77184(G77184,G81069,G75612);
  nand GNAME77185(G77185,G77184,G77183);
  or GNAME77186(G77186,G81067,G75584);
  or GNAME77187(G77187,G81076,G75619);
  nand GNAME77188(G77188,G77187,G77186);
  or GNAME77189(G77189,G81001,G75583);
  or GNAME77190(G77190,G81052,G75618);
  nand GNAME77191(G77191,G77190,G77189);
  or GNAME77192(G77192,G81064,G75582);
  or GNAME77193(G77193,G81070,G75617);
  nand GNAME77194(G77194,G77193,G77192);
  or GNAME77195(G77195,G81068,G75591);
  or GNAME77196(G77196,G81077,G75626);
  nand GNAME77197(G77197,G77196,G77195);
  or GNAME77198(G77198,G81002,G75590);
  or GNAME77199(G77199,G81053,G75625);
  nand GNAME77200(G77200,G77199,G77198);
  or GNAME77201(G77201,G81065,G75589);
  or GNAME77202(G77202,G81071,G75624);
  nand GNAME77203(G77203,G77202,G77201);
  or GNAME77204(G77204,G81067,G75619);
  or GNAME77205(G77205,G81076,G75633);
  nand GNAME77206(G77206,G77205,G77204);
  or GNAME77207(G77207,G81001,G75618);
  or GNAME77208(G77208,G81052,G75632);
  nand GNAME77209(G77209,G77208,G77207);
  or GNAME77210(G77210,G81064,G75617);
  or GNAME77211(G77211,G81070,G75631);
  nand GNAME77212(G77212,G77211,G77210);
  or GNAME77213(G77213,G81068,G75626);
  or GNAME77214(G77214,G81077,G75638);
  nand GNAME77215(G77215,G77214,G77213);
  or GNAME77216(G77216,G81002,G75625);
  or GNAME77217(G77217,G81053,G75637);
  nand GNAME77218(G77218,G77217,G77216);
  or GNAME77219(G77219,G81065,G75624);
  or GNAME77220(G77220,G81071,G75636);
  nand GNAME77221(G77221,G77220,G77219);
  or GNAME77222(G77222,G81033,G75567);
  or GNAME77223(G77223,G81015,G75611);
  nand GNAME77224(G77224,G77223,G77222);
  or GNAME77225(G77225,G75597,G81018);
  or GNAME77226(G77226,G81012,G75641);
  nand GNAME77227(G77227,G77226,G77225);
  or GNAME77228(G77228,G81034,G75588);
  or GNAME77229(G77229,G81016,G75623);
  nand GNAME77230(G77230,G77229,G77228);
  or GNAME77231(G77231,G75600,G81019);
  or GNAME77232(G77232,G81013,G75642);
  nand GNAME77233(G77233,G77232,G77231);
  or GNAME77234(G77234,G81035,G75595);
  or GNAME77235(G77235,G81017,G75630);
  nand GNAME77236(G77236,G77235,G77234);
  or GNAME77237(G77237,G75601,G81020);
  or GNAME77238(G77238,G81014,G75643);
  nand GNAME77239(G77239,G77238,G77237);
  or GNAME77240(G77240,G81078,G75566);
  or GNAME77241(G77241,G81072,G75610);
  nand GNAME77242(G77242,G77241,G77240);
  or GNAME77243(G77243,G80985,G75565);
  or GNAME77244(G77244,G81042,G75609);
  nand GNAME77245(G77245,G77244,G77243);
  or GNAME77246(G77246,G80991,G75564);
  or GNAME77247(G77247,G81043,G75608);
  nand GNAME77248(G77248,G77247,G77246);
  or GNAME77249(G77249,G81027,G75610);
  or GNAME77250(G77250,G81072,G75602);
  nand GNAME77251(G77251,G77250,G77249);
  or GNAME77252(G77252,G80985,G75609);
  or GNAME77253(G77253,G81042,G75653);
  nand GNAME77254(G77254,G77253,G77252);
  or GNAME77255(G77255,G80991,G75608);
  or GNAME77256(G77256,G81043,G75615);
  nand GNAME77257(G77257,G77256,G77255);
  or GNAME77258(G77258,G81079,G75587);
  or GNAME77259(G77259,G81073,G75622);
  nand GNAME77260(G77260,G77259,G77258);
  or GNAME77261(G77261,G80986,G75586);
  or GNAME77262(G77262,G81044,G75621);
  nand GNAME77263(G77263,G77262,G77261);
  or GNAME77264(G77264,G80992,G75585);
  or GNAME77265(G77265,G81046,G75620);
  nand GNAME77266(G77266,G77265,G77264);
  or GNAME77267(G77267,G81080,G75594);
  or GNAME77268(G77268,G81074,G75629);
  nand GNAME77269(G77269,G77268,G77267);
  or GNAME77270(G77270,G80987,G75593);
  or GNAME77271(G77271,G81045,G75628);
  nand GNAME77272(G77272,G77271,G77270);
  or GNAME77273(G77273,G80993,G75592);
  or GNAME77274(G77274,G81047,G75627);
  nand GNAME77275(G77275,G77274,G77273);
  or GNAME77276(G77276,G81029,G75622);
  or GNAME77277(G77277,G81073,G75603);
  nand GNAME77278(G77278,G77277,G77276);
  or GNAME77279(G77279,G80986,G75621);
  or GNAME77280(G77280,G81044,G75666);
  nand GNAME77281(G77281,G77280,G77279);
  or GNAME77282(G77282,G80992,G75620);
  or GNAME77283(G77283,G81046,G75634);
  nand GNAME77284(G77284,G77283,G77282);
  or GNAME77285(G77285,G81031,G75629);
  or GNAME77286(G77286,G81074,G75604);
  nand GNAME77287(G77287,G77286,G77285);
  or GNAME77288(G77288,G80987,G75628);
  or GNAME77289(G77289,G81045,G75672);
  nand GNAME77290(G77290,G77289,G77288);
  or GNAME77291(G77291,G80993,G75627);
  or GNAME77292(G77292,G81047,G75639);
  nand GNAME77293(G77293,G77292,G77291);
  or GNAME77294(G77294,G81000,G75613);
  or GNAME77295(G77295,G81051,G75656);
  nand GNAME77296(G77296,G77295,G77294);
  or GNAME77297(G77297,G81033,G75616);
  or GNAME77298(G77298,G81024,G75655);
  nand GNAME77299(G77299,G77298,G77297);
  or GNAME77300(G77300,G81066,G75614);
  or GNAME77301(G77301,G81075,G75654);
  nand GNAME77302(G77302,G77301,G77300);
  or GNAME77303(G77303,G81001,G75632);
  or GNAME77304(G77304,G81052,G75669);
  nand GNAME77305(G77305,G77304,G77303);
  or GNAME77306(G77306,G81034,G75635);
  or GNAME77307(G77307,G81025,G75668);
  nand GNAME77308(G77308,G77307,G77306);
  or GNAME77309(G77309,G81067,G75633);
  or GNAME77310(G77310,G81076,G75667);
  nand GNAME77311(G77311,G77310,G77309);
  or GNAME77312(G77312,G81002,G75637);
  or GNAME77313(G77313,G81053,G75675);
  nand GNAME77314(G77314,G77313,G77312);
  or GNAME77315(G77315,G81035,G75640);
  or GNAME77316(G77316,G81026,G75674);
  nand GNAME77317(G77317,G77316,G77315);
  or GNAME77318(G77318,G81068,G75638);
  or GNAME77319(G77319,G81077,G75673);
  nand GNAME77320(G77320,G77319,G77318);
  or GNAME77321(G77321,G81066,G75654);
  or GNAME77322(G77322,G81075,G75665);
  nand GNAME77323(G77323,G77322,G77321);
  or GNAME77324(G77324,G81063,G75658);
  or GNAME77325(G77325,G81069,G75664);
  nand GNAME77326(G77326,G77325,G77324);
  or GNAME77327(G77327,G81067,G75667);
  or GNAME77328(G77328,G81076,G75684);
  nand GNAME77329(G77329,G77328,G77327);
  or GNAME77330(G77330,G81064,G75671);
  or GNAME77331(G77331,G81070,G75683);
  nand GNAME77332(G77332,G77331,G77330);
  or GNAME77333(G77333,G81068,G75673);
  or GNAME77334(G77334,G81077,G75691);
  nand GNAME77335(G77335,G77334,G77333);
  or GNAME77336(G77336,G81065,G75677);
  or GNAME77337(G77337,G81071,G75690);
  nand GNAME77338(G77338,G77337,G77336);
  or GNAME77339(G77339,G81027,G75602);
  or GNAME77340(G77340,G81072,G75662);
  nand GNAME77341(G77341,G77340,G77339);
  or GNAME77342(G77342,G81029,G75603);
  or GNAME77343(G77343,G81073,G75681);
  nand GNAME77344(G77344,G77343,G77342);
  or GNAME77345(G77345,G81031,G75604);
  or GNAME77346(G77346,G81074,G75688);
  nand GNAME77347(G77347,G77346,G77345);
  or GNAME77348(G77348,G81063,G75612);
  or GNAME77349(G77349,G81069,G75658);
  nand GNAME77350(G77350,G77349,G77348);
  or GNAME77351(G77351,G80991,G75615);
  or GNAME77352(G77352,G81043,G75657);
  nand GNAME77353(G77353,G77352,G77351);
  or GNAME77354(G77354,G81048,G74115);
  or GNAME77355(G77355,G80980,G77767);
  nand GNAME77356(G77356,G77355,G77354);
  or GNAME77357(G77357,G81027,G75662);
  or GNAME77358(G77358,G81072,G75663);
  nand GNAME77359(G77359,G77358,G77357);
  or GNAME77360(G77360,G80991,G75657);
  or GNAME77361(G77361,G81043,G75661);
  nand GNAME77362(G77362,G77361,G77360);
  or GNAME77363(G77363,G81000,G75656);
  or GNAME77364(G77364,G81051,G75660);
  nand GNAME77365(G77365,G77364,G77363);
  or GNAME77366(G77366,G81064,G75631);
  or GNAME77367(G77367,G81070,G75671);
  nand GNAME77368(G77368,G77367,G77366);
  or GNAME77369(G77369,G80992,G75634);
  or GNAME77370(G77370,G81046,G75670);
  nand GNAME77371(G77371,G77370,G77369);
  or GNAME77372(G77372,G81049,G74118);
  or GNAME77373(G77373,G80981,G77766);
  nand GNAME77374(G77374,G77373,G77372);
  or GNAME77375(G77375,G81065,G75636);
  or GNAME77376(G77376,G81071,G75677);
  nand GNAME77377(G77377,G77376,G77375);
  or GNAME77378(G77378,G80993,G75639);
  or GNAME77379(G77379,G81047,G75676);
  nand GNAME77380(G77380,G77379,G77378);
  or GNAME77381(G77381,G81050,G74121);
  or GNAME77382(G77382,G80982,G77768);
  nand GNAME77383(G77383,G77382,G77381);
  or GNAME77384(G77384,G81029,G75681);
  or GNAME77385(G77385,G81073,G75682);
  nand GNAME77386(G77386,G77385,G77384);
  or GNAME77387(G77387,G80992,G75670);
  or GNAME77388(G77388,G81046,G75680);
  nand GNAME77389(G77389,G77388,G77387);
  or GNAME77390(G77390,G81001,G75669);
  or GNAME77391(G77391,G81052,G75679);
  nand GNAME77392(G77392,G77391,G77390);
  or GNAME77393(G77393,G81031,G75688);
  or GNAME77394(G77394,G81074,G75689);
  nand GNAME77395(G77395,G77394,G77393);
  or GNAME77396(G77396,G80993,G75676);
  or GNAME77397(G77397,G81047,G75687);
  nand GNAME77398(G77398,G77397,G77396);
  or GNAME77399(G77399,G81002,G75675);
  or GNAME77400(G77400,G81053,G75686);
  nand GNAME77401(G77401,G77400,G77399);
  or GNAME77402(G77402,G81063,G75664);
  or GNAME77403(G77403,G81069,G75719);
  nand GNAME77404(G77404,G77403,G77402);
  or GNAME77405(G77405,G81028,G75659);
  or GNAME77406(G77406,G81024,G75718);
  nand GNAME77407(G77407,G77406,G77405);
  or GNAME77408(G77408,G81027,G75663);
  or GNAME77409(G77409,G81072,G75717);
  nand GNAME77410(G77410,G77409,G77408);
  or GNAME77411(G77411,G81027,G75717);
  or GNAME77412(G77412,G81072,G75703);
  nand GNAME77413(G77413,G77412,G77411);
  or GNAME77414(G77414,G81000,G75716);
  or GNAME77415(G77415,G81051,G75720);
  nand GNAME77416(G77416,G77415,G77414);
  or GNAME77417(G77417,G81063,G75719);
  or GNAME77418(G77418,G81069,G75701);
  nand GNAME77419(G77419,G77418,G77417);
  or GNAME77420(G77420,G81064,G75683);
  or GNAME77421(G77421,G81070,G75726);
  nand GNAME77422(G77422,G77421,G77420);
  or GNAME77423(G77423,G81030,G75678);
  or GNAME77424(G77424,G81025,G75725);
  nand GNAME77425(G77425,G77424,G77423);
  or GNAME77426(G77426,G81029,G75682);
  or GNAME77427(G77427,G81073,G75724);
  nand GNAME77428(G77428,G77427,G77426);
  or GNAME77429(G77429,G81065,G75690);
  or GNAME77430(G77430,G81071,G75730);
  nand GNAME77431(G77431,G77430,G77429);
  or GNAME77432(G77432,G81032,G75685);
  or GNAME77433(G77433,G81026,G75729);
  nand GNAME77434(G77434,G77433,G77432);
  or GNAME77435(G77435,G81031,G75689);
  or GNAME77436(G77436,G81074,G75728);
  nand GNAME77437(G77437,G77436,G77435);
  or GNAME77438(G77438,G81029,G75724);
  or GNAME77439(G77439,G81073,G75708);
  nand GNAME77440(G77440,G77439,G77438);
  or GNAME77441(G77441,G81001,G75723);
  or GNAME77442(G77442,G81052,G75731);
  nand GNAME77443(G77443,G77442,G77441);
  or GNAME77444(G77444,G81064,G75726);
  or GNAME77445(G77445,G81070,G75706);
  nand GNAME77446(G77446,G77445,G77444);
  or GNAME77447(G77447,G81031,G75728);
  or GNAME77448(G77448,G81074,G75713);
  nand GNAME77449(G77449,G77448,G77447);
  or GNAME77450(G77450,G81002,G75727);
  or GNAME77451(G77451,G81053,G75734);
  nand GNAME77452(G77452,G77451,G77450);
  or GNAME77453(G77453,G81065,G75730);
  or GNAME77454(G77454,G81071,G75711);
  nand GNAME77455(G77455,G77454,G77453);
  or GNAME77456(G77456,G81066,G75650);
  or GNAME77457(G77457,G81075,G75722);
  nand GNAME77458(G77458,G77457,G77456);
  or GNAME77459(G77459,G81027,G75703);
  or GNAME77460(G77460,G81072,G75704);
  nand GNAME77461(G77461,G77460,G77459);
  or GNAME77462(G77462,G81063,G75701);
  or GNAME77463(G77463,G81069,G75702);
  nand GNAME77464(G77464,G77463,G77462);
  or GNAME77465(G77465,G81067,G75651);
  or GNAME77466(G77466,G81076,G75733);
  nand GNAME77467(G77467,G77466,G77465);
  or GNAME77468(G77468,G81068,G75652);
  or GNAME77469(G77469,G81077,G75736);
  nand GNAME77470(G77470,G77469,G77468);
  or GNAME77471(G77471,G81029,G75708);
  or GNAME77472(G77472,G81073,G75709);
  nand GNAME77473(G77473,G77472,G77471);
  or GNAME77474(G77474,G81064,G75706);
  or GNAME77475(G77475,G81070,G75707);
  nand GNAME77476(G77476,G77475,G77474);
  or GNAME77477(G77477,G81031,G75713);
  or GNAME77478(G77478,G81074,G75714);
  nand GNAME77479(G77479,G77478,G77477);
  or GNAME77480(G77480,G81065,G75711);
  or GNAME77481(G77481,G81071,G75712);
  nand GNAME77482(G77482,G77481,G77480);
  or GNAME77483(G77483,G81066,G75665);
  or GNAME77484(G77484,G81075,G75650);
  nand GNAME77485(G77485,G77484,G77483);
  or GNAME77486(G77486,G81000,G75660);
  or GNAME77487(G77487,G81051,G75716);
  nand GNAME77488(G77488,G77487,G77486);
  or GNAME77489(G77489,G81054,G74124);
  or GNAME77490(G77490,G80988,G77769);
  nand GNAME77491(G77491,G77490,G77489);
  or GNAME77492(G77492,G81067,G75684);
  or GNAME77493(G77493,G81076,G75651);
  nand GNAME77494(G77494,G77493,G77492);
  or GNAME77495(G77495,G81001,G75679);
  or GNAME77496(G77496,G81052,G75723);
  nand GNAME77497(G77497,G77496,G77495);
  or GNAME77498(G77498,G81055,G74127);
  or GNAME77499(G77499,G80989,G77770);
  nand GNAME77500(G77500,G77499,G77498);
  or GNAME77501(G77501,G81068,G75691);
  or GNAME77502(G77502,G81077,G75652);
  nand GNAME77503(G77503,G77502,G77501);
  or GNAME77504(G77504,G81002,G75686);
  or GNAME77505(G77505,G81053,G75727);
  nand GNAME77506(G77506,G77505,G77504);
  or GNAME77507(G77507,G81056,G74130);
  or GNAME77508(G77508,G80990,G77771);
  nand GNAME77509(G77509,G77508,G77507);
  or GNAME77510(G77510,G81066,G75722);
  or GNAME77511(G77511,G81075,G75705);
  nand GNAME77512(G77512,G77511,G77510);
  or GNAME77513(G77513,G81028,G75721);
  or GNAME77514(G77514,G81024,G75761);
  nand GNAME77515(G77515,G77514,G77513);
  or GNAME77516(G77516,G81003,G74133);
  or GNAME77517(G77517,G80994,G77774);
  nand GNAME77518(G77518,G77517,G77516);
  or GNAME77519(G77519,G81067,G75733);
  or GNAME77520(G77520,G81076,G75710);
  nand GNAME77521(G77521,G77520,G77519);
  or GNAME77522(G77522,G81030,G75732);
  or GNAME77523(G77523,G81025,G75767);
  nand GNAME77524(G77524,G77523,G77522);
  or GNAME77525(G77525,G81005,G74136);
  or GNAME77526(G77526,G80996,G77776);
  nand GNAME77527(G77527,G77526,G77525);
  or GNAME77528(G77528,G81068,G75736);
  or GNAME77529(G77529,G81077,G75715);
  nand GNAME77530(G77530,G77529,G77528);
  or GNAME77531(G77531,G81032,G75735);
  or GNAME77532(G77532,G81026,G75771);
  nand GNAME77533(G77533,G77532,G77531);
  or GNAME77534(G77534,G81006,G74139);
  or GNAME77535(G77535,G80997,G77777);
  nand GNAME77536(G77536,G77535,G77534);
  or GNAME77537(G77537,G81066,G75758);
  or GNAME77538(G77538,G81075,G75750);
  nand GNAME77539(G77539,G77538,G77537);
  or GNAME77540(G77540,G81027,G75760);
  or GNAME77541(G77541,G81072,G75751);
  nand GNAME77542(G77542,G77541,G77540);
  or GNAME77543(G77543,G81004,G74142);
  or GNAME77544(G77544,G80995,G77775);
  nand GNAME77545(G77545,G77544,G77543);
  or GNAME77546(G77546,G81067,G75764);
  or GNAME77547(G77547,G81076,G75754);
  nand GNAME77548(G77548,G77547,G77546);
  or GNAME77549(G77549,G81029,G75766);
  or GNAME77550(G77550,G81073,G75755);
  nand GNAME77551(G77551,G77550,G77549);
  or GNAME77552(G77552,G81007,G74145);
  or GNAME77553(G77553,G80998,G77778);
  nand GNAME77554(G77554,G77553,G77552);
  or GNAME77555(G77555,G81068,G75768);
  or GNAME77556(G77556,G81077,G75756);
  nand GNAME77557(G77557,G77556,G77555);
  or GNAME77558(G77558,G81031,G75770);
  or GNAME77559(G77559,G81074,G75757);
  nand GNAME77560(G77560,G77559,G77558);
  or GNAME77561(G77561,G81008,G74148);
  or GNAME77562(G77562,G80999,G77779);
  nand GNAME77563(G77563,G77562,G77561);
  or GNAME77564(G77564,G81027,G75704);
  or GNAME77565(G77565,G81072,G75760);
  nand GNAME77566(G77566,G77565,G77564);
  or GNAME77567(G77567,G81063,G75702);
  or GNAME77568(G77568,G81069,G75759);
  nand GNAME77569(G77569,G77568,G77567);
  or GNAME77570(G77570,G81066,G75705);
  or GNAME77571(G77571,G81075,G75758);
  nand GNAME77572(G77572,G77571,G77570);
  or GNAME77573(G77573,G81029,G75709);
  or GNAME77574(G77574,G81073,G75766);
  nand GNAME77575(G77575,G77574,G77573);
  or GNAME77576(G77576,G81064,G75707);
  or GNAME77577(G77577,G81070,G75765);
  nand GNAME77578(G77578,G77577,G77576);
  or GNAME77579(G77579,G81067,G75710);
  or GNAME77580(G77580,G81076,G75764);
  nand GNAME77581(G77581,G77580,G77579);
  or GNAME77582(G77582,G81031,G75714);
  or GNAME77583(G77583,G81074,G75770);
  nand GNAME77584(G77584,G77583,G77582);
  or GNAME77585(G77585,G81065,G75712);
  or GNAME77586(G77586,G81071,G75769);
  nand GNAME77587(G77587,G77586,G77585);
  or GNAME77588(G77588,G81068,G75715);
  or GNAME77589(G77589,G81077,G75768);
  nand GNAME77590(G77590,G77589,G77588);
  or GNAME77591(G77591,G81028,G75796);
  or GNAME77592(G77592,G81024,G75797);
  nand GNAME77593(G77593,G77592,G77591);
  or GNAME77594(G77594,G81027,G75795);
  or GNAME77595(G77595,G81072,G75794);
  nand GNAME77596(G77596,G77595,G77594);
  or GNAME77597(G77597,G81081,G74151);
  or GNAME77598(G77598,G81057,G77780);
  nand GNAME77599(G77599,G77598,G77597);
  or GNAME77600(G77600,G81030,G75800);
  or GNAME77601(G77601,G81025,G75801);
  nand GNAME77602(G77602,G77601,G77600);
  or GNAME77603(G77603,G81029,G75798);
  or GNAME77604(G77604,G81073,G75799);
  nand GNAME77605(G77605,G77604,G77603);
  or GNAME77606(G77606,G81082,G74154);
  or GNAME77607(G77607,G81058,G77781);
  nand GNAME77608(G77608,G77607,G77606);
  or GNAME77609(G77609,G81032,G75804);
  or GNAME77610(G77610,G81026,G75805);
  nand GNAME77611(G77611,G77610,G77609);
  or GNAME77612(G77612,G81031,G75802);
  or GNAME77613(G77613,G81074,G75803);
  nand GNAME77614(G77614,G77613,G77612);
  or GNAME77615(G77615,G81083,G74157);
  or GNAME77616(G77616,G81059,G77782);
  nand GNAME77617(G77617,G77616,G77615);
  or GNAME77618(G77618,G81027,G75751);
  or GNAME77619(G77619,G81072,G75795);
  nand GNAME77620(G77620,G77619,G77618);
  or GNAME77621(G77621,G81066,G75750);
  or GNAME77622(G77622,G81075,G75763);
  nand GNAME77623(G77623,G77622,G77621);
  or GNAME77624(G77624,G81029,G75755);
  or GNAME77625(G77625,G81073,G75798);
  nand GNAME77626(G77626,G77625,G77624);
  or GNAME77627(G77627,G81067,G75754);
  or GNAME77628(G77628,G81076,G75774);
  nand GNAME77629(G77629,G77628,G77627);
  or GNAME77630(G77630,G81031,G75757);
  or GNAME77631(G77631,G81074,G75802);
  nand GNAME77632(G77632,G77631,G77630);
  or GNAME77633(G77633,G81068,G75756);
  or GNAME77634(G77634,G81077,G75775);
  nand GNAME77635(G77635,G77634,G77633);
  or GNAME77636(G77636,G81028,G75749);
  or GNAME77637(G77637,G81024,G75762);
  nand GNAME77638(G77638,G77637,G77636);
  or GNAME77639(G77639,G81030,G75752);
  or GNAME77640(G77640,G81025,G75772);
  nand GNAME77641(G77641,G77640,G77639);
  or GNAME77642(G77642,G81032,G75753);
  or GNAME77643(G77643,G81026,G75773);
  nand GNAME77644(G77644,G77643,G77642);
  or GNAME77645(G77645,G81027,G75794);
  or GNAME77646(G77646,G81072,G75807);
  nand GNAME77647(G77647,G77646,G77645);
  or GNAME77648(G77648,G81029,G75799);
  or GNAME77649(G77649,G81073,G75809);
  nand GNAME77650(G77650,G77649,G77648);
  or GNAME77651(G77651,G81031,G75803);
  or GNAME77652(G77652,G81074,G75811);
  nand GNAME77653(G77653,G77652,G77651);
  or GNAME77654(G77654,G81033,G74160);
  or GNAME77655(G77655,G81015,G77785);
  nand GNAME77656(G77656,G77655,G77654);
  or GNAME77657(G77657,G81034,G74163);
  or GNAME77658(G77658,G81016,G77787);
  nand GNAME77659(G77659,G77658,G77657);
  or GNAME77660(G77660,G81035,G74166);
  or GNAME77661(G77661,G81017,G77788);
  nand GNAME77662(G77662,G77661,G77660);
  or GNAME77663(G77663,G81028,G75806);
  or GNAME77664(G77664,G81024,G75818);
  nand GNAME77665(G77665,G77664,G77663);
  or GNAME77666(G77666,G75812,G81009);
  or GNAME77667(G77667,G81021,G75824);
  nand GNAME77668(G77668,G77667,G77666);
  or GNAME77669(G77669,G81030,G75808);
  or GNAME77670(G77670,G81025,G75820);
  nand GNAME77671(G77671,G77670,G77669);
  or GNAME77672(G77672,G75816,G81010);
  or GNAME77673(G77673,G81022,G75826);
  nand GNAME77674(G77674,G77673,G77672);
  or GNAME77675(G77675,G81032,G75810);
  or GNAME77676(G77676,G81026,G75822);
  nand GNAME77677(G77677,G77676,G77675);
  or GNAME77678(G77678,G75817,G81011);
  or GNAME77679(G77679,G81023,G75828);
  nand GNAME77680(G77680,G77679,G77678);
  or GNAME77681(G77681,G75825,G81009);
  or GNAME77682(G77682,G81021,G75830);
  nand GNAME77683(G77683,G77682,G77681);
  or GNAME77684(G77684,G75827,G81010);
  or GNAME77685(G77685,G81022,G75832);
  nand GNAME77686(G77686,G77685,G77684);
  or GNAME77687(G77687,G75829,G81011);
  or GNAME77688(G77688,G81023,G75834);
  nand GNAME77689(G77689,G77688,G77687);
  not GNAME77690(G77690,G79117);
  not GNAME77691(G77691,G77882);
  not GNAME77692(G77692,G77895);
  not GNAME77693(G77693,G2344);
  not GNAME77694(G77694,G1928);
  not GNAME77695(G77695,G1512);
  not GNAME77696(G77696,G80851);
  not GNAME77697(G77697,G80856);
  not GNAME77698(G77698,G80855);
  not GNAME77699(G77699,G80857);
  not GNAME77700(G77700,G80865);
  not GNAME77701(G77701,G80864);
  not GNAME77702(G77702,G80866);
  not GNAME77703(G77703,G80861);
  not GNAME77704(G77704,G80862);
  not GNAME77705(G77705,G80863);
  not GNAME77706(G77706,G80873);
  not GNAME77707(G77707,G80874);
  not GNAME77708(G77708,G80875);
  not GNAME77709(G77709,G80870);
  not GNAME77710(G77710,G80871);
  not GNAME77711(G77711,G80872);
  not GNAME77712(G77712,G80882);
  not GNAME77713(G77713,G80883);
  not GNAME77714(G77714,G80884);
  not GNAME77715(G77715,G80879);
  not GNAME77716(G77716,G80880);
  not GNAME77717(G77717,G80881);
  not GNAME77718(G77718,G80891);
  not GNAME77719(G77719,G80892);
  not GNAME77720(G77720,G80893);
  not GNAME77721(G77721,G80888);
  not GNAME77722(G77722,G80889);
  not GNAME77723(G77723,G80890);
  not GNAME77724(G77724,G80898);
  not GNAME77725(G77725,G80900);
  not GNAME77726(G77726,G80902);
  not GNAME77727(G77727,G80897);
  not GNAME77728(G77728,G80899);
  not GNAME77729(G77729,G80901);
  not GNAME77730(G77730,G80916);
  not GNAME77731(G77731,G80919);
  not GNAME77732(G77732,G80921);
  not GNAME77733(G77733,G80935);
  not GNAME77734(G77734,G80937);
  not GNAME77735(G77735,G80939);
  not GNAME77736(G77736,G80917);
  not GNAME77737(G77737,G80920);
  not GNAME77738(G77738,G80922);
  not GNAME77739(G77739,G80918);
  not GNAME77740(G77740,G80923);
  not GNAME77741(G77741,G80924);
  not GNAME77742(G77742,G80940);
  not GNAME77743(G77743,G80941);
  not GNAME77744(G77744,G80942);
  not GNAME77745(G77745,G80934);
  not GNAME77746(G77746,G80949);
  not GNAME77747(G77747,G80936);
  not GNAME77748(G77748,G80938);
  not GNAME77749(G77749,G80950);
  not GNAME77750(G77750,G80951);
  not GNAME77751(G77751,G80946);
  not GNAME77752(G77752,G80947);
  not GNAME77753(G77753,G80954);
  not GNAME77754(G77754,G80957);
  not GNAME77755(G77755,G80953);
  not GNAME77756(G77756,G80956);
  not GNAME77757(G77757,G80948);
  not GNAME77758(G77758,G80967);
  not GNAME77759(G77759,G80952);
  not GNAME77760(G77760,G80955);
  not GNAME77761(G77761,G80969);
  not GNAME77762(G77762,G80971);
  not GNAME77763(G77763,G80968);
  not GNAME77764(G77764,G80970);
  not GNAME77765(G77765,G80972);
  not GNAME77766(G77766,G80909);
  not GNAME77767(G77767,G80908);
  not GNAME77768(G77768,G80910);
  not GNAME77769(G77769,G80911);
  not GNAME77770(G77770,G80912);
  not GNAME77771(G77771,G80913);
  not GNAME77772(G77772,G80914);
  not GNAME77773(G77773,G80915);
  not GNAME77774(G77774,G80928);
  not GNAME77775(G77775,G80943);
  not GNAME77776(G77776,G80929);
  not GNAME77777(G77777,G80930);
  not GNAME77778(G77778,G80944);
  not GNAME77779(G77779,G80945);
  not GNAME77780(G77780,G80958);
  not GNAME77781(G77781,G80959);
  not GNAME77782(G77782,G80960);
  not GNAME77783(G77783,G80962);
  not GNAME77784(G77784,G80963);
  not GNAME77785(G77785,G80973);
  not GNAME77786(G77786,G80961);
  not GNAME77787(G77787,G80974);
  not GNAME77788(G77788,G80975);
  not GNAME77789(G77789,G80976);
  not GNAME77790(G77790,G80977);
  not GNAME77791(G77791,G80978);
  not GNAME77792(G77792,G75176);
  not GNAME77793(G77793,G75175);
  not GNAME77794(G77794,G75177);
  not GNAME77795(G77795,G75181);
  not GNAME77796(G77796,G75182);
  not GNAME77797(G77797,G75183);
  not GNAME77798(G77798,G75187);
  not GNAME77799(G77799,G75188);
  not GNAME77800(G77800,G75189);
  not GNAME77801(G77801,G75193);
  not GNAME77802(G77802,G75194);
  not GNAME77803(G77803,G75195);
  not GNAME77804(G77804,G75199);
  not GNAME77805(G77805,G75200);
  not GNAME77806(G77806,G75201);
  not GNAME77807(G77807,G75205);
  not GNAME77808(G77808,G75206);
  not GNAME77809(G77809,G75207);
  not GNAME77810(G77810,G75214);
  not GNAME77811(G77811,G75215);
  not GNAME77812(G77812,G75216);
  nand GNAME77813(G77813,G75245,G77842);
  nand GNAME77814(G77814,G75246,G77843);
  nand GNAME77815(G77815,G75247,G77844);
  nand GNAME77816(G77816,G75248,G77845);
  nand GNAME77817(G77817,G75249,G77846);
  nand GNAME77818(G77818,G75250,G77847);
  nand GNAME77819(G77819,G75251,G77848);
  nand GNAME77820(G77820,G75252,G77849);
  nand GNAME77821(G77821,G75253,G77850);
  nand GNAME77822(G77822,G75254,G77851);
  nand GNAME77823(G77823,G75255,G77852);
  nand GNAME77824(G77824,G75256,G77853);
  nand GNAME77825(G77825,G75260,G77854);
  nand GNAME77826(G77826,G75257,G77855);
  nand GNAME77827(G77827,G75258,G77856);
  nand GNAME77828(G77828,G75259,G77857);
  nand GNAME77829(G77829,G75261,G77858);
  nand GNAME77830(G77830,G75262,G77859);
  nand GNAME77831(G77831,G77860,G77693);
  nand GNAME77832(G77832,G77861,G77694);
  nand GNAME77833(G77833,G77862,G77695);
  nand GNAME77834(G77834,G75263,G77863);
  nand GNAME77835(G77835,G75264,G77864);
  nand GNAME77836(G77836,G75265,G77865);
  xor GNAME77837(G77837,G77960,G77934);
  xor GNAME77838(G77838,G74855,G80599);
  xor GNAME77839(G77839,G74837,G80586);
  xor GNAME77840(G77840,G74843,G80612);
  xor GNAME77841(G77841,G80846,G72455);
  xor GNAME77842(G77842,G2678,G2699);
  xor GNAME77843(G77843,G2262,G2283);
  xor GNAME77844(G77844,G1846,G1867);
  xor GNAME77845(G77845,G2636,G2657);
  xor GNAME77846(G77846,G2220,G2241);
  xor GNAME77847(G77847,G1804,G1825);
  xor GNAME77848(G77848,G2552,G2573);
  xor GNAME77849(G77849,G2136,G2157);
  xor GNAME77850(G77850,G1720,G1741);
  xor GNAME77851(G77851,G2594,G2615);
  xor GNAME77852(G77852,G2178,G2199);
  xor GNAME77853(G77853,G1762,G1783);
  xor GNAME77854(G77854,G2428,G2449);
  xor GNAME77855(G77855,G2470,G2491);
  xor GNAME77856(G77856,G2054,G2075);
  xor GNAME77857(G77857,G1638,G1659);
  xor GNAME77858(G77858,G2012,G2033);
  xor GNAME77859(G77859,G1596,G1617);
  xor GNAME77860(G77860,G2344,G2365);
  xor GNAME77861(G77861,G1928,G1949);
  xor GNAME77862(G77862,G1512,G1533);
  xor GNAME77863(G77863,G2386,G2407);
  xor GNAME77864(G77864,G1970,G1991);
  xor GNAME77865(G77865,G1554,G1575);
  xor GNAME77866(G77866,G74111,G74114);
  xor GNAME77867(G77867,G64175,G74187);
  xor GNAME77868(G77868,G70430,G77867);
  xor GNAME77869(G77869,G64160,G74189);
  xor GNAME77870(G77870,G70415,G77869);
  xor GNAME77871(G77871,G64190,G74191);
  xor GNAME77872(G77872,G70445,G77871);
  dff DFF_77881(CK,G77880,G70395);
  and GNAME77882(G77882,G77880,G77883);
  nand GNAME77883(G77883,G80,G77885);
  buf GNAME77884(G77884,G77880);
  buf GNAME77885(G77885,G77875);
  dff DFF_77894(CK,G77893,G70380);
  and GNAME77895(G77895,G77893,G77896);
  nand GNAME77896(G77896,G80,G77898);
  buf GNAME77897(G77897,G77893);
  buf GNAME77898(G77898,G77888);
  dff DFF_77907(CK,G77906,G68100);
  and GNAME77908(G77908,G77906,G77909);
  nand GNAME77909(G77909,G80,G77911);
  buf GNAME77910(G77910,G77906);
  buf GNAME77911(G77911,G77901);
  dff DFF_77920(CK,G77919,G68070);
  and GNAME77921(G77921,G77919,G77922);
  nand GNAME77922(G77922,G80,G77924);
  buf GNAME77923(G77923,G77919);
  buf GNAME77924(G77924,G77914);
  dff DFF_77933(CK,G77932,G73841);
  and GNAME77934(G77934,G77932,G77935);
  nand GNAME77935(G77935,G80,G77937);
  buf GNAME77936(G77936,G77932);
  buf GNAME77937(G77937,G77927);
  dff DFF_77946(CK,G77945,G77837);
  and GNAME77947(G77947,G77945,G77948);
  nand GNAME77948(G77948,G80,G77950);
  buf GNAME77949(G77949,G77945);
  buf GNAME77950(G77950,G77940);
  dff DFF_77959(CK,G77958,G77866);
  and GNAME77960(G77960,G77958,G77961);
  nand GNAME77961(G77961,G80,G77963);
  buf GNAME77962(G77962,G77958);
  buf GNAME77963(G77963,G77953);
  dff DFF_77972(CK,G77971,G70365);
  and GNAME77973(G77973,G77971,G77974);
  nand GNAME77974(G77974,G80,G77976);
  buf GNAME77975(G77975,G77971);
  buf GNAME77976(G77976,G77966);
  dff DFF_77985(CK,G77984,G72060);
  and GNAME77986(G77986,G77984,G77987);
  nand GNAME77987(G77987,G80,G77989);
  buf GNAME77988(G77988,G77984);
  buf GNAME77989(G77989,G77979);
  dff DFF_77998(CK,G77997,G70350);
  and GNAME77999(G77999,G77997,G78000);
  nand GNAME78000(G78000,G80,G78002);
  buf GNAME78001(G78001,G77997);
  buf GNAME78002(G78002,G77992);
  dff DFF_78011(CK,G78010,G72045);
  and GNAME78012(G78012,G78010,G78013);
  nand GNAME78013(G78013,G80,G78015);
  buf GNAME78014(G78014,G78010);
  buf GNAME78015(G78015,G78005);
  dff DFF_78024(CK,G78023,G72480);
  and GNAME78025(G78025,G78023,G78026);
  nand GNAME78026(G78026,G80,G78028);
  buf GNAME78027(G78027,G78023);
  buf GNAME78028(G78028,G78018);
  dff DFF_78037(CK,G78036,G72945);
  and GNAME78038(G78038,G78036,G78039);
  nand GNAME78039(G78039,G80,G78041);
  buf GNAME78040(G78040,G78036);
  buf GNAME78041(G78041,G78031);
  dff DFF_78050(CK,G78049,G72495);
  and GNAME78051(G78051,G78049,G78052);
  nand GNAME78052(G78052,G80,G78054);
  buf GNAME78053(G78053,G78049);
  buf GNAME78054(G78054,G78044);
  dff DFF_78063(CK,G78062,G73838);
  and GNAME78064(G78064,G78062,G78065);
  nand GNAME78065(G78065,G80,G78067);
  buf GNAME78066(G78066,G78062);
  buf GNAME78067(G78067,G78057);
  dff DFF_78076(CK,G78075,G72030);
  and GNAME78077(G78077,G78075,G78078);
  nand GNAME78078(G78078,G80,G78080);
  buf GNAME78079(G78079,G78075);
  buf GNAME78080(G78080,G78070);
  dff DFF_78089(CK,G78088,G72015);
  and GNAME78090(G78090,G78088,G78091);
  nand GNAME78091(G78091,G80,G78093);
  buf GNAME78092(G78092,G78088);
  buf GNAME78093(G78093,G78083);
  dff DFF_78102(CK,G78101,G72000);
  and GNAME78103(G78103,G78101,G78104);
  nand GNAME78104(G78104,G80,G78106);
  buf GNAME78105(G78105,G78101);
  buf GNAME78106(G78106,G78096);
  dff DFF_78115(CK,G78114,G71985);
  and GNAME78116(G78116,G78114,G78117);
  nand GNAME78117(G78117,G80,G78119);
  buf GNAME78118(G78118,G78114);
  buf GNAME78119(G78119,G78109);
  dff DFF_78128(CK,G78127,G72960);
  and GNAME78129(G78129,G78127,G78130);
  nand GNAME78130(G78130,G80,G78132);
  buf GNAME78131(G78131,G78127);
  buf GNAME78132(G78132,G78122);
  dff DFF_78141(CK,G78140,G72975);
  and GNAME78142(G78142,G78140,G78143);
  nand GNAME78143(G78143,G80,G78145);
  buf GNAME78144(G78144,G78140);
  buf GNAME78145(G78145,G78135);
  dff DFF_78154(CK,G78153,G72990);
  and GNAME78155(G78155,G78153,G78156);
  nand GNAME78156(G78156,G80,G78158);
  buf GNAME78157(G78157,G78153);
  buf GNAME78158(G78158,G78148);
  dff DFF_78167(CK,G78166,G73035);
  and GNAME78168(G78168,G78166,G78169);
  nand GNAME78169(G78169,G80,G78171);
  buf GNAME78170(G78170,G78166);
  buf GNAME78171(G78171,G78161);
  dff DFF_78180(CK,G78179,G73835);
  and GNAME78181(G78181,G78179,G78182);
  nand GNAME78182(G78182,G80,G78184);
  buf GNAME78183(G78183,G78179);
  buf GNAME78184(G78184,G78174);
  dff DFF_78193(CK,G78192,G73832);
  and GNAME78194(G78194,G78192,G78195);
  nand GNAME78195(G78195,G80,G78197);
  buf GNAME78196(G78196,G78192);
  buf GNAME78197(G78197,G78187);
  dff DFF_78206(CK,G78205,G71970);
  and GNAME78207(G78207,G78205,G78208);
  nand GNAME78208(G78208,G80,G78210);
  buf GNAME78209(G78209,G78205);
  buf GNAME78210(G78210,G78200);
  dff DFF_78219(CK,G78218,G71955);
  and GNAME78220(G78220,G78218,G78221);
  nand GNAME78221(G78221,G80,G78223);
  buf GNAME78222(G78222,G78218);
  buf GNAME78223(G78223,G78213);
  dff DFF_78232(CK,G78231,G71940);
  and GNAME78233(G78233,G78231,G78234);
  nand GNAME78234(G78234,G80,G78236);
  buf GNAME78235(G78235,G78231);
  buf GNAME78236(G78236,G78226);
  dff DFF_78245(CK,G78244,G71925);
  and GNAME78246(G78246,G78244,G78247);
  nand GNAME78247(G78247,G80,G78249);
  buf GNAME78248(G78248,G78244);
  buf GNAME78249(G78249,G78239);
  dff DFF_78258(CK,G78257,G73005);
  and GNAME78259(G78259,G78257,G78260);
  nand GNAME78260(G78260,G80,G78262);
  buf GNAME78261(G78261,G78257);
  buf GNAME78262(G78262,G78252);
  dff DFF_78271(CK,G78270,G73020);
  and GNAME78272(G78272,G78270,G78273);
  nand GNAME78273(G78273,G80,G78275);
  buf GNAME78274(G78274,G78270);
  buf GNAME78275(G78275,G78265);
  dff DFF_78284(CK,G78283,G73050);
  and GNAME78285(G78285,G78283,G78286);
  nand GNAME78286(G78286,G80,G78288);
  buf GNAME78287(G78287,G78283);
  buf GNAME78288(G78288,G78278);
  dff DFF_78297(CK,G78296,G73095);
  and GNAME78298(G78298,G78296,G78299);
  nand GNAME78299(G78299,G80,G78301);
  buf GNAME78300(G78300,G78296);
  buf GNAME78301(G78301,G78291);
  dff DFF_78310(CK,G78309,G73829);
  and GNAME78311(G78311,G78309,G78312);
  nand GNAME78312(G78312,G80,G78314);
  buf GNAME78313(G78313,G78309);
  buf GNAME78314(G78314,G78304);
  dff DFF_78323(CK,G78322,G73850);
  and GNAME78324(G78324,G78322,G78325);
  nand GNAME78325(G78325,G80,G78327);
  buf GNAME78326(G78326,G78322);
  buf GNAME78327(G78327,G78317);
  dff DFF_78336(CK,G78335,G71910);
  and GNAME78337(G78337,G78335,G78338);
  nand GNAME78338(G78338,G80,G78340);
  buf GNAME78339(G78339,G78335);
  buf GNAME78340(G78340,G78330);
  dff DFF_78349(CK,G78348,G71895);
  and GNAME78350(G78350,G78348,G78351);
  nand GNAME78351(G78351,G80,G78353);
  buf GNAME78352(G78352,G78348);
  buf GNAME78353(G78353,G78343);
  dff DFF_78362(CK,G78361,G71880);
  and GNAME78363(G78363,G78361,G78364);
  nand GNAME78364(G78364,G80,G78366);
  buf GNAME78365(G78365,G78361);
  buf GNAME78366(G78366,G78356);
  dff DFF_78375(CK,G78374,G71865);
  and GNAME78376(G78376,G78374,G78377);
  nand GNAME78377(G78377,G80,G78379);
  buf GNAME78378(G78378,G78374);
  buf GNAME78379(G78379,G78369);
  dff DFF_78388(CK,G78387,G73065);
  and GNAME78389(G78389,G78387,G78390);
  nand GNAME78390(G78390,G80,G78392);
  buf GNAME78391(G78391,G78387);
  buf GNAME78392(G78392,G78382);
  dff DFF_78401(CK,G78400,G73080);
  and GNAME78402(G78402,G78400,G78403);
  nand GNAME78403(G78403,G80,G78405);
  buf GNAME78404(G78404,G78400);
  buf GNAME78405(G78405,G78395);
  dff DFF_78414(CK,G78413,G73110);
  and GNAME78415(G78415,G78413,G78416);
  nand GNAME78416(G78416,G80,G78418);
  buf GNAME78417(G78417,G78413);
  buf GNAME78418(G78418,G78408);
  dff DFF_78427(CK,G78426,G73155);
  and GNAME78428(G78428,G78426,G78429);
  nand GNAME78429(G78429,G80,G78431);
  buf GNAME78430(G78430,G78426);
  buf GNAME78431(G78431,G78421);
  dff DFF_78440(CK,G78439,G73847);
  and GNAME78441(G78441,G78439,G78442);
  nand GNAME78442(G78442,G80,G78444);
  buf GNAME78443(G78443,G78439);
  buf GNAME78444(G78444,G78434);
  dff DFF_78453(CK,G78452,G73844);
  and GNAME78454(G78454,G78452,G78455);
  nand GNAME78455(G78455,G80,G78457);
  buf GNAME78456(G78456,G78452);
  buf GNAME78457(G78457,G78447);
  dff DFF_78466(CK,G78465,G71850);
  and GNAME78467(G78467,G78465,G78468);
  nand GNAME78468(G78468,G80,G78470);
  buf GNAME78469(G78469,G78465);
  buf GNAME78470(G78470,G78460);
  dff DFF_78479(CK,G78478,G72420);
  and GNAME78480(G78480,G78478,G78481);
  nand GNAME78481(G78481,G80,G78483);
  buf GNAME78482(G78482,G78478);
  buf GNAME78483(G78483,G78473);
  dff DFF_78492(CK,G78491,G71835);
  and GNAME78493(G78493,G78491,G78494);
  nand GNAME78494(G78494,G80,G78496);
  buf GNAME78495(G78495,G78491);
  buf GNAME78496(G78496,G78486);
  dff DFF_78505(CK,G78504,G72405);
  and GNAME78506(G78506,G78504,G78507);
  nand GNAME78507(G78507,G80,G78509);
  buf GNAME78508(G78508,G78504);
  buf GNAME78509(G78509,G78499);
  dff DFF_78518(CK,G78517,G73125);
  and GNAME78519(G78519,G78517,G78520);
  nand GNAME78520(G78520,G80,G78522);
  buf GNAME78521(G78521,G78517);
  buf GNAME78522(G78522,G78512);
  dff DFF_78531(CK,G78530,G73140);
  and GNAME78532(G78532,G78530,G78533);
  nand GNAME78533(G78533,G80,G78535);
  buf GNAME78534(G78534,G78530);
  buf GNAME78535(G78535,G78525);
  dff DFF_78544(CK,G78543,G73170);
  and GNAME78545(G78545,G78543,G78546);
  nand GNAME78546(G78546,G80,G78548);
  buf GNAME78547(G78547,G78543);
  buf GNAME78548(G78548,G78538);
  dff DFF_78557(CK,G78556,G73185);
  and GNAME78558(G78558,G78556,G78559);
  nand GNAME78559(G78559,G80,G78561);
  buf GNAME78560(G78560,G78556);
  buf GNAME78561(G78561,G78551);
  dff DFF_78570(CK,G78569,G73853);
  and GNAME78571(G78571,G78569,G78572);
  nand GNAME78572(G78572,G80,G78574);
  buf GNAME78573(G78573,G78569);
  buf GNAME78574(G78574,G78564);
  dff DFF_78583(CK,G78582,G73856);
  and GNAME78584(G78584,G78582,G78585);
  nand GNAME78585(G78585,G80,G78587);
  buf GNAME78586(G78586,G78582);
  buf GNAME78587(G78587,G78577);
  dff DFF_78596(CK,G78595,G72390);
  and GNAME78597(G78597,G78595,G78598);
  nand GNAME78598(G78598,G80,G78600);
  buf GNAME78599(G78599,G78595);
  buf GNAME78600(G78600,G78590);
  dff DFF_78609(CK,G78608,G72375);
  and GNAME78610(G78610,G78608,G78611);
  nand GNAME78611(G78611,G80,G78613);
  buf GNAME78612(G78612,G78608);
  buf GNAME78613(G78613,G78603);
  dff DFF_78622(CK,G78621,G72360);
  and GNAME78623(G78623,G78621,G78624);
  nand GNAME78624(G78624,G80,G78626);
  buf GNAME78625(G78625,G78621);
  buf GNAME78626(G78626,G78616);
  dff DFF_78635(CK,G78634,G72345);
  and GNAME78636(G78636,G78634,G78637);
  nand GNAME78637(G78637,G80,G78639);
  buf GNAME78638(G78638,G78634);
  buf GNAME78639(G78639,G78629);
  dff DFF_78648(CK,G78647,G73200);
  and GNAME78649(G78649,G78647,G78650);
  nand GNAME78650(G78650,G80,G78652);
  buf GNAME78651(G78651,G78647);
  buf GNAME78652(G78652,G78642);
  dff DFF_78661(CK,G78660,G73215);
  and GNAME78662(G78662,G78660,G78663);
  nand GNAME78663(G78663,G80,G78665);
  buf GNAME78664(G78664,G78660);
  buf GNAME78665(G78665,G78655);
  dff DFF_78674(CK,G78673,G73230);
  and GNAME78675(G78675,G78673,G78676);
  nand GNAME78676(G78676,G80,G78678);
  buf GNAME78677(G78677,G78673);
  buf GNAME78678(G78678,G78668);
  dff DFF_78687(CK,G78686,G73245);
  and GNAME78688(G78688,G78686,G78689);
  nand GNAME78689(G78689,G80,G78691);
  buf GNAME78690(G78690,G78686);
  buf GNAME78691(G78691,G78681);
  dff DFF_78700(CK,G78699,G73868);
  and GNAME78701(G78701,G78699,G78702);
  nand GNAME78702(G78702,G80,G78704);
  buf GNAME78703(G78703,G78699);
  buf GNAME78704(G78704,G78694);
  dff DFF_78713(CK,G78712,G73865);
  and GNAME78714(G78714,G78712,G78715);
  nand GNAME78715(G78715,G80,G78717);
  buf GNAME78716(G78716,G78712);
  buf GNAME78717(G78717,G78707);
  dff DFF_78726(CK,G78725,G72330);
  and GNAME78727(G78727,G78725,G78728);
  nand GNAME78728(G78728,G80,G78730);
  buf GNAME78729(G78729,G78725);
  buf GNAME78730(G78730,G78720);
  dff DFF_78739(CK,G78738,G72315);
  and GNAME78740(G78740,G78738,G78741);
  nand GNAME78741(G78741,G80,G78743);
  buf GNAME78742(G78742,G78738);
  buf GNAME78743(G78743,G78733);
  dff DFF_78752(CK,G78751,G72300);
  and GNAME78753(G78753,G78751,G78754);
  nand GNAME78754(G78754,G80,G78756);
  buf GNAME78755(G78755,G78751);
  buf GNAME78756(G78756,G78746);
  dff DFF_78765(CK,G78764,G72285);
  and GNAME78766(G78766,G78764,G78767);
  nand GNAME78767(G78767,G80,G78769);
  buf GNAME78768(G78768,G78764);
  buf GNAME78769(G78769,G78759);
  dff DFF_78778(CK,G78777,G73260);
  and GNAME78779(G78779,G78777,G78780);
  nand GNAME78780(G78780,G80,G78782);
  buf GNAME78781(G78781,G78777);
  buf GNAME78782(G78782,G78772);
  dff DFF_78791(CK,G78790,G73275);
  and GNAME78792(G78792,G78790,G78793);
  nand GNAME78793(G78793,G80,G78795);
  buf GNAME78794(G78794,G78790);
  buf GNAME78795(G78795,G78785);
  dff DFF_78804(CK,G78803,G73290);
  and GNAME78805(G78805,G78803,G78806);
  nand GNAME78806(G78806,G80,G78808);
  buf GNAME78807(G78807,G78803);
  buf GNAME78808(G78808,G78798);
  dff DFF_78817(CK,G78816,G73305);
  and GNAME78818(G78818,G78816,G78819);
  nand GNAME78819(G78819,G80,G78821);
  buf GNAME78820(G78820,G78816);
  buf GNAME78821(G78821,G78811);
  dff DFF_78830(CK,G78829,G73862);
  and GNAME78831(G78831,G78829,G78832);
  nand GNAME78832(G78832,G80,G78834);
  buf GNAME78833(G78833,G78829);
  buf GNAME78834(G78834,G78824);
  dff DFF_78843(CK,G78842,G73859);
  and GNAME78844(G78844,G78842,G78845);
  nand GNAME78845(G78845,G80,G78847);
  buf GNAME78846(G78846,G78842);
  buf GNAME78847(G78847,G78837);
  dff DFF_78856(CK,G78855,G72270);
  and GNAME78857(G78857,G78855,G78858);
  nand GNAME78858(G78858,G80,G78860);
  buf GNAME78859(G78859,G78855);
  buf GNAME78860(G78860,G78850);
  dff DFF_78869(CK,G78868,G72255);
  and GNAME78870(G78870,G78868,G78871);
  nand GNAME78871(G78871,G80,G78873);
  buf GNAME78872(G78872,G78868);
  buf GNAME78873(G78873,G78863);
  dff DFF_78882(CK,G78881,G72240);
  and GNAME78883(G78883,G78881,G78884);
  nand GNAME78884(G78884,G80,G78886);
  buf GNAME78885(G78885,G78881);
  buf GNAME78886(G78886,G78876);
  dff DFF_78895(CK,G78894,G72225);
  and GNAME78896(G78896,G78894,G78897);
  nand GNAME78897(G78897,G80,G78899);
  buf GNAME78898(G78898,G78894);
  buf GNAME78899(G78899,G78889);
  dff DFF_78908(CK,G78907,G73320);
  and GNAME78909(G78909,G78907,G78910);
  nand GNAME78910(G78910,G80,G78912);
  buf GNAME78911(G78911,G78907);
  buf GNAME78912(G78912,G78902);
  dff DFF_78921(CK,G78920,G73335);
  and GNAME78922(G78922,G78920,G78923);
  nand GNAME78923(G78923,G80,G78925);
  buf GNAME78924(G78924,G78920);
  buf GNAME78925(G78925,G78915);
  dff DFF_78934(CK,G78933,G73350);
  and GNAME78935(G78935,G78933,G78936);
  nand GNAME78936(G78936,G80,G78938);
  buf GNAME78937(G78937,G78933);
  buf GNAME78938(G78938,G78928);
  dff DFF_78947(CK,G78946,G73365);
  and GNAME78948(G78948,G78946,G78949);
  nand GNAME78949(G78949,G80,G78951);
  buf GNAME78950(G78950,G78946);
  buf GNAME78951(G78951,G78941);
  dff DFF_78960(CK,G78959,G73883);
  and GNAME78961(G78961,G78959,G78962);
  nand GNAME78962(G78962,G80,G78964);
  buf GNAME78963(G78963,G78959);
  buf GNAME78964(G78964,G78954);
  dff DFF_78973(CK,G78972,G73880);
  and GNAME78974(G78974,G78972,G78975);
  nand GNAME78975(G78975,G80,G78977);
  buf GNAME78976(G78976,G78972);
  buf GNAME78977(G78977,G78967);
  dff DFF_78986(CK,G78985,G72210);
  and GNAME78987(G78987,G78985,G78988);
  nand GNAME78988(G78988,G80,G78990);
  buf GNAME78989(G78989,G78985);
  buf GNAME78990(G78990,G78980);
  dff DFF_78999(CK,G78998,G71820);
  and GNAME79000(G79000,G78998,G79001);
  nand GNAME79001(G79001,G80,G79003);
  buf GNAME79002(G79002,G78998);
  buf GNAME79003(G79003,G78993);
  dff DFF_79012(CK,G79011,G72195);
  and GNAME79013(G79013,G79011,G79014);
  nand GNAME79014(G79014,G80,G79016);
  buf GNAME79015(G79015,G79011);
  buf GNAME79016(G79016,G79006);
  dff DFF_79025(CK,G79024,G71805);
  and GNAME79026(G79026,G79024,G79027);
  nand GNAME79027(G79027,G80,G79029);
  buf GNAME79028(G79028,G79024);
  buf GNAME79029(G79029,G79019);
  dff DFF_79038(CK,G79037,G73380);
  and GNAME79039(G79039,G79037,G79040);
  nand GNAME79040(G79040,G80,G79042);
  buf GNAME79041(G79041,G79037);
  buf GNAME79042(G79042,G79032);
  dff DFF_79051(CK,G79050,G73395);
  and GNAME79052(G79052,G79050,G79053);
  nand GNAME79053(G79053,G80,G79055);
  buf GNAME79054(G79054,G79050);
  buf GNAME79055(G79055,G79045);
  dff DFF_79064(CK,G79063,G73410);
  and GNAME79065(G79065,G79063,G79066);
  nand GNAME79066(G79066,G80,G79068);
  buf GNAME79067(G79067,G79063);
  buf GNAME79068(G79068,G79058);
  dff DFF_79077(CK,G79076,G73425);
  and GNAME79078(G79078,G79076,G79079);
  nand GNAME79079(G79079,G80,G79081);
  buf GNAME79080(G79080,G79076);
  buf GNAME79081(G79081,G79071);
  dff DFF_79090(CK,G79089,G73877);
  and GNAME79091(G79091,G79089,G79092);
  nand GNAME79092(G79092,G80,G79094);
  buf GNAME79093(G79093,G79089);
  buf GNAME79094(G79094,G79084);
  dff DFF_79103(CK,G79102,G73874);
  and GNAME79104(G79104,G79102,G79105);
  nand GNAME79105(G79105,G80,G79107);
  buf GNAME79106(G79106,G79102);
  buf GNAME79107(G79107,G79097);
  dff DFF_79116(CK,G79115,G70335);
  and GNAME79117(G79117,G79115,G79118);
  nand GNAME79118(G79118,G80,G79120);
  buf GNAME79119(G79119,G79115);
  buf GNAME79120(G79120,G79110);
  dff DFF_79129(CK,G79128,G71790);
  and GNAME79130(G79130,G79128,G79131);
  nand GNAME79131(G79131,G80,G79133);
  buf GNAME79132(G79132,G79128);
  buf GNAME79133(G79133,G79123);
  dff DFF_79142(CK,G79141,G71775);
  and GNAME79143(G79143,G79141,G79144);
  nand GNAME79144(G79144,G80,G79146);
  buf GNAME79145(G79145,G79141);
  buf GNAME79146(G79146,G79136);
  dff DFF_79155(CK,G79154,G70320);
  and GNAME79156(G79156,G79154,G79157);
  nand GNAME79157(G79157,G80,G79159);
  buf GNAME79158(G79158,G79154);
  buf GNAME79159(G79159,G79149);
  dff DFF_79168(CK,G79167,G71760);
  and GNAME79169(G79169,G79167,G79170);
  nand GNAME79170(G79170,G80,G79172);
  buf GNAME79171(G79171,G79167);
  buf GNAME79172(G79172,G79162);
  dff DFF_79181(CK,G79180,G71745);
  and GNAME79182(G79182,G79180,G79183);
  nand GNAME79183(G79183,G80,G79185);
  buf GNAME79184(G79184,G79180);
  buf GNAME79185(G79185,G79175);
  dff DFF_79194(CK,G79193,G71730);
  and GNAME79195(G79195,G79193,G79196);
  nand GNAME79196(G79196,G80,G79198);
  buf GNAME79197(G79197,G79193);
  buf GNAME79198(G79198,G79188);
  dff DFF_79207(CK,G79206,G71715);
  and GNAME79208(G79208,G79206,G79209);
  nand GNAME79209(G79209,G80,G79211);
  buf GNAME79210(G79210,G79206);
  buf GNAME79211(G79211,G79201);
  dff DFF_79220(CK,G79219,G71700);
  and GNAME79221(G79221,G79219,G79222);
  nand GNAME79222(G79222,G80,G79224);
  buf GNAME79223(G79223,G79219);
  buf GNAME79224(G79224,G79214);
  dff DFF_79233(CK,G79232,G73440);
  and GNAME79234(G79234,G79232,G79235);
  nand GNAME79235(G79235,G80,G79237);
  buf GNAME79236(G79236,G79232);
  buf GNAME79237(G79237,G79227);
  dff DFF_79246(CK,G79245,G73455);
  and GNAME79247(G79247,G79245,G79248);
  nand GNAME79248(G79248,G80,G79250);
  buf GNAME79249(G79249,G79245);
  buf GNAME79250(G79250,G79240);
  dff DFF_79259(CK,G79258,G73485);
  and GNAME79260(G79260,G79258,G79261);
  nand GNAME79261(G79261,G80,G79263);
  buf GNAME79262(G79262,G79258);
  buf GNAME79263(G79263,G79253);
  dff DFF_79272(CK,G79271,G73500);
  and GNAME79273(G79273,G79271,G79274);
  nand GNAME79274(G79274,G80,G79276);
  buf GNAME79275(G79275,G79271);
  buf GNAME79276(G79276,G79266);
  dff DFF_79285(CK,G79284,G73871);
  and GNAME79286(G79286,G79284,G79287);
  nand GNAME79287(G79287,G80,G79289);
  buf GNAME79288(G79288,G79284);
  buf GNAME79289(G79289,G79279);
  dff DFF_79298(CK,G79297,G73895);
  and GNAME79299(G79299,G79297,G79300);
  nand GNAME79300(G79300,G80,G79302);
  buf GNAME79301(G79301,G79297);
  buf GNAME79302(G79302,G79292);
  dff DFF_79311(CK,G79310,G71685);
  and GNAME79312(G79312,G79310,G79313);
  nand GNAME79313(G79313,G80,G79315);
  buf GNAME79314(G79314,G79310);
  buf GNAME79315(G79315,G79305);
  dff DFF_79324(CK,G79323,G71670);
  and GNAME79325(G79325,G79323,G79326);
  nand GNAME79326(G79326,G80,G79328);
  buf GNAME79327(G79327,G79323);
  buf GNAME79328(G79328,G79318);
  dff DFF_79337(CK,G79336,G71655);
  and GNAME79338(G79338,G79336,G79339);
  nand GNAME79339(G79339,G80,G79341);
  buf GNAME79340(G79340,G79336);
  buf GNAME79341(G79341,G79331);
  dff DFF_79350(CK,G79349,G71640);
  and GNAME79351(G79351,G79349,G79352);
  nand GNAME79352(G79352,G80,G79354);
  buf GNAME79353(G79353,G79349);
  buf GNAME79354(G79354,G79344);
  dff DFF_79363(CK,G79362,G71625);
  and GNAME79364(G79364,G79362,G79365);
  nand GNAME79365(G79365,G80,G79367);
  buf GNAME79366(G79366,G79362);
  buf GNAME79367(G79367,G79357);
  dff DFF_79376(CK,G79375,G71610);
  and GNAME79377(G79377,G79375,G79378);
  nand GNAME79378(G79378,G80,G79380);
  buf GNAME79379(G79379,G79375);
  buf GNAME79380(G79380,G79370);
  dff DFF_79389(CK,G79388,G71595);
  and GNAME79390(G79390,G79388,G79391);
  nand GNAME79391(G79391,G80,G79393);
  buf GNAME79392(G79392,G79388);
  buf GNAME79393(G79393,G79383);
  dff DFF_79402(CK,G79401,G71580);
  and GNAME79403(G79403,G79401,G79404);
  nand GNAME79404(G79404,G80,G79406);
  buf GNAME79405(G79405,G79401);
  buf GNAME79406(G79406,G79396);
  dff DFF_79415(CK,G79414,G73470);
  and GNAME79416(G79416,G79414,G79417);
  nand GNAME79417(G79417,G80,G79419);
  buf GNAME79418(G79418,G79414);
  buf GNAME79419(G79419,G79409);
  dff DFF_79428(CK,G79427,G73515);
  and GNAME79429(G79429,G79427,G79430);
  nand GNAME79430(G79430,G80,G79432);
  buf GNAME79431(G79431,G79427);
  buf GNAME79432(G79432,G79422);
  dff DFF_79441(CK,G79440,G73530);
  and GNAME79442(G79442,G79440,G79443);
  nand GNAME79443(G79443,G80,G79445);
  buf GNAME79444(G79444,G79440);
  buf GNAME79445(G79445,G79435);
  dff DFF_79454(CK,G79453,G73545);
  and GNAME79455(G79455,G79453,G79456);
  nand GNAME79456(G79456,G80,G79458);
  buf GNAME79457(G79457,G79453);
  buf GNAME79458(G79458,G79448);
  dff DFF_79467(CK,G79466,G73560);
  and GNAME79468(G79468,G79466,G79469);
  nand GNAME79469(G79469,G80,G79471);
  buf GNAME79470(G79470,G79466);
  buf GNAME79471(G79471,G79461);
  dff DFF_79480(CK,G79479,G73892);
  and GNAME79481(G79481,G79479,G79482);
  nand GNAME79482(G79482,G80,G79484);
  buf GNAME79483(G79483,G79479);
  buf GNAME79484(G79484,G79474);
  dff DFF_79493(CK,G79492,G73889);
  and GNAME79494(G79494,G79492,G79495);
  nand GNAME79495(G79495,G80,G79497);
  buf GNAME79496(G79496,G79492);
  buf GNAME79497(G79497,G79487);
  dff DFF_79506(CK,G79505,G71565);
  and GNAME79507(G79507,G79505,G79508);
  nand GNAME79508(G79508,G80,G79510);
  buf GNAME79509(G79509,G79505);
  buf GNAME79510(G79510,G79500);
  dff DFF_79519(CK,G79518,G71550);
  and GNAME79520(G79520,G79518,G79521);
  nand GNAME79521(G79521,G80,G79523);
  buf GNAME79522(G79522,G79518);
  buf GNAME79523(G79523,G79513);
  dff DFF_79532(CK,G79531,G71535);
  and GNAME79533(G79533,G79531,G79534);
  nand GNAME79534(G79534,G80,G79536);
  buf GNAME79535(G79535,G79531);
  buf GNAME79536(G79536,G79526);
  dff DFF_79545(CK,G79544,G72180);
  and GNAME79546(G79546,G79544,G79547);
  nand GNAME79547(G79547,G80,G79549);
  buf GNAME79548(G79548,G79544);
  buf GNAME79549(G79549,G79539);
  dff DFF_79558(CK,G79557,G72165);
  and GNAME79559(G79559,G79557,G79560);
  nand GNAME79560(G79560,G80,G79562);
  buf GNAME79561(G79561,G79557);
  buf GNAME79562(G79562,G79552);
  dff DFF_79571(CK,G79570,G72150);
  and GNAME79572(G79572,G79570,G79573);
  nand GNAME79573(G79573,G80,G79575);
  buf GNAME79574(G79574,G79570);
  buf GNAME79575(G79575,G79565);
  dff DFF_79584(CK,G79583,G72135);
  and GNAME79585(G79585,G79583,G79586);
  nand GNAME79586(G79586,G80,G79588);
  buf GNAME79587(G79587,G79583);
  buf GNAME79588(G79588,G79578);
  dff DFF_79597(CK,G79596,G71520);
  and GNAME79598(G79598,G79596,G79599);
  nand GNAME79599(G79599,G80,G79601);
  buf GNAME79600(G79600,G79596);
  buf GNAME79601(G79601,G79591);
  dff DFF_79610(CK,G79609,G71505);
  and GNAME79611(G79611,G79609,G79612);
  nand GNAME79612(G79612,G80,G79614);
  buf GNAME79613(G79613,G79609);
  buf GNAME79614(G79614,G79604);
  dff DFF_79623(CK,G79622,G73575);
  and GNAME79624(G79624,G79622,G79625);
  nand GNAME79625(G79625,G80,G79627);
  buf GNAME79626(G79626,G79622);
  buf GNAME79627(G79627,G79617);
  dff DFF_79636(CK,G79635,G73590);
  and GNAME79637(G79637,G79635,G79638);
  nand GNAME79638(G79638,G80,G79640);
  buf GNAME79639(G79639,G79635);
  buf GNAME79640(G79640,G79630);
  dff DFF_79649(CK,G79648,G73605);
  and GNAME79650(G79650,G79648,G79651);
  nand GNAME79651(G79651,G80,G79653);
  buf GNAME79652(G79652,G79648);
  buf GNAME79653(G79653,G79643);
  dff DFF_79662(CK,G79661,G73620);
  and GNAME79663(G79663,G79661,G79664);
  nand GNAME79664(G79664,G80,G79666);
  buf GNAME79665(G79665,G79661);
  buf GNAME79666(G79666,G79656);
  dff DFF_79675(CK,G79674,G73886);
  and GNAME79676(G79676,G79674,G79677);
  nand GNAME79677(G79677,G80,G79679);
  buf GNAME79678(G79678,G79674);
  buf GNAME79679(G79679,G79669);
  dff DFF_79688(CK,G79687,G73910);
  and GNAME79689(G79689,G79687,G79690);
  nand GNAME79690(G79690,G80,G79692);
  buf GNAME79691(G79691,G79687);
  buf GNAME79692(G79692,G79682);
  dff DFF_79701(CK,G79700,G71490);
  and GNAME79702(G79702,G79700,G79703);
  nand GNAME79703(G79703,G80,G79705);
  buf GNAME79704(G79704,G79700);
  buf GNAME79705(G79705,G79695);
  dff DFF_79714(CK,G79713,G71475);
  and GNAME79715(G79715,G79713,G79716);
  nand GNAME79716(G79716,G80,G79718);
  buf GNAME79717(G79717,G79713);
  buf GNAME79718(G79718,G79708);
  dff DFF_79727(CK,G79726,G72120);
  and GNAME79728(G79728,G79726,G79729);
  nand GNAME79729(G79729,G80,G79731);
  buf GNAME79730(G79730,G79726);
  buf GNAME79731(G79731,G79721);
  dff DFF_79740(CK,G79739,G72105);
  and GNAME79741(G79741,G79739,G79742);
  nand GNAME79742(G79742,G80,G79744);
  buf GNAME79743(G79743,G79739);
  buf GNAME79744(G79744,G79734);
  dff DFF_79753(CK,G79752,G72090);
  and GNAME79754(G79754,G79752,G79755);
  nand GNAME79755(G79755,G80,G79757);
  buf GNAME79756(G79756,G79752);
  buf GNAME79757(G79757,G79747);
  dff DFF_79766(CK,G79765,G72075);
  and GNAME79767(G79767,G79765,G79768);
  nand GNAME79768(G79768,G80,G79770);
  buf GNAME79769(G79769,G79765);
  buf GNAME79770(G79770,G79760);
  dff DFF_79779(CK,G79778,G71460);
  and GNAME79780(G79780,G79778,G79781);
  nand GNAME79781(G79781,G80,G79783);
  buf GNAME79782(G79782,G79778);
  buf GNAME79783(G79783,G79773);
  dff DFF_79792(CK,G79791,G71445);
  and GNAME79793(G79793,G79791,G79794);
  nand GNAME79794(G79794,G80,G79796);
  buf GNAME79795(G79795,G79791);
  buf GNAME79796(G79796,G79786);
  dff DFF_79805(CK,G79804,G73635);
  and GNAME79806(G79806,G79804,G79807);
  nand GNAME79807(G79807,G80,G79809);
  buf GNAME79808(G79808,G79804);
  buf GNAME79809(G79809,G79799);
  dff DFF_79818(CK,G79817,G73650);
  and GNAME79819(G79819,G79817,G79820);
  nand GNAME79820(G79820,G80,G79822);
  buf GNAME79821(G79821,G79817);
  buf GNAME79822(G79822,G79812);
  dff DFF_79831(CK,G79830,G73665);
  and GNAME79832(G79832,G79830,G79833);
  nand GNAME79833(G79833,G80,G79835);
  buf GNAME79834(G79834,G79830);
  buf GNAME79835(G79835,G79825);
  dff DFF_79844(CK,G79843,G73680);
  and GNAME79845(G79845,G79843,G79846);
  nand GNAME79846(G79846,G80,G79848);
  buf GNAME79847(G79847,G79843);
  buf GNAME79848(G79848,G79838);
  dff DFF_79857(CK,G79856,G73907);
  and GNAME79858(G79858,G79856,G79859);
  nand GNAME79859(G79859,G80,G79861);
  buf GNAME79860(G79860,G79856);
  buf GNAME79861(G79861,G79851);
  dff DFF_79870(CK,G79869,G73904);
  and GNAME79871(G79871,G79869,G79872);
  nand GNAME79872(G79872,G80,G79874);
  buf GNAME79873(G79873,G79869);
  buf GNAME79874(G79874,G79864);
  dff DFF_79883(CK,G79882,G70305);
  and GNAME79884(G79884,G79882,G79885);
  nand GNAME79885(G79885,G80,G79887);
  buf GNAME79886(G79886,G79882);
  buf GNAME79887(G79887,G79877);
  dff DFF_79896(CK,G79895,G70290);
  and GNAME79897(G79897,G79895,G79898);
  nand GNAME79898(G79898,G80,G79900);
  buf GNAME79899(G79899,G79895);
  buf GNAME79900(G79900,G79890);
  dff DFF_79909(CK,G79908,G71430);
  and GNAME79910(G79910,G79908,G79911);
  nand GNAME79911(G79911,G80,G79913);
  buf GNAME79912(G79912,G79908);
  buf GNAME79913(G79913,G79903);
  dff DFF_79922(CK,G79921,G71415);
  and GNAME79923(G79923,G79921,G79924);
  nand GNAME79924(G79924,G80,G79926);
  buf GNAME79925(G79925,G79921);
  buf GNAME79926(G79926,G79916);
  dff DFF_79935(CK,G79934,G71400);
  and GNAME79936(G79936,G79934,G79937);
  nand GNAME79937(G79937,G80,G79939);
  buf GNAME79938(G79938,G79934);
  buf GNAME79939(G79939,G79929);
  dff DFF_79948(CK,G79947,G71385);
  and GNAME79949(G79949,G79947,G79950);
  nand GNAME79950(G79950,G80,G79952);
  buf GNAME79951(G79951,G79947);
  buf GNAME79952(G79952,G79942);
  dff DFF_79961(CK,G79960,G71370);
  and GNAME79962(G79962,G79960,G79963);
  nand GNAME79963(G79963,G80,G79965);
  buf GNAME79964(G79964,G79960);
  buf GNAME79965(G79965,G79955);
  dff DFF_79974(CK,G79973,G70275);
  and GNAME79975(G79975,G79973,G79976);
  nand GNAME79976(G79976,G80,G79978);
  buf GNAME79977(G79977,G79973);
  buf GNAME79978(G79978,G79968);
  dff DFF_79987(CK,G79986,G70260);
  and GNAME79988(G79988,G79986,G79989);
  nand GNAME79989(G79989,G80,G79991);
  buf GNAME79990(G79990,G79986);
  buf GNAME79991(G79991,G79981);
  dff DFF_80000(CK,G79999,G73695);
  and GNAME80001(G80001,G79999,G80002);
  nand GNAME80002(G80002,G80,G80004);
  buf GNAME80003(G80003,G79999);
  buf GNAME80004(G80004,G79994);
  dff DFF_80013(CK,G80012,G73710);
  and GNAME80014(G80014,G80012,G80015);
  nand GNAME80015(G80015,G80,G80017);
  buf GNAME80016(G80016,G80012);
  buf GNAME80017(G80017,G80007);
  dff DFF_80026(CK,G80025,G73725);
  and GNAME80027(G80027,G80025,G80028);
  nand GNAME80028(G80028,G80,G80030);
  buf GNAME80029(G80029,G80025);
  buf GNAME80030(G80030,G80020);
  dff DFF_80039(CK,G80038,G73740);
  and GNAME80040(G80040,G80038,G80041);
  nand GNAME80041(G80041,G80,G80043);
  buf GNAME80042(G80042,G80038);
  buf GNAME80043(G80043,G80033);
  dff DFF_80052(CK,G80051,G73901);
  and GNAME80053(G80053,G80051,G80054);
  nand GNAME80054(G80054,G80,G80056);
  buf GNAME80055(G80055,G80051);
  buf GNAME80056(G80056,G80046);
  dff DFF_80065(CK,G80064,G73898);
  and GNAME80066(G80066,G80064,G80067);
  nand GNAME80067(G80067,G80,G80069);
  buf GNAME80068(G80068,G80064);
  buf GNAME80069(G80069,G80059);
  dff DFF_80078(CK,G80077,G70245);
  and GNAME80079(G80079,G80077,G80080);
  nand GNAME80080(G80080,G80,G80082);
  buf GNAME80081(G80081,G80077);
  buf GNAME80082(G80082,G80072);
  dff DFF_80091(CK,G80090,G70440);
  and GNAME80092(G80092,G80090,G80093);
  nand GNAME80093(G80093,G80,G80095);
  buf GNAME80094(G80094,G80090);
  buf GNAME80095(G80095,G80085);
  dff DFF_80104(CK,G80103,G71355);
  and GNAME80105(G80105,G80103,G80106);
  nand GNAME80106(G80106,G80,G80108);
  buf GNAME80107(G80107,G80103);
  buf GNAME80108(G80108,G80098);
  dff DFF_80117(CK,G80116,G71340);
  and GNAME80118(G80118,G80116,G80119);
  nand GNAME80119(G80119,G80,G80121);
  buf GNAME80120(G80120,G80116);
  buf GNAME80121(G80121,G80111);
  dff DFF_80130(CK,G80129,G71325);
  and GNAME80131(G80131,G80129,G80132);
  nand GNAME80132(G80132,G80,G80134);
  buf GNAME80133(G80133,G80129);
  buf GNAME80134(G80134,G80124);
  dff DFF_80143(CK,G80142,G71310);
  and GNAME80144(G80144,G80142,G80145);
  nand GNAME80145(G80145,G80,G80147);
  buf GNAME80146(G80146,G80142);
  buf GNAME80147(G80147,G80137);
  dff DFF_80156(CK,G80155,G70230);
  and GNAME80157(G80157,G80155,G80158);
  nand GNAME80158(G80158,G80,G80160);
  buf GNAME80159(G80159,G80155);
  buf GNAME80160(G80160,G80150);
  dff DFF_80169(CK,G80168,G70425);
  and GNAME80170(G80170,G80168,G80171);
  nand GNAME80171(G80171,G80,G80173);
  buf GNAME80172(G80172,G80168);
  buf GNAME80173(G80173,G80163);
  dff DFF_80182(CK,G80181,G73755);
  and GNAME80183(G80183,G80181,G80184);
  nand GNAME80184(G80184,G80,G80186);
  buf GNAME80185(G80185,G80181);
  buf GNAME80186(G80186,G80176);
  dff DFF_80195(CK,G80194,G72450);
  and GNAME80196(G80196,G80194,G80197);
  nand GNAME80197(G80197,G80,G80199);
  buf GNAME80198(G80198,G80194);
  buf GNAME80199(G80199,G80189);
  dff DFF_80208(CK,G80207,G73770);
  and GNAME80209(G80209,G80207,G80210);
  nand GNAME80210(G80210,G80,G80212);
  buf GNAME80211(G80211,G80207);
  buf GNAME80212(G80212,G80202);
  dff DFF_80221(CK,G80220,G73785);
  and GNAME80222(G80222,G80220,G80223);
  nand GNAME80223(G80223,G80,G80225);
  buf GNAME80224(G80224,G80220);
  buf GNAME80225(G80225,G80215);
  dff DFF_80234(CK,G80233,G73922);
  and GNAME80235(G80235,G80233,G80236);
  nand GNAME80236(G80236,G80,G80238);
  buf GNAME80237(G80237,G80233);
  buf GNAME80238(G80238,G80228);
  dff DFF_80247(CK,G80246,G73919);
  and GNAME80248(G80248,G80246,G80249);
  nand GNAME80249(G80249,G80,G80251);
  buf GNAME80250(G80250,G80246);
  buf GNAME80251(G80251,G80241);
  dff DFF_80260(CK,G80259,G68040);
  and GNAME80261(G80261,G80259,G80262);
  nand GNAME80262(G80262,G80,G80264);
  buf GNAME80263(G80263,G80259);
  buf GNAME80264(G80264,G80254);
  dff DFF_80273(CK,G80272,G75174);
  and GNAME80274(G80274,G80272,G80275);
  nand GNAME80275(G80275,G80,G80277);
  buf GNAME80276(G80276,G80272);
  buf GNAME80277(G80277,G80267);
  dff DFF_80286(CK,G80285,G74300);
  and GNAME80287(G80287,G80285,G80288);
  nand GNAME80288(G80288,G80,G80290);
  buf GNAME80289(G80289,G80285);
  buf GNAME80290(G80290,G80280);
  dff DFF_80299(CK,G80298,G74297);
  and GNAME80300(G80300,G80298,G80301);
  nand GNAME80301(G80301,G80,G80303);
  buf GNAME80302(G80302,G80298);
  buf GNAME80303(G80303,G80293);
  dff DFF_80312(CK,G80311,G74294);
  and GNAME80313(G80313,G80311,G80314);
  nand GNAME80314(G80314,G80,G80316);
  buf GNAME80315(G80315,G80311);
  buf GNAME80316(G80316,G80306);
  dff DFF_80325(CK,G80324,G74291);
  and GNAME80326(G80326,G80324,G80327);
  nand GNAME80327(G80327,G80,G80329);
  buf GNAME80328(G80328,G80324);
  buf GNAME80329(G80329,G80319);
  dff DFF_80338(CK,G80337,G74288);
  and GNAME80339(G80339,G80337,G80340);
  nand GNAME80340(G80340,G80,G80342);
  buf GNAME80341(G80341,G80337);
  buf GNAME80342(G80342,G80332);
  dff DFF_80351(CK,G80350,G74285);
  and GNAME80352(G80352,G80350,G80353);
  nand GNAME80353(G80353,G80,G80355);
  buf GNAME80354(G80354,G80350);
  buf GNAME80355(G80355,G80345);
  dff DFF_80364(CK,G80363,G74282);
  and GNAME80365(G80365,G80363,G80366);
  nand GNAME80366(G80366,G80,G80368);
  buf GNAME80367(G80367,G80363);
  buf GNAME80368(G80368,G80358);
  dff DFF_80377(CK,G80376,G74234);
  and GNAME80378(G80378,G80376,G80379);
  nand GNAME80379(G80379,G80,G80381);
  buf GNAME80380(G80380,G80376);
  buf GNAME80381(G80381,G80371);
  dff DFF_80390(CK,G80389,G74231);
  and GNAME80391(G80391,G80389,G80392);
  nand GNAME80392(G80392,G80,G80394);
  buf GNAME80393(G80393,G80389);
  buf GNAME80394(G80394,G80384);
  dff DFF_80403(CK,G80402,G74228);
  and GNAME80404(G80404,G80402,G80405);
  nand GNAME80405(G80405,G80,G80407);
  buf GNAME80406(G80406,G80402);
  buf GNAME80407(G80407,G80397);
  dff DFF_80416(CK,G80415,G74225);
  and GNAME80417(G80417,G80415,G80418);
  nand GNAME80418(G80418,G80,G80420);
  buf GNAME80419(G80419,G80415);
  buf GNAME80420(G80420,G80410);
  dff DFF_80429(CK,G80428,G74222);
  and GNAME80430(G80430,G80428,G80431);
  nand GNAME80431(G80431,G80,G80433);
  buf GNAME80432(G80432,G80428);
  buf GNAME80433(G80433,G80423);
  dff DFF_80442(CK,G80441,G74219);
  and GNAME80443(G80443,G80441,G80444);
  nand GNAME80444(G80444,G80,G80446);
  buf GNAME80445(G80445,G80441);
  buf GNAME80446(G80446,G80436);
  dff DFF_80455(CK,G80454,G74216);
  and GNAME80456(G80456,G80454,G80457);
  nand GNAME80457(G80457,G80,G80459);
  buf GNAME80458(G80458,G80454);
  buf GNAME80459(G80459,G80449);
  dff DFF_80468(CK,G80467,G74213);
  and GNAME80469(G80469,G80467,G80470);
  nand GNAME80470(G80470,G80,G80472);
  buf GNAME80471(G80471,G80467);
  buf GNAME80472(G80472,G80462);
  dff DFF_80481(CK,G80480,G74258);
  and GNAME80482(G80482,G80480,G80483);
  nand GNAME80483(G80483,G80,G80485);
  buf GNAME80484(G80484,G80480);
  buf GNAME80485(G80485,G80475);
  dff DFF_80494(CK,G80493,G74255);
  and GNAME80495(G80495,G80493,G80496);
  nand GNAME80496(G80496,G80,G80498);
  buf GNAME80497(G80497,G80493);
  buf GNAME80498(G80498,G80488);
  dff DFF_80507(CK,G80506,G74252);
  and GNAME80508(G80508,G80506,G80509);
  nand GNAME80509(G80509,G80,G80511);
  buf GNAME80510(G80510,G80506);
  buf GNAME80511(G80511,G80501);
  dff DFF_80520(CK,G80519,G74249);
  and GNAME80521(G80521,G80519,G80522);
  nand GNAME80522(G80522,G80,G80524);
  buf GNAME80523(G80523,G80519);
  buf GNAME80524(G80524,G80514);
  dff DFF_80533(CK,G80532,G74246);
  and GNAME80534(G80534,G80532,G80535);
  nand GNAME80535(G80535,G80,G80537);
  buf GNAME80536(G80536,G80532);
  buf GNAME80537(G80537,G80527);
  dff DFF_80546(CK,G80545,G74243);
  and GNAME80547(G80547,G80545,G80548);
  nand GNAME80548(G80548,G80,G80550);
  buf GNAME80549(G80549,G80545);
  buf GNAME80550(G80550,G80540);
  dff DFF_80559(CK,G80558,G74240);
  and GNAME80560(G80560,G80558,G80561);
  nand GNAME80561(G80561,G80,G80563);
  buf GNAME80562(G80562,G80558);
  buf GNAME80563(G80563,G80553);
  dff DFF_80572(CK,G80571,G74237);
  and GNAME80573(G80573,G80571,G80574);
  nand GNAME80574(G80574,G80,G80576);
  buf GNAME80575(G80575,G80571);
  buf GNAME80576(G80576,G80566);
  dff DFF_80585(CK,G80584,G77872);
  and GNAME80586(G80586,G80584,G80587);
  nand GNAME80587(G80587,G80,G80589);
  buf GNAME80588(G80588,G80584);
  buf GNAME80589(G80589,G80579);
  dff DFF_80598(CK,G80597,G77870);
  and GNAME80599(G80599,G80597,G80600);
  nand GNAME80600(G80600,G80,G80602);
  buf GNAME80601(G80601,G80597);
  buf GNAME80602(G80602,G80592);
  dff DFF_80611(CK,G80610,G77868);
  and GNAME80612(G80612,G80610,G80613);
  nand GNAME80613(G80613,G80,G80615);
  buf GNAME80614(G80614,G80610);
  buf GNAME80615(G80615,G80605);
  dff DFF_80624(CK,G80623,G70215);
  and GNAME80625(G80625,G80623,G80626);
  nand GNAME80626(G80626,G80,G80628);
  buf GNAME80627(G80627,G80623);
  buf GNAME80628(G80628,G80618);
  dff DFF_80637(CK,G80636,G70200);
  and GNAME80638(G80638,G80636,G80639);
  nand GNAME80639(G80639,G80,G80641);
  buf GNAME80640(G80640,G80636);
  buf GNAME80641(G80641,G80631);
  dff DFF_80650(CK,G80649,G70185);
  and GNAME80651(G80651,G80649,G80652);
  nand GNAME80652(G80652,G80,G80654);
  buf GNAME80653(G80653,G80649);
  buf GNAME80654(G80654,G80644);
  dff DFF_80663(CK,G80662,G70410);
  and GNAME80664(G80664,G80662,G80665);
  nand GNAME80665(G80665,G80,G80667);
  buf GNAME80666(G80666,G80662);
  buf GNAME80667(G80667,G80657);
  dff DFF_80676(CK,G80675,G73800);
  and GNAME80677(G80677,G80675,G80678);
  nand GNAME80678(G80678,G80,G80680);
  buf GNAME80679(G80679,G80675);
  buf GNAME80680(G80680,G80670);
  dff DFF_80689(CK,G80688,G73815);
  and GNAME80690(G80690,G80688,G80691);
  nand GNAME80691(G80691,G80,G80693);
  buf GNAME80692(G80692,G80688);
  buf GNAME80693(G80693,G80683);
  dff DFF_80702(CK,G80701,G73916);
  and GNAME80703(G80703,G80701,G80704);
  nand GNAME80704(G80704,G80,G80706);
  buf GNAME80705(G80705,G80701);
  buf GNAME80706(G80706,G80696);
  dff DFF_80715(CK,G80714,G73913);
  and GNAME80716(G80716,G80714,G80717);
  nand GNAME80717(G80717,G80,G80719);
  buf GNAME80718(G80718,G80714);
  buf GNAME80719(G80719,G80709);
  dff DFF_80728(CK,G80727,G77841);
  and GNAME80729(G80729,G80727,G80730);
  nand GNAME80730(G80730,G80,G80732);
  buf GNAME80731(G80731,G80727);
  buf GNAME80732(G80732,G80722);
  dff DFF_80741(CK,G80740,G74279);
  and GNAME80742(G80742,G80740,G80743);
  nand GNAME80743(G80743,G80,G80745);
  buf GNAME80744(G80744,G80740);
  buf GNAME80745(G80745,G80735);
  dff DFF_80754(CK,G80753,G74276);
  and GNAME80755(G80755,G80753,G80756);
  nand GNAME80756(G80756,G80,G80758);
  buf GNAME80757(G80757,G80753);
  buf GNAME80758(G80758,G80748);
  dff DFF_80767(CK,G80766,G74273);
  and GNAME80768(G80768,G80766,G80769);
  nand GNAME80769(G80769,G80,G80771);
  buf GNAME80770(G80770,G80766);
  buf GNAME80771(G80771,G80761);
  dff DFF_80780(CK,G80779,G74270);
  and GNAME80781(G80781,G80779,G80782);
  nand GNAME80782(G80782,G80,G80784);
  buf GNAME80783(G80783,G80779);
  buf GNAME80784(G80784,G80774);
  dff DFF_80793(CK,G80792,G74267);
  and GNAME80794(G80794,G80792,G80795);
  nand GNAME80795(G80795,G80,G80797);
  buf GNAME80796(G80796,G80792);
  buf GNAME80797(G80797,G80787);
  dff DFF_80806(CK,G80805,G74264);
  and GNAME80807(G80807,G80805,G80808);
  nand GNAME80808(G80808,G80,G80810);
  buf GNAME80809(G80809,G80805);
  buf GNAME80810(G80810,G80800);
  dff DFF_80819(CK,G80818,G74261);
  and GNAME80820(G80820,G80818,G80821);
  nand GNAME80821(G80821,G80,G80823);
  buf GNAME80822(G80822,G80818);
  buf GNAME80823(G80823,G80813);
  dff DFF_80832(CK,G80831,G80979);
  and GNAME80833(G80833,G80831,G80834);
  nand GNAME80834(G80834,G80,G80836);
  buf GNAME80835(G80835,G80831);
  buf GNAME80836(G80836,G80826);
  dff DFF_80845(CK,G80844,G73820);
  and GNAME80846(G80846,G80844,G80847);
  nand GNAME80847(G80847,G80,G80849);
  buf GNAME80848(G80848,G80844);
  buf GNAME80849(G80849,G80839);
  buf GNAME80850(G80850,G80261);
  buf GNAME80851(G80851,G80261);
  buf GNAME80852(G80852,G2699);
  buf GNAME80853(G80853,G2283);
  buf GNAME80854(G80854,G1867);
  buf GNAME80855(G80855,G10874);
  buf GNAME80856(G80856,G9002);
  buf GNAME80857(G80857,G7130);
  buf GNAME80858(G80858,G2657);
  buf GNAME80859(G80859,G2241);
  buf GNAME80860(G80860,G1825);
  buf GNAME80861(G80861,G10832);
  buf GNAME80862(G80862,G8960);
  buf GNAME80863(G80863,G7088);
  buf GNAME80864(G80864,G10853);
  buf GNAME80865(G80865,G8981);
  buf GNAME80866(G80866,G7109);
  buf GNAME80867(G80867,G2615);
  buf GNAME80868(G80868,G2199);
  buf GNAME80869(G80869,G1783);
  buf GNAME80870(G80870,G10790);
  buf GNAME80871(G80871,G8918);
  buf GNAME80872(G80872,G7046);
  buf GNAME80873(G80873,G10811);
  buf GNAME80874(G80874,G8939);
  buf GNAME80875(G80875,G7067);
  buf GNAME80876(G80876,G2573);
  buf GNAME80877(G80877,G2157);
  buf GNAME80878(G80878,G1741);
  buf GNAME80879(G80879,G10748);
  buf GNAME80880(G80880,G8876);
  buf GNAME80881(G80881,G7004);
  buf GNAME80882(G80882,G10769);
  buf GNAME80883(G80883,G8897);
  buf GNAME80884(G80884,G7025);
  buf GNAME80885(G80885,G2491);
  buf GNAME80886(G80886,G2075);
  buf GNAME80887(G80887,G1659);
  buf GNAME80888(G80888,G10666);
  buf GNAME80889(G80889,G8794);
  buf GNAME80890(G80890,G6922);
  buf GNAME80891(G80891,G10727);
  buf GNAME80892(G80892,G8855);
  buf GNAME80893(G80893,G6983);
  buf GNAME80894(G80894,G2449);
  buf GNAME80895(G80895,G2033);
  buf GNAME80896(G80896,G1617);
  buf GNAME80897(G80897,G10624);
  buf GNAME80898(G80898,G10645);
  buf GNAME80899(G80899,G8752);
  buf GNAME80900(G80900,G8773);
  buf GNAME80901(G80901,G6880);
  buf GNAME80902(G80902,G6901);
  buf GNAME80903(G80903,G2407);
  buf GNAME80904(G80904,G1991);
  buf GNAME80905(G80905,G1575);
  buf GNAME80906(G80906,G77921);
  buf GNAME80907(G80907,G77908);
  buf GNAME80908(G80908,G2699);
  buf GNAME80909(G80909,G2283);
  buf GNAME80910(G80910,G1867);
  buf GNAME80911(G80911,G2657);
  buf GNAME80912(G80912,G2241);
  buf GNAME80913(G80913,G1825);
  buf GNAME80914(G80914,G77921);
  buf GNAME80915(G80915,G77908);
  buf GNAME80916(G80916,G10603);
  buf GNAME80917(G80917,G10582);
  buf GNAME80918(G80918,G10561);
  buf GNAME80919(G80919,G8731);
  buf GNAME80920(G80920,G8710);
  buf GNAME80921(G80921,G6859);
  buf GNAME80922(G80922,G6838);
  buf GNAME80923(G80923,G8689);
  buf GNAME80924(G80924,G6817);
  buf GNAME80925(G80925,G2365);
  buf GNAME80926(G80926,G1949);
  buf GNAME80927(G80927,G1533);
  buf GNAME80928(G80928,G2615);
  buf GNAME80929(G80929,G2199);
  buf GNAME80930(G80930,G1783);
  buf GNAME80931(G80931,G10311);
  buf GNAME80932(G80932,G8439);
  buf GNAME80933(G80933,G6567);
  buf GNAME80934(G80934,G10458);
  buf GNAME80935(G80935,G10519);
  buf GNAME80936(G80936,G8586);
  buf GNAME80937(G80937,G8647);
  buf GNAME80938(G80938,G6714);
  buf GNAME80939(G80939,G6775);
  buf GNAME80940(G80940,G10540);
  buf GNAME80941(G80941,G8668);
  buf GNAME80942(G80942,G6796);
  buf GNAME80943(G80943,G2573);
  buf GNAME80944(G80944,G2157);
  buf GNAME80945(G80945,G1741);
  buf GNAME80946(G80946,G10416);
  buf GNAME80947(G80947,G10395);
  buf GNAME80948(G80948,G10374);
  buf GNAME80949(G80949,G10437);
  buf GNAME80950(G80950,G8565);
  buf GNAME80951(G80951,G6693);
  buf GNAME80952(G80952,G8502);
  buf GNAME80953(G80953,G8523);
  buf GNAME80954(G80954,G8544);
  buf GNAME80955(G80955,G6630);
  buf GNAME80956(G80956,G6651);
  buf GNAME80957(G80957,G6672);
  buf GNAME80958(G80958,G2491);
  buf GNAME80959(G80959,G2075);
  buf GNAME80960(G80960,G1659);
  buf GNAME80961(G80961,G2449);
  buf GNAME80962(G80962,G2033);
  buf GNAME80963(G80963,G1617);
  buf GNAME80964(G80964,G10311);
  buf GNAME80965(G80965,G8439);
  buf GNAME80966(G80966,G6567);
  buf GNAME80967(G80967,G10353);
  buf GNAME80968(G80968,G10332);
  buf GNAME80969(G80969,G8481);
  buf GNAME80970(G80970,G8460);
  buf GNAME80971(G80971,G6609);
  buf GNAME80972(G80972,G6588);
  buf GNAME80973(G80973,G2407);
  buf GNAME80974(G80974,G1991);
  buf GNAME80975(G80975,G1575);
  buf GNAME80976(G80976,G2365);
  buf GNAME80977(G80977,G1949);
  buf GNAME80978(G80978,G1533);
  buf GNAME80979(G80979,G74357);
  buf GNAME80980(G80980,G77813);
  buf GNAME80981(G80981,G77814);
  buf GNAME80982(G80982,G77815);
  buf GNAME80983(G80983,G74357);
  buf GNAME80984(G80984,G74357);
  buf GNAME80985(G80985,G75245);
  buf GNAME80986(G80986,G75246);
  buf GNAME80987(G80987,G75247);
  buf GNAME80988(G80988,G77816);
  buf GNAME80989(G80989,G77817);
  buf GNAME80990(G80990,G77818);
  buf GNAME80991(G80991,G75248);
  buf GNAME80992(G80992,G75249);
  buf GNAME80993(G80993,G75250);
  buf GNAME80994(G80994,G77822);
  buf GNAME80995(G80995,G77819);
  buf GNAME80996(G80996,G77823);
  buf GNAME80997(G80997,G77824);
  buf GNAME80998(G80998,G77820);
  buf GNAME80999(G80999,G77821);
  buf GNAME81000(G81000,G75254);
  buf GNAME81001(G81001,G75255);
  buf GNAME81002(G81002,G75256);
  buf GNAME81003(G81003,G75254);
  buf GNAME81004(G81004,G75251);
  buf GNAME81005(G81005,G75255);
  buf GNAME81006(G81006,G75256);
  buf GNAME81007(G81007,G75252);
  buf GNAME81008(G81008,G75253);
  buf GNAME81009(G81009,G77693);
  buf GNAME81010(G81010,G77694);
  buf GNAME81011(G81011,G77695);
  buf GNAME81012(G81012,G77831);
  buf GNAME81013(G81013,G77832);
  buf GNAME81014(G81014,G77833);
  buf GNAME81015(G81015,G77834);
  buf GNAME81016(G81016,G77835);
  buf GNAME81017(G81017,G77836);
  buf GNAME81018(G81018,G77693);
  buf GNAME81019(G81019,G77694);
  buf GNAME81020(G81020,G77695);
  buf GNAME81021(G81021,G77831);
  buf GNAME81022(G81022,G77832);
  buf GNAME81023(G81023,G77833);
  buf GNAME81024(G81024,G77834);
  buf GNAME81025(G81025,G77835);
  buf GNAME81026(G81026,G77836);
  buf GNAME81027(G81027,G75260);
  buf GNAME81028(G81028,G75263);
  buf GNAME81029(G81029,G75261);
  buf GNAME81030(G81030,G75264);
  buf GNAME81031(G81031,G75262);
  buf GNAME81032(G81032,G75265);
  buf GNAME81033(G81033,G75263);
  buf GNAME81034(G81034,G75264);
  buf GNAME81035(G81035,G75265);
  buf GNAME81036(G81036,G77766);
  buf GNAME81037(G81037,G77767);
  buf GNAME81038(G81038,G77768);
  buf GNAME81039(G81039,G77767);
  buf GNAME81040(G81040,G77766);
  buf GNAME81041(G81041,G77768);
  buf GNAME81042(G81042,G77813);
  buf GNAME81043(G81043,G77816);
  buf GNAME81044(G81044,G77814);
  buf GNAME81045(G81045,G77815);
  buf GNAME81046(G81046,G77817);
  buf GNAME81047(G81047,G77818);
  buf GNAME81048(G81048,G75245);
  buf GNAME81049(G81049,G75246);
  buf GNAME81050(G81050,G75247);
  buf GNAME81051(G81051,G77822);
  buf GNAME81052(G81052,G77823);
  buf GNAME81053(G81053,G77824);
  buf GNAME81054(G81054,G75248);
  buf GNAME81055(G81055,G75249);
  buf GNAME81056(G81056,G75250);
  buf GNAME81057(G81057,G77826);
  buf GNAME81058(G81058,G77827);
  buf GNAME81059(G81059,G77828);
  buf GNAME81060(G81060,G77825);
  buf GNAME81061(G81061,G77829);
  buf GNAME81062(G81062,G77830);
  buf GNAME81063(G81063,G75251);
  buf GNAME81064(G81064,G75252);
  buf GNAME81065(G81065,G75253);
  buf GNAME81066(G81066,G75257);
  buf GNAME81067(G81067,G75258);
  buf GNAME81068(G81068,G75259);
  buf GNAME81069(G81069,G77819);
  buf GNAME81070(G81070,G77820);
  buf GNAME81071(G81071,G77821);
  buf GNAME81072(G81072,G77825);
  buf GNAME81073(G81073,G77829);
  buf GNAME81074(G81074,G77830);
  buf GNAME81075(G81075,G77826);
  buf GNAME81076(G81076,G77827);
  buf GNAME81077(G81077,G77828);
  buf GNAME81078(G81078,G75260);
  buf GNAME81079(G81079,G75261);
  buf GNAME81080(G81080,G75262);
  buf GNAME81081(G81081,G75257);
  buf GNAME81082(G81082,G75258);
  buf GNAME81083(G81083,G75259);

endmodule
