
module b15s_1 ( G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, 
        G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, 
        G29, G30, G31, G32, G33, G34, G35, G36, G21356, G21357, G21358, G21359, 
        G21360, G21361, G21362, G21363, G21364, G21365, G21366, G21367, G21368, 
        G21369, G21370, G21371, G21372, G21373, G21374, G21375, G21376, G21377, 
        G21378, G21379, G21380, G21381, G21382, G21383, G21384, G21385, G21386, 
        G21387, G21388, G21389, G21390, G21391, G21392, G21393, G21394, G21395, 
        G21396, G21397, G21398, G21399, G21400, G21401, G21402, G21403, G21404, 
        G21405, G21406, G21407, G21408, G21409, G21410, G21411, G21412, G21413, 
        G21414, G21415, G21416, G21417, G21418, G21419, G21420, G21421, G21422, 
        G21423, G21424, G21425, G21426, G21427, G21428, G21429, G21430, G21431, 
        G21432, G21433, G21434, G21435, G21436, G21437, G21438, G21439, G21440, 
        G21441, G21442, G21443, G21444, G21445, G21446, G21447, G21448, G21449, 
        G21450, G21451, G21452, G21453, G21454, G21455, G21456, G21457, G21458, 
        G21459, G21460, G21461, G21462, G21463, G21464, G21465, G21466, G21467, 
        G21468, G21469, G21470, G21471, G21472, G21473, G21474, G21475, G21476, 
        G21477, G21478, G21479, G21480, G21481, G21482, G21483, G21484, G21485, 
        G21486, G21487, G21488, G21489, G21490, G21491, G21492, G21493, G21494, 
        G21495, G21496, G21497, G21498, G21499, G21500, G21501, G21502, G21503, 
        G21504, G21505, G21506, G21507, G21508, G21509, G21510, G21511, G21512, 
        G21513, G21514, G21515, G21516, G21517, G21518, G21519, G21520, G21521, 
        G21522, G21523, G21524, G21525, G21526, G21527, G21528, G21529, G21530, 
        G21531, G21532, G21533, G21534, G21535, G21536, G21537, G21538, G21539, 
        G21540, G21541, G21542, G21543, G21544, G21545, G21546, G21547, G21548, 
        G21549, G21550, G21551, G21552, G21553, G21554, G21555, G21556, G21557, 
        G21558, G21559, G21560, G21561, G21562, G21563, G21564, G21565, G21566, 
        G21567, G21568, G21569, G21570, G21571, G21572, G21573, G21574, G21575, 
        G21576, G21577, G21578, G21579, G21580, G21581, G21582, G21583, G21584, 
        G21585, G21586, G21587, G21588, G21589, G21590, G21591, G21592, G21593, 
        G21594, G21595, G21596, G21597, G21598, G21599, G21600, G21601, G21602, 
        G21603, G21604, G21605, G21606, G21607, G21608, G21609, G21610, G21611, 
        G21612, G21613, G21614, G21615, G21616, G21617, G21618, G21619, G21620, 
        G21621, G21622, G21623, G21624, G21625, G21626, G21627, G21628, G21629, 
        G21630, G21631, G21632, G21633, G21634, G21635, G21636, G21637, G21638, 
        G21639, G21640, G21641, G21642, G21643, G21644, G21645, G21646, G21647, 
        G21648, G21649, G21650, G21651, G21652, G21653, G21654, G21655, G21656, 
        G21657, G21658, G21659, G21660, G21661, G21662, G21663, G21664, G21665, 
        G21666, G21667, G21668, G21669, G21670, G21671, G21672, G21673, G21674, 
        G21675, G21676, G21677, G21678, G21679, G21680, G21681, G21682, G21683, 
        G21684, G21685, G21686, G21687, G21688, G21689, G21690, G21691, G21692, 
        G21693, G21694, G21695, G21696, G21697, G21698, G21699, G21700, G21701, 
        G21702, G21703, G21704, G21705, G21706, G21707, G21708, G21709, G21710, 
        G21711, G21712, G21713, G21714, G21715, G21716, G21717, G21718, G21719, 
        G21720, G21721, G21722, G21723, G21724, G21725, G21726, G21727, G21728, 
        G21729, G21730, G21731, G21732, G21733, G21734, G21735, G21736, G21737, 
        G21738, G21739, G21740, G21741, G21742, G21743, G21744, G21745, G21746, 
        G21747, G21748, G21749, G21750, G21751, G21752, G21753, G21754, G21755, 
        G21756, G21757, G21758, G21759, G21760, G21761, G21762, G21763, G21764, 
        G21765, G21766, G21767, G21768, G21769, G21770, G21771, G21772, G21773, 
        G21774, G21775, G21776, G21777, G21778, G21779, G21780, G21781, G21782, 
        G21783, G21784, G21785, G21786, G21787, G21788, G21789, G21790, G21791, 
        G21792, G21793, G21794, G21795, G21796, G21797, G21798, G21799, G21800, 
        G21801, G21802, G21803, G21804, G1732, G1733, G1734, G1735, G757, G758, 
        G759, G760, G761, G762, G763, G764, G765, G766, G767, G768, G769, G770, 
        G771, G772, G773, G774, G775, G776, G777, G778, G779, G780, G781, G782, 
        G783, G784, G785, G786, G787, G789, G790, G1737, G1738, G791, G792, 
        G793, G794, G795, G796, G797, G798, G799, G800, G801, G802, G803, G804, 
        G805, G806, G807, G808, G809, G810, G811, G812, G813, G814, G815, G816, 
        G817, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, 
        G829, G830, G831, G832, G833, G834, G835, G836, G837, G838, G839, G840, 
        G841, G842, G843, G844, G845, G846, G847, G848, G849, G850, G851, G852, 
        G853, G854, G855, G856, G857, G858, G859, G860, G861, G862, G863, G864, 
        G865, G866, G867, G868, G869, G870, G871, G872, G873, G874, G875, G876, 
        G877, G878, G879, G880, G881, G882, G883, G884, G885, G886, G887, G888, 
        G889, G890, G891, G892, G893, G894, G895, G896, G897, G898, G899, G900, 
        G901, G902, G903, G904, G905, G906, G907, G908, G909, G910, G911, G912, 
        G913, G914, G915, G916, G917, G918, G919, G920, G921, G922, G923, G924, 
        G925, G926, G927, G928, G929, G930, G931, G932, G933, G934, G935, G936, 
        G937, G938, G939, G940, G941, G942, G943, G944, G945, G946, G947, G948, 
        G949, G950, G951, G952, G1740, G1742, G1743, G1744, G1745, G953, G954, 
        G955, G956, G1746, G957, G958, G959, G960, G961, G962, G963, G964, 
        G965, G966, G967, G968, G969, G970, G971, G972, G973, G974, G975, G976, 
        G977, G978, G979, G980, G981, G982, G983, G984, G985, G986, G987, G988, 
        G989, G990, G991, G992, G993, G994, G995, G996, G997, G998, G999, 
        G1000, G1001, G1002, G1003, G1004, G1005, G1006, G1007, G1008, G1009, 
        G1010, G1011, G1012, G1013, G1014, G1015, G1016, G1017, G1018, G1019, 
        G1020, G1021, G1022, G1023, G1024, G1025, G1026, G1027, G1028, G1029, 
        G1030, G1031, G1032, G1033, G1034, G1035, G1036, G1037, G1038, G1039, 
        G1040, G1041, G1042, G1043, G1044, G1045, G1046, G1047, G1048, G1049, 
        G1050, G1051, G1052, G1053, G1054, G1055, G1056, G1057, G1058, G1059, 
        G1060, G1061, G1062, G1063, G1064, G1065, G1066, G1067, G1068, G1069, 
        G1070, G1071, G1072, G1073, G1074, G1075, G1076, G1077, G1078, G1079, 
        G1080, G1081, G1082, G1083, G1084, G1085, G1086, G1087, G1088, G1089, 
        G1090, G1091, G1092, G1093, G1094, G1095, G1096, G1097, G1098, G1099, 
        G1100, G1101, G1102, G1103, G1104, G1105, G1106, G1107, G1108, G1109, 
        G1110, G1111, G1112, G1113, G1114, G1115, G1116, G1117, G1118, G1119, 
        G1120, G1121, G1122, G1123, G1124, G1125, G1126, G1127, G1128, G1129, 
        G1130, G1131, G1132, G1133, G1134, G1135, G1136, G1137, G1138, G1139, 
        G1140, G1141, G1142, G1143, G1144, G1145, G1146, G1147, G1148, G1149, 
        G1150, G1151, G1152, G1153, G1154, G1155, G1156, G1157, G1158, G1159, 
        G1160, G1161, G1162, G1163, G1164, G1165, G1166, G1167, G1168, G1169, 
        G1170, G1171, G1172, G1173, G1174, G1175, G1176, G1177, G1178, G1179, 
        G1180, G1181, G1182, G1183, G1747, G1184, G1185, G1186, G1748, G1187, 
        G1749, G1188, G1189, G1750, G1751 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16,
         G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30,
         G31, G32, G33, G34, G35, G36, G21390, G21391, G21392, G21393, G21394,
         G21395, G21396, G21397, G21398, G21399, G21400, G21401, G21402,
         G21403, G21404, G21405, G21406, G21407, G21408, G21409, G21410,
         G21411, G21412, G21413, G21414, G21415, G21416, G21417, G21418,
         G21419, G21420, G21421, G21422, G21423, G21424, G21425, G21426,
         G21427, G21428, G21429, G21430, G21431, G21432, G21433, G21434,
         G21435, G21436, G21437, G21438, G21439, G21440, G21441, G21442,
         G21443, G21444, G21445, G21446, G21447, G21448, G21449, G21450,
         G21451, G21452, G21453, G21454, G21455, G21456, G21457, G21458,
         G21459, G21460, G21461, G21462, G21463, G21464, G21465, G21466,
         G21467, G21468, G21469, G21470, G21471, G21472, G21473, G21474,
         G21475, G21476, G21477, G21478, G21479, G21480, G21481, G21482,
         G21483, G21484, G21485, G21486, G21487, G21488, G21489, G21490,
         G21491, G21492, G21493, G21494, G21495, G21496, G21497, G21498,
         G21499, G21500, G21501, G21502, G21503, G21504, G21505, G21506,
         G21507, G21508, G21509, G21510, G21511, G21512, G21513, G21514,
         G21515, G21516, G21517, G21518, G21519, G21520, G21521, G21522,
         G21523, G21524, G21525, G21526, G21527, G21528, G21529, G21530,
         G21531, G21532, G21533, G21534, G21535, G21536, G21537, G21538,
         G21539, G21540, G21541, G21542, G21543, G21544, G21545, G21546,
         G21547, G21548, G21549, G21550, G21551, G21552, G21553, G21554,
         G21555, G21556, G21557, G21558, G21559, G21560, G21561, G21562,
         G21563, G21564, G21565, G21566, G21567, G21568, G21569, G21570,
         G21571, G21572, G21573, G21574, G21575, G21576, G21577, G21578,
         G21579, G21580, G21581, G21582, G21583, G21584, G21585, G21586,
         G21587, G21588, G21589, G21590, G21591, G21592, G21593, G21594,
         G21595, G21596, G21597, G21598, G21599, G21600, G21601, G21602,
         G21603, G21604, G21605, G21606, G21607, G21608, G21609, G21610,
         G21611, G21612, G21613, G21614, G21615, G21616, G21617, G21618,
         G21619, G21620, G21621, G21622, G21623, G21624, G21625, G21626,
         G21627, G21628, G21629, G21630, G21631, G21632, G21633, G21634,
         G21635, G21636, G21637, G21638, G21639, G21640, G21641, G21642,
         G21643, G21644, G21645, G21646, G21647, G21648, G21649, G21650,
         G21651, G21652, G21653, G21654, G21655, G21656, G21657, G21658,
         G21659, G21660, G21661, G21694, G21695, G21696, G21697, G21698,
         G21699, G21700, G21701, G21702, G21703, G21704, G21705, G21706,
         G21707, G21708, G21709, G21710, G21711, G21712, G21713, G21714,
         G21715, G21716, G21717, G21718, G21719, G21720, G21721, G21722,
         G21723, G21724, G21725, G21726, G21727, G21728, G21729, G21730,
         G21731, G21732, G21733, G21734, G21735, G21736, G21737, G21738,
         G21739, G21740, G21741, G21742, G21743, G21744, G21745, G21746,
         G21747, G21748, G21749, G21750, G21751, G21752, G21753, G21754,
         G21755, G21756, G21757, G21758, G21759, G21760, G21761, G21762,
         G21763, G21764, G21765, G21766, G21767, G21768, G21769, G21770,
         G21771, G21772, G21773, G21774, G21775, G21776, G21777, G21778,
         G21779, G21780, G21781, G21782, G21783, G21784, G21785, G21786,
         G21787, G21788, G21789, G21790, G21791, G21792, G21793, G21795,
         G21796, G21797, G21798, G21801, G21803, G21804;
  output G1732, G1733, G1734, G1735, G757, G758, G759, G760, G761, G762, G763,
         G764, G765, G766, G767, G768, G769, G770, G771, G772, G773, G774,
         G775, G776, G777, G778, G779, G780, G781, G782, G783, G784, G785,
         G786, G787, G789, G790, G1737, G1738, G791, G792, G793, G794, G795,
         G796, G797, G798, G799, G800, G801, G802, G803, G804, G805, G806,
         G807, G808, G809, G810, G811, G812, G813, G814, G815, G816, G817,
         G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828,
         G829, G830, G831, G832, G833, G834, G835, G836, G837, G838, G839,
         G840, G841, G842, G843, G844, G845, G846, G847, G848, G849, G850,
         G851, G852, G853, G854, G855, G856, G857, G858, G859, G860, G861,
         G862, G863, G864, G865, G866, G867, G868, G869, G870, G871, G872,
         G873, G874, G875, G876, G877, G878, G879, G880, G881, G882, G883,
         G884, G885, G886, G887, G888, G889, G890, G891, G892, G893, G894,
         G895, G896, G897, G898, G899, G900, G901, G902, G903, G904, G905,
         G906, G907, G908, G909, G910, G911, G912, G913, G914, G915, G916,
         G917, G918, G919, G920, G921, G922, G923, G924, G925, G926, G927,
         G928, G929, G930, G931, G932, G933, G934, G935, G936, G937, G938,
         G939, G940, G941, G942, G943, G944, G945, G946, G947, G948, G949,
         G950, G951, G952, G1740, G1742, G1743, G1744, G1745, G953, G954, G955,
         G956, G1746, G957, G958, G959, G960, G961, G962, G963, G964, G965,
         G966, G967, G968, G969, G970, G971, G972, G973, G974, G975, G976,
         G977, G978, G979, G980, G981, G982, G983, G984, G985, G986, G987,
         G988, G989, G990, G991, G992, G993, G994, G995, G996, G997, G998,
         G999, G1000, G1001, G1002, G1003, G1004, G1005, G1006, G1007, G1008,
         G1009, G1010, G1011, G1012, G1013, G1014, G1015, G1016, G1017, G1018,
         G1019, G1020, G1021, G1022, G1023, G1024, G1025, G1026, G1027, G1028,
         G1029, G1030, G1031, G1032, G1033, G1034, G1035, G1036, G1037, G1038,
         G1039, G1040, G1041, G1042, G1043, G1044, G1045, G1046, G1047, G1048,
         G1049, G1050, G1051, G1052, G1053, G1054, G1055, G1056, G1057, G1058,
         G1059, G1060, G1061, G1062, G1063, G1064, G1065, G1066, G1067, G1068,
         G1069, G1070, G1071, G1072, G1073, G1074, G1075, G1076, G1077, G1078,
         G1079, G1080, G1081, G1082, G1083, G1084, G1085, G1086, G1087, G1088,
         G1089, G1090, G1091, G1092, G1093, G1094, G1095, G1096, G1097, G1098,
         G1099, G1100, G1101, G1102, G1103, G1104, G1105, G1106, G1107, G1108,
         G1109, G1110, G1111, G1112, G1113, G1114, G1115, G1116, G1117, G1118,
         G1119, G1120, G1121, G1122, G1123, G1124, G1125, G1126, G1127, G1128,
         G1129, G1130, G1131, G1132, G1133, G1134, G1135, G1136, G1137, G1138,
         G1139, G1140, G1141, G1142, G1143, G1144, G1145, G1146, G1147, G1148,
         G1149, G1150, G1151, G1152, G1153, G1154, G1155, G1156, G1157, G1158,
         G1159, G1160, G1161, G1162, G1163, G1164, G1165, G1166, G1167, G1168,
         G1169, G1170, G1171, G1172, G1173, G1174, G1175, G1176, G1177, G1178,
         G1179, G1180, G1181, G1182, G1183, G1747, G1184, G1185, G1186, G1748,
         G1187, G1749, G1188, G1189, G1750, G1751;
  inout G21356,  G21357,  G21358,  G21359,  G21360,  G21361,  G21362,  G21363, 
     G21364,  G21365,  G21366,  G21367,  G21368,  G21369,  G21370,  G21371, 
     G21372,  G21373,  G21374,  G21375,  G21376,  G21377,  G21378,  G21379, 
     G21380,  G21381,  G21382,  G21383,  G21384,  G21385,  G21386,  G21387, 
     G21388,  G21389,  G21662,  G21663,  G21664,  G21665,  G21666,  G21667, 
     G21668,  G21669,  G21670,  G21671,  G21672,  G21673,  G21674,  G21675, 
     G21676,  G21677,  G21678,  G21679,  G21680,  G21681,  G21682,  G21683, 
     G21684,  G21685,  G21686,  G21687,  G21688,  G21689,  G21690,  G21691, 
     G21692,  G21693,  G21794,  G21799,  G21800,  G21802;
  wire   n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529;

  NOR2X2 U7327 ( .A(n10015), .B(G21428), .Y(n10020) );
  AND2X2 U7328 ( .A(n7564), .B(n6891), .Y(n6882) );
  INVX3 U7329 ( .A(n6889), .Y(n6903) );
  NOR2X2 U7330 ( .A(n9651), .B(n9751), .Y(n9655) );
  NOR2X2 U7331 ( .A(n7444), .B(n10120), .Y(n10121) );
  NOR2X2 U7332 ( .A(n9651), .B(n8743), .Y(n9650) );
  NOR2X4 U7333 ( .A(n8804), .B(n8784), .Y(n7569) );
  INVX3 U7334 ( .A(n7564), .Y(n9085) );
  NOR2X4 U7335 ( .A(n9093), .B(G21797), .Y(n7564) );
  NAND3X2 U7336 ( .A(n9623), .B(n7430), .C(G21428), .Y(n9319) );
  NAND2X2 U7337 ( .A(n8818), .B(n9752), .Y(n9651) );
  NAND2X2 U7338 ( .A(n9269), .B(n12912), .Y(n6891) );
  NAND2X2 U7339 ( .A(n9637), .B(n9638), .Y(n9325) );
  AND2X2 U7340 ( .A(n10198), .B(n9644), .Y(n10120) );
  NOR2X2 U7341 ( .A(n8932), .B(G21390), .Y(n8946) );
  NOR2X2 U7342 ( .A(n9759), .B(n9192), .Y(n9772) );
  NOR2X2 U7343 ( .A(n8932), .B(n8955), .Y(n8928) );
  NOR2X2 U7344 ( .A(n7428), .B(n8817), .Y(n9755) );
  NOR2XL U7345 ( .A(n6901), .B(n7198), .Y(n11326) );
  NAND2X2 U7346 ( .A(n9625), .B(n9626), .Y(n9321) );
  INVX3 U7347 ( .A(n6887), .Y(n6905) );
  NAND2XL U7348 ( .A(n6891), .B(n10225), .Y(n6887) );
  INVX3 U7349 ( .A(n9926), .Y(n9908) );
  NOR2X4 U7350 ( .A(n12706), .B(n12707), .Y(n9926) );
  INVX3 U7351 ( .A(n7300), .Y(n7020) );
  AND2X2 U7352 ( .A(n10112), .B(n10113), .Y(n10015) );
  INVX2 U7353 ( .A(n8711), .Y(n9076) );
  NAND4X2 U7354 ( .A(n13509), .B(n13510), .C(n13511), .D(n13512), .Y(n8711) );
  NAND2X2 U7355 ( .A(n8818), .B(n10008), .Y(n9759) );
  NAND4XL U7356 ( .A(n10009), .B(n10010), .C(n10011), .D(n10012), .Y(n10008)
         );
  INVX3 U7357 ( .A(n9623), .Y(n9324) );
  NOR4XL U7358 ( .A(n9441), .B(n9558), .C(n9559), .D(n9560), .Y(n9557) );
  NOR4XL U7359 ( .A(n9441), .B(n9549), .C(n9550), .D(n9551), .Y(n9548) );
  NOR4XL U7360 ( .A(n9441), .B(n9541), .C(n9542), .D(n9543), .Y(n9540) );
  NAND2X2 U7361 ( .A(n7411), .B(n7420), .Y(n7011) );
  INVX3 U7362 ( .A(n8947), .Y(n8932) );
  INVXL U7363 ( .A(n10256), .Y(n9192) );
  NAND2XL U7364 ( .A(n11339), .B(n10256), .Y(n11405) );
  NAND2XL U7365 ( .A(n11492), .B(n10256), .Y(n11487) );
  NAND2XL U7366 ( .A(n11575), .B(n10256), .Y(n11570) );
  NAND2XL U7367 ( .A(n11706), .B(n10256), .Y(n11700) );
  NAND2XL U7368 ( .A(n12697), .B(n10256), .Y(n12692) );
  NAND3XL U7369 ( .A(n10254), .B(n10255), .C(n10256), .Y(n10249) );
  NAND3XL U7370 ( .A(n10359), .B(n10360), .C(n10256), .Y(n10353) );
  NAND3XL U7371 ( .A(n12680), .B(n12681), .C(n10256), .Y(n12675) );
  NAND2XL U7372 ( .A(n10256), .B(n10527), .Y(n10528) );
  NAND2XL U7373 ( .A(n10256), .B(n10529), .Y(n10695) );
  NAND2XL U7374 ( .A(n10256), .B(n9406), .Y(n10778) );
  NAND2XL U7375 ( .A(n10256), .B(n10696), .Y(n11003) );
  NAND2XL U7376 ( .A(n10256), .B(n9436), .Y(n11068) );
  NAND2XL U7377 ( .A(n10256), .B(n11004), .Y(n11205) );
  INVX3 U7378 ( .A(n9260), .Y(n10227) );
  NOR2X2 U7379 ( .A(n7429), .B(n8817), .Y(n9260) );
  NAND4X1 U7380 ( .A(n6878), .B(n6879), .C(n6880), .D(n6881), .Y(G999) );
  NAND2X1 U7381 ( .A(n6882), .B(n6883), .Y(n6881) );
  NOR2X1 U7382 ( .A(n6884), .B(n6885), .Y(n6880) );
  NOR2X1 U7383 ( .A(n6886), .B(n6887), .Y(n6885) );
  NOR2X1 U7384 ( .A(n6888), .B(n6889), .Y(n6884) );
  NAND2X1 U7385 ( .A(n6890), .B(G21768), .Y(n6879) );
  OR2X1 U7386 ( .A(n6891), .B(n6892), .Y(n6878) );
  NAND4X1 U7387 ( .A(n6893), .B(n6894), .C(n6895), .D(n6896), .Y(G998) );
  NOR2X1 U7388 ( .A(n6897), .B(n6898), .Y(n6896) );
  NOR2X1 U7389 ( .A(n6899), .B(n6891), .Y(n6898) );
  NOR2X1 U7390 ( .A(n6900), .B(n6901), .Y(n6897) );
  NAND2X1 U7391 ( .A(n6882), .B(n6902), .Y(n6895) );
  NAND2X1 U7392 ( .A(n6903), .B(n6904), .Y(n6894) );
  NAND2X1 U7393 ( .A(n6905), .B(n6906), .Y(n6893) );
  NAND4X1 U7394 ( .A(n6907), .B(n6908), .C(n6909), .D(n6910), .Y(G997) );
  NOR2X1 U7395 ( .A(n6911), .B(n6912), .Y(n6910) );
  NOR2X1 U7396 ( .A(n6913), .B(n6891), .Y(n6912) );
  NOR2X1 U7397 ( .A(n6914), .B(n6901), .Y(n6911) );
  NAND2X1 U7398 ( .A(n6882), .B(n6915), .Y(n6909) );
  NAND2X1 U7399 ( .A(n6903), .B(n6916), .Y(n6908) );
  NAND2X1 U7400 ( .A(n6905), .B(n6917), .Y(n6907) );
  NAND4X1 U7401 ( .A(n6918), .B(n6919), .C(n6920), .D(n6921), .Y(G996) );
  NOR2X1 U7402 ( .A(n6922), .B(n6923), .Y(n6921) );
  NOR2X1 U7403 ( .A(n6924), .B(n6891), .Y(n6923) );
  NOR2X1 U7404 ( .A(n6925), .B(n6901), .Y(n6922) );
  NAND2X1 U7405 ( .A(n6882), .B(n6926), .Y(n6920) );
  NAND2X1 U7406 ( .A(n6927), .B(n6903), .Y(n6919) );
  NAND2X1 U7407 ( .A(n6905), .B(n6928), .Y(n6918) );
  NAND4X1 U7408 ( .A(n6929), .B(n6930), .C(n6931), .D(n6932), .Y(G995) );
  NOR2X1 U7409 ( .A(n6933), .B(n6934), .Y(n6932) );
  NOR2X1 U7410 ( .A(n6935), .B(n6891), .Y(n6934) );
  NOR2X1 U7411 ( .A(n6936), .B(n6901), .Y(n6933) );
  NAND2X1 U7412 ( .A(n6882), .B(n6937), .Y(n6931) );
  NAND2X1 U7413 ( .A(n6938), .B(n6903), .Y(n6930) );
  NAND2X1 U7414 ( .A(n6905), .B(n6939), .Y(n6929) );
  NAND4X1 U7415 ( .A(n6940), .B(n6941), .C(n6942), .D(n6943), .Y(G994) );
  NOR2X1 U7416 ( .A(n6944), .B(n6945), .Y(n6943) );
  NOR2X1 U7417 ( .A(n6946), .B(n6891), .Y(n6945) );
  NOR2X1 U7418 ( .A(n6947), .B(n6901), .Y(n6944) );
  NAND2X1 U7419 ( .A(n6882), .B(n6948), .Y(n6942) );
  NAND2X1 U7420 ( .A(n6949), .B(n6903), .Y(n6941) );
  NAND2X1 U7421 ( .A(n6905), .B(n6950), .Y(n6940) );
  NAND4X1 U7422 ( .A(n6951), .B(n6952), .C(n6953), .D(n6954), .Y(G993) );
  NOR2X1 U7423 ( .A(n6955), .B(n6956), .Y(n6954) );
  NOR2X1 U7424 ( .A(n6957), .B(n6891), .Y(n6956) );
  NOR2X1 U7425 ( .A(n6958), .B(n6901), .Y(n6955) );
  NAND2X1 U7426 ( .A(n6882), .B(n6959), .Y(n6953) );
  NAND2X1 U7427 ( .A(n6960), .B(n6903), .Y(n6952) );
  NAND2X1 U7428 ( .A(n6905), .B(n6961), .Y(n6951) );
  NAND4X1 U7429 ( .A(n6962), .B(n6963), .C(n6964), .D(n6965), .Y(G992) );
  NOR2X1 U7430 ( .A(n6966), .B(n6967), .Y(n6965) );
  NOR2X1 U7431 ( .A(n6968), .B(n6891), .Y(n6967) );
  AND2X1 U7432 ( .A(G21761), .B(n6890), .Y(n6966) );
  NAND2X1 U7433 ( .A(n6882), .B(n6969), .Y(n6964) );
  NAND2X1 U7434 ( .A(n6970), .B(n6903), .Y(n6963) );
  NAND2X1 U7435 ( .A(n6905), .B(n6971), .Y(n6962) );
  NAND4X1 U7436 ( .A(n6972), .B(n6973), .C(n6974), .D(n6975), .Y(G991) );
  NOR2X1 U7437 ( .A(n6976), .B(n6977), .Y(n6975) );
  NOR2X1 U7438 ( .A(n6978), .B(n6891), .Y(n6977) );
  AND2X1 U7439 ( .A(G21760), .B(n6890), .Y(n6976) );
  NAND2X1 U7440 ( .A(n6882), .B(n6979), .Y(n6974) );
  NAND2X1 U7441 ( .A(n6980), .B(n6903), .Y(n6973) );
  NAND2X1 U7442 ( .A(n6905), .B(n6981), .Y(n6972) );
  NAND4X1 U7443 ( .A(n6982), .B(n6983), .C(n6984), .D(n6985), .Y(G990) );
  NOR2X1 U7444 ( .A(n6986), .B(n6987), .Y(n6985) );
  NOR2X1 U7445 ( .A(n6988), .B(n6891), .Y(n6987) );
  NOR2X1 U7446 ( .A(n6989), .B(n6901), .Y(n6986) );
  NAND2X1 U7447 ( .A(n6882), .B(n6990), .Y(n6984) );
  NAND2X1 U7448 ( .A(n6991), .B(n6903), .Y(n6983) );
  NAND2X1 U7449 ( .A(n6905), .B(n6992), .Y(n6982) );
  NAND4X1 U7450 ( .A(n6993), .B(n6994), .C(n6995), .D(n6996), .Y(G989) );
  NOR2X1 U7451 ( .A(n6997), .B(n6998), .Y(n6996) );
  NOR2X1 U7452 ( .A(n6999), .B(n6891), .Y(n6998) );
  NOR2X1 U7453 ( .A(n7000), .B(n6901), .Y(n6997) );
  NAND2X1 U7454 ( .A(n6882), .B(n7001), .Y(n6995) );
  NAND2X1 U7455 ( .A(n6903), .B(n7002), .Y(n6994) );
  NAND2X1 U7456 ( .A(n6905), .B(n7003), .Y(n6993) );
  NAND4X1 U7457 ( .A(n7004), .B(n7005), .C(n7006), .D(n7007), .Y(G988) );
  NOR3X1 U7458 ( .A(n7008), .B(n7009), .C(n7010), .Y(n7007) );
  NOR3X1 U7459 ( .A(G21598), .B(n7011), .C(n7012), .Y(n7010) );
  NOR2X1 U7460 ( .A(n7013), .B(n7014), .Y(n7009) );
  NOR2X1 U7461 ( .A(n7015), .B(n7016), .Y(n7013) );
  NOR2X1 U7462 ( .A(n7017), .B(n7011), .Y(n7015) );
  NOR2X1 U7463 ( .A(n7018), .B(n7019), .Y(n7008) );
  NAND2X1 U7464 ( .A(n7020), .B(n7021), .Y(n7006) );
  NAND2X1 U7465 ( .A(n7022), .B(n7023), .Y(n7005) );
  NAND2X1 U7466 ( .A(n7024), .B(n7025), .Y(n7004) );
  NAND4X1 U7467 ( .A(n7026), .B(n7027), .C(n7028), .D(n7029), .Y(G987) );
  NOR3X1 U7468 ( .A(n7030), .B(n7031), .C(n7032), .Y(n7029) );
  NOR2X1 U7469 ( .A(n7033), .B(n7019), .Y(n7032) );
  NOR2X1 U7470 ( .A(n7034), .B(n7011), .Y(n7031) );
  NOR2X1 U7471 ( .A(n7035), .B(n7036), .Y(n7030) );
  NAND2X1 U7472 ( .A(n7020), .B(n7037), .Y(n7028) );
  NAND2X1 U7473 ( .A(n7038), .B(n7022), .Y(n7027) );
  NAND2X1 U7474 ( .A(n7024), .B(n7039), .Y(n7026) );
  NAND4X1 U7475 ( .A(n7040), .B(n7041), .C(n7042), .D(n7043), .Y(G986) );
  NOR3X1 U7476 ( .A(n7044), .B(n7045), .C(n7046), .Y(n7043) );
  NOR2X1 U7477 ( .A(n7047), .B(n7048), .Y(n7046) );
  NOR3X1 U7478 ( .A(n7011), .B(n7049), .C(n7050), .Y(n7045) );
  NOR2X1 U7479 ( .A(n7051), .B(n7052), .Y(n7044) );
  NAND2X1 U7480 ( .A(n7016), .B(G21596), .Y(n7042) );
  NAND2X1 U7481 ( .A(n7020), .B(n7053), .Y(n7041) );
  NAND2X1 U7482 ( .A(n7054), .B(G21787), .Y(n7040) );
  NAND4X1 U7483 ( .A(n7055), .B(n7056), .C(n7057), .D(n7058), .Y(G985) );
  NOR3X1 U7484 ( .A(n7059), .B(n7060), .C(n7061), .Y(n7058) );
  NOR2X1 U7485 ( .A(n7062), .B(n7019), .Y(n7061) );
  NOR2X1 U7486 ( .A(n7063), .B(n7011), .Y(n7060) );
  NOR2X1 U7487 ( .A(n7064), .B(n7036), .Y(n7059) );
  NAND2X1 U7488 ( .A(n7020), .B(n7065), .Y(n7057) );
  NAND2X1 U7489 ( .A(n7066), .B(n7022), .Y(n7056) );
  NAND2X1 U7490 ( .A(n7024), .B(n7067), .Y(n7055) );
  NAND4X1 U7491 ( .A(n7068), .B(n7069), .C(n7070), .D(n7071), .Y(G984) );
  NOR3X1 U7492 ( .A(n7072), .B(n7073), .C(n7074), .Y(n7071) );
  NOR2X1 U7493 ( .A(n7047), .B(n7075), .Y(n7074) );
  NOR3X1 U7494 ( .A(n7011), .B(n7076), .C(n7077), .Y(n7073) );
  NOR2X1 U7495 ( .A(n7078), .B(n7052), .Y(n7072) );
  NAND2X1 U7496 ( .A(n7016), .B(G21594), .Y(n7070) );
  NAND2X1 U7497 ( .A(n7020), .B(n7079), .Y(n7069) );
  NAND2X1 U7498 ( .A(n7054), .B(G21785), .Y(n7068) );
  NAND4X1 U7499 ( .A(n7080), .B(n7081), .C(n7082), .D(n7083), .Y(G983) );
  NOR3X1 U7500 ( .A(n7084), .B(n7085), .C(n7086), .Y(n7083) );
  NOR2X1 U7501 ( .A(n7047), .B(n7087), .Y(n7086) );
  NOR3X1 U7502 ( .A(n7011), .B(n7088), .C(n7089), .Y(n7085) );
  NOR2X1 U7503 ( .A(n7090), .B(n7052), .Y(n7084) );
  NAND2X1 U7504 ( .A(n7016), .B(G21593), .Y(n7082) );
  NAND2X1 U7505 ( .A(n7020), .B(n7091), .Y(n7081) );
  NAND2X1 U7506 ( .A(n7054), .B(G21784), .Y(n7080) );
  NAND4X1 U7507 ( .A(n7092), .B(n7093), .C(n7094), .D(n7095), .Y(G982) );
  NOR3X1 U7508 ( .A(n7096), .B(n7097), .C(n7098), .Y(n7095) );
  NOR2X1 U7509 ( .A(n7099), .B(n7019), .Y(n7098) );
  NOR2X1 U7510 ( .A(n7100), .B(n7011), .Y(n7097) );
  NOR2X1 U7511 ( .A(n7101), .B(n7036), .Y(n7096) );
  NAND2X1 U7512 ( .A(n7020), .B(n7102), .Y(n7094) );
  NAND2X1 U7513 ( .A(n7103), .B(n7022), .Y(n7093) );
  NAND2X1 U7514 ( .A(n7024), .B(n7104), .Y(n7092) );
  NAND4X1 U7515 ( .A(n7105), .B(n7106), .C(n7107), .D(n7108), .Y(G981) );
  NOR3X1 U7516 ( .A(n7109), .B(n7110), .C(n7111), .Y(n7108) );
  NOR2X1 U7517 ( .A(n7047), .B(n7112), .Y(n7111) );
  NOR2X1 U7518 ( .A(n7113), .B(n7011), .Y(n7110) );
  NOR2X1 U7519 ( .A(n7114), .B(n7052), .Y(n7109) );
  NAND2X1 U7520 ( .A(n7016), .B(G21591), .Y(n7107) );
  NAND2X1 U7521 ( .A(n7020), .B(n7115), .Y(n7106) );
  NAND2X1 U7522 ( .A(n7054), .B(G21782), .Y(n7105) );
  NAND4X1 U7523 ( .A(n7116), .B(n7117), .C(n7118), .D(n7119), .Y(G980) );
  NOR3X1 U7524 ( .A(n7120), .B(n7121), .C(n7122), .Y(n7119) );
  NOR2X1 U7525 ( .A(n7123), .B(n7019), .Y(n7122) );
  NOR2X1 U7526 ( .A(n7124), .B(n7011), .Y(n7121) );
  AND2X1 U7527 ( .A(G21590), .B(n7016), .Y(n7120) );
  NAND2X1 U7528 ( .A(n7020), .B(n7125), .Y(n7118) );
  NAND2X1 U7529 ( .A(n7126), .B(n7022), .Y(n7117) );
  NAND2X1 U7530 ( .A(n7024), .B(n7127), .Y(n7116) );
  NAND4X1 U7531 ( .A(n7128), .B(n7129), .C(n7130), .D(n7131), .Y(G979) );
  NOR3X1 U7532 ( .A(n7132), .B(n7133), .C(n7134), .Y(n7131) );
  NOR2X1 U7533 ( .A(n7135), .B(n7019), .Y(n7134) );
  NOR2X1 U7534 ( .A(n7136), .B(n7011), .Y(n7133) );
  NOR2X1 U7535 ( .A(n7137), .B(n7036), .Y(n7132) );
  NAND2X1 U7536 ( .A(n7020), .B(n7138), .Y(n7130) );
  NAND2X1 U7537 ( .A(n7139), .B(n7022), .Y(n7129) );
  NAND2X1 U7538 ( .A(n7024), .B(n7140), .Y(n7128) );
  NAND4X1 U7539 ( .A(n7141), .B(n7142), .C(n7143), .D(n7144), .Y(G978) );
  NOR3X1 U7540 ( .A(n7145), .B(n7146), .C(n7147), .Y(n7144) );
  NOR2X1 U7541 ( .A(n7148), .B(n7019), .Y(n7147) );
  NOR2X1 U7542 ( .A(n7149), .B(n7011), .Y(n7146) );
  NOR2X1 U7543 ( .A(n7150), .B(n7036), .Y(n7145) );
  NAND2X1 U7544 ( .A(n7020), .B(n7151), .Y(n7143) );
  NAND2X1 U7545 ( .A(n7152), .B(n7022), .Y(n7142) );
  NAND2X1 U7546 ( .A(n7024), .B(n7153), .Y(n7141) );
  NAND4X1 U7547 ( .A(n7154), .B(n7155), .C(n7156), .D(n7157), .Y(G977) );
  NOR3X1 U7548 ( .A(n7158), .B(n7159), .C(n7160), .Y(n7157) );
  NOR2X1 U7549 ( .A(n7161), .B(n7019), .Y(n7160) );
  NOR2X1 U7550 ( .A(n7162), .B(n7011), .Y(n7159) );
  AND2X1 U7551 ( .A(G21587), .B(n7016), .Y(n7158) );
  NAND2X1 U7552 ( .A(n7020), .B(n7163), .Y(n7156) );
  NAND2X1 U7553 ( .A(n7164), .B(n7022), .Y(n7155) );
  NAND2X1 U7554 ( .A(n7024), .B(n7165), .Y(n7154) );
  NAND4X1 U7555 ( .A(n7166), .B(n7167), .C(n7168), .D(n7169), .Y(G976) );
  NOR3X1 U7556 ( .A(n7170), .B(n7171), .C(n7172), .Y(n7169) );
  NOR2X1 U7557 ( .A(n7173), .B(n7019), .Y(n7172) );
  NOR2X1 U7558 ( .A(n7174), .B(n7011), .Y(n7171) );
  NOR2X1 U7559 ( .A(n7175), .B(n7036), .Y(n7170) );
  NAND2X1 U7560 ( .A(n7020), .B(n7176), .Y(n7168) );
  NAND2X1 U7561 ( .A(n7177), .B(n7022), .Y(n7167) );
  NAND2X1 U7562 ( .A(n7024), .B(n7178), .Y(n7166) );
  NAND4X1 U7563 ( .A(n7179), .B(n7180), .C(n7181), .D(n7182), .Y(G975) );
  NOR3X1 U7564 ( .A(n7183), .B(n7184), .C(n7185), .Y(n7182) );
  NOR2X1 U7565 ( .A(n7186), .B(n7019), .Y(n7185) );
  NOR2X1 U7566 ( .A(n7187), .B(n7011), .Y(n7184) );
  AND2X1 U7567 ( .A(G21585), .B(n7016), .Y(n7183) );
  NAND2X1 U7568 ( .A(n7020), .B(n7188), .Y(n7181) );
  NAND2X1 U7569 ( .A(n7189), .B(n7022), .Y(n7180) );
  NAND2X1 U7570 ( .A(n7024), .B(n7190), .Y(n7179) );
  NAND4X1 U7571 ( .A(n7191), .B(n7192), .C(n7193), .D(n7194), .Y(G974) );
  NOR3X1 U7572 ( .A(n7195), .B(n7196), .C(n7197), .Y(n7194) );
  NOR2X1 U7573 ( .A(n7198), .B(n7019), .Y(n7197) );
  NOR2X1 U7574 ( .A(n7199), .B(n7011), .Y(n7196) );
  NOR2X1 U7575 ( .A(n7200), .B(n7036), .Y(n7195) );
  NAND2X1 U7576 ( .A(n7020), .B(n7201), .Y(n7193) );
  NAND2X1 U7577 ( .A(n7202), .B(n7022), .Y(n7192) );
  NAND2X1 U7578 ( .A(n7024), .B(n7203), .Y(n7191) );
  NAND4X1 U7579 ( .A(n7204), .B(n7205), .C(n7206), .D(n7207), .Y(G973) );
  NOR3X1 U7580 ( .A(n7208), .B(n7209), .C(n7210), .Y(n7207) );
  NOR2X1 U7581 ( .A(n7211), .B(n7019), .Y(n7210) );
  NOR2X1 U7582 ( .A(n7212), .B(n7011), .Y(n7209) );
  NOR2X1 U7583 ( .A(n7213), .B(n7036), .Y(n7208) );
  NAND2X1 U7584 ( .A(n7020), .B(n7214), .Y(n7206) );
  NAND2X1 U7585 ( .A(n7022), .B(n7215), .Y(n7205) );
  NAND2X1 U7586 ( .A(n7024), .B(n7216), .Y(n7204) );
  NAND4X1 U7587 ( .A(n7217), .B(n7218), .C(n7219), .D(n7220), .Y(G972) );
  NOR3X1 U7588 ( .A(n7221), .B(n7222), .C(n7223), .Y(n7220) );
  NOR4X1 U7589 ( .A(G21582), .B(n7011), .C(n7224), .D(n7225), .Y(n7223) );
  NOR2X1 U7590 ( .A(n7226), .B(n7227), .Y(n7222) );
  NOR2X1 U7591 ( .A(n7228), .B(n7229), .Y(n7226) );
  NOR2X1 U7592 ( .A(G21581), .B(n7011), .Y(n7228) );
  NOR2X1 U7593 ( .A(n7230), .B(n7019), .Y(n7221) );
  NAND2X1 U7594 ( .A(n7020), .B(n7231), .Y(n7219) );
  NAND2X1 U7595 ( .A(n7232), .B(n7022), .Y(n7218) );
  NAND2X1 U7596 ( .A(n7024), .B(n7233), .Y(n7217) );
  NAND4X1 U7597 ( .A(n7234), .B(n7235), .C(n7236), .D(n7237), .Y(G971) );
  NOR3X1 U7598 ( .A(n7238), .B(n7239), .C(n7240), .Y(n7237) );
  NOR3X1 U7599 ( .A(G21581), .B(n7225), .C(n7011), .Y(n7240) );
  AND2X1 U7600 ( .A(n7229), .B(G21581), .Y(n7239) );
  NAND2X1 U7601 ( .A(n7036), .B(n7241), .Y(n7229) );
  NAND2X1 U7602 ( .A(n7242), .B(n7225), .Y(n7241) );
  NOR2X1 U7603 ( .A(n7243), .B(n7019), .Y(n7238) );
  NAND2X1 U7604 ( .A(n7020), .B(n7244), .Y(n7236) );
  NAND2X1 U7605 ( .A(n7245), .B(n7022), .Y(n7235) );
  NAND2X1 U7606 ( .A(n7024), .B(n7246), .Y(n7234) );
  NAND4X1 U7607 ( .A(n7247), .B(n7248), .C(n7249), .D(n7250), .Y(G970) );
  NOR3X1 U7608 ( .A(n7251), .B(n7252), .C(n7253), .Y(n7250) );
  NOR4X1 U7609 ( .A(G21580), .B(n7011), .C(n7254), .D(n7255), .Y(n7253) );
  NOR2X1 U7610 ( .A(n7256), .B(n7257), .Y(n7252) );
  NOR2X1 U7611 ( .A(n7258), .B(n7259), .Y(n7256) );
  NOR2X1 U7612 ( .A(G21579), .B(n7011), .Y(n7258) );
  NOR2X1 U7613 ( .A(n7260), .B(n7019), .Y(n7251) );
  NAND2X1 U7614 ( .A(n7020), .B(n7261), .Y(n7249) );
  NAND2X1 U7615 ( .A(n7262), .B(n7022), .Y(n7248) );
  NAND2X1 U7616 ( .A(n7024), .B(n7263), .Y(n7247) );
  NAND4X1 U7617 ( .A(n7264), .B(n7265), .C(n7266), .D(n7267), .Y(G969) );
  NOR3X1 U7618 ( .A(n7268), .B(n7269), .C(n7270), .Y(n7267) );
  NOR3X1 U7619 ( .A(G21579), .B(n7255), .C(n7011), .Y(n7270) );
  AND2X1 U7620 ( .A(n7259), .B(G21579), .Y(n7269) );
  NAND2X1 U7621 ( .A(n7036), .B(n7271), .Y(n7259) );
  NAND2X1 U7622 ( .A(n7242), .B(n7255), .Y(n7271) );
  NOR2X1 U7623 ( .A(n7272), .B(n7019), .Y(n7268) );
  NAND2X1 U7624 ( .A(n7020), .B(n7273), .Y(n7266) );
  NAND2X1 U7625 ( .A(n7274), .B(n7022), .Y(n7265) );
  NAND2X1 U7626 ( .A(n7024), .B(n7275), .Y(n7264) );
  NAND4X1 U7627 ( .A(n7276), .B(n7277), .C(n7278), .D(n7279), .Y(G968) );
  NOR3X1 U7628 ( .A(n7280), .B(n7281), .C(n7282), .Y(n7279) );
  NOR4X1 U7629 ( .A(G21578), .B(n7011), .C(n7283), .D(n7284), .Y(n7282) );
  NOR2X1 U7630 ( .A(n7285), .B(n7286), .Y(n7281) );
  INVX1 U7631 ( .A(G21578), .Y(n7286) );
  NOR2X1 U7632 ( .A(n7287), .B(n7288), .Y(n7285) );
  NOR2X1 U7633 ( .A(G21577), .B(n7011), .Y(n7287) );
  AND2X1 U7634 ( .A(G21769), .B(n7054), .Y(n7280) );
  NAND2X1 U7635 ( .A(n7289), .B(n7020), .Y(n7278) );
  NAND2X1 U7636 ( .A(n7290), .B(n7022), .Y(n7277) );
  NAND2X1 U7637 ( .A(n7024), .B(n7291), .Y(n7276) );
  NAND4X1 U7638 ( .A(n7292), .B(n7293), .C(n7294), .D(n7295), .Y(G967) );
  NOR3X1 U7639 ( .A(n7296), .B(n7297), .C(n7298), .Y(n7295) );
  NOR2X1 U7640 ( .A(n7299), .B(n7052), .Y(n7298) );
  NOR2X1 U7641 ( .A(n6886), .B(n7047), .Y(n7297) );
  NOR2X1 U7642 ( .A(n6888), .B(n7300), .Y(n7296) );
  NAND2X1 U7643 ( .A(n7054), .B(G21768), .Y(n7294) );
  NAND2X1 U7644 ( .A(G21577), .B(n7288), .Y(n7293) );
  NAND2X1 U7645 ( .A(n7036), .B(n7301), .Y(n7288) );
  NAND2X1 U7646 ( .A(n7242), .B(n7284), .Y(n7301) );
  INVX1 U7647 ( .A(n7302), .Y(n7284) );
  NAND3X1 U7648 ( .A(n7242), .B(n7302), .C(n7283), .Y(n7292) );
  INVX1 U7649 ( .A(G21577), .Y(n7283) );
  NAND4X1 U7650 ( .A(n7303), .B(n7304), .C(n7305), .D(n7306), .Y(G966) );
  NOR3X1 U7651 ( .A(n7307), .B(n7308), .C(n7309), .Y(n7306) );
  NOR2X1 U7652 ( .A(n7310), .B(n7047), .Y(n7309) );
  AND2X1 U7653 ( .A(n7311), .B(n7242), .Y(n7308) );
  ADDHXL U7654 ( .A(n7312), .B(n7313), .S(n7311) );
  NOR2X1 U7655 ( .A(n7314), .B(n7052), .Y(n7307) );
  NAND2X1 U7656 ( .A(n7016), .B(G21576), .Y(n7305) );
  NAND2X1 U7657 ( .A(n7020), .B(n6904), .Y(n7304) );
  NAND2X1 U7658 ( .A(n7054), .B(G21767), .Y(n7303) );
  NAND4X1 U7659 ( .A(n7315), .B(n7316), .C(n7317), .D(n7318), .Y(G965) );
  NOR3X1 U7660 ( .A(n7319), .B(n7320), .C(n7321), .Y(n7318) );
  AND3X1 U7661 ( .A(n7322), .B(n7323), .C(n7242), .Y(n7321) );
  NOR2X1 U7662 ( .A(n7324), .B(n7322), .Y(n7320) );
  INVX1 U7663 ( .A(G21575), .Y(n7322) );
  NOR2X1 U7664 ( .A(n7325), .B(n7016), .Y(n7324) );
  NOR2X1 U7665 ( .A(n7323), .B(n7011), .Y(n7325) );
  NOR2X1 U7666 ( .A(n6914), .B(n7019), .Y(n7319) );
  INVX1 U7667 ( .A(G21766), .Y(n6914) );
  NAND2X1 U7668 ( .A(n7020), .B(n6916), .Y(n7317) );
  NAND2X1 U7669 ( .A(n7022), .B(n6917), .Y(n7316) );
  NAND2X1 U7670 ( .A(n7024), .B(n6915), .Y(n7315) );
  NAND4X1 U7671 ( .A(n7326), .B(n7327), .C(n7328), .D(n7329), .Y(G964) );
  NOR3X1 U7672 ( .A(n7330), .B(n7331), .C(n7332), .Y(n7329) );
  NOR4X1 U7673 ( .A(G21574), .B(n7011), .C(n7333), .D(n7334), .Y(n7332) );
  NOR2X1 U7674 ( .A(n7335), .B(n7336), .Y(n7331) );
  NOR2X1 U7675 ( .A(n7337), .B(n7338), .Y(n7335) );
  NOR2X1 U7676 ( .A(G21573), .B(n7011), .Y(n7337) );
  NOR2X1 U7677 ( .A(n6925), .B(n7019), .Y(n7330) );
  INVX1 U7678 ( .A(G21765), .Y(n6925) );
  NAND2X1 U7679 ( .A(n7020), .B(n6927), .Y(n7328) );
  NAND2X1 U7680 ( .A(n7022), .B(n6928), .Y(n7327) );
  NAND2X1 U7681 ( .A(n7024), .B(n6926), .Y(n7326) );
  NAND4X1 U7682 ( .A(n7339), .B(n7340), .C(n7341), .D(n7342), .Y(G963) );
  NOR3X1 U7683 ( .A(n7343), .B(n7344), .C(n7345), .Y(n7342) );
  NOR3X1 U7684 ( .A(G21573), .B(n7334), .C(n7011), .Y(n7345) );
  AND2X1 U7685 ( .A(n7338), .B(G21573), .Y(n7344) );
  NAND2X1 U7686 ( .A(n7036), .B(n7346), .Y(n7338) );
  NAND2X1 U7687 ( .A(n7242), .B(n7334), .Y(n7346) );
  NOR2X1 U7688 ( .A(n6936), .B(n7019), .Y(n7343) );
  INVX1 U7689 ( .A(G21764), .Y(n6936) );
  NAND2X1 U7690 ( .A(n7020), .B(n6938), .Y(n7341) );
  NAND2X1 U7691 ( .A(n7022), .B(n6939), .Y(n7340) );
  NAND2X1 U7692 ( .A(n7024), .B(n6937), .Y(n7339) );
  NAND4X1 U7693 ( .A(n7347), .B(n7348), .C(n7349), .D(n7350), .Y(G962) );
  NOR3X1 U7694 ( .A(n7351), .B(n7352), .C(n7353), .Y(n7350) );
  NOR4X1 U7695 ( .A(G21572), .B(n7011), .C(n7354), .D(n7355), .Y(n7353) );
  NOR2X1 U7696 ( .A(n7356), .B(n7357), .Y(n7352) );
  INVX1 U7697 ( .A(G21572), .Y(n7357) );
  NOR2X1 U7698 ( .A(n7358), .B(n7359), .Y(n7356) );
  NOR2X1 U7699 ( .A(G21571), .B(n7011), .Y(n7358) );
  NOR2X1 U7700 ( .A(n6947), .B(n7019), .Y(n7351) );
  INVX1 U7701 ( .A(G21763), .Y(n6947) );
  NAND2X1 U7702 ( .A(n7020), .B(n6949), .Y(n7349) );
  NAND2X1 U7703 ( .A(n7022), .B(n6950), .Y(n7348) );
  NAND2X1 U7704 ( .A(n7024), .B(n6948), .Y(n7347) );
  NAND4X1 U7705 ( .A(n7360), .B(n7361), .C(n7362), .D(n7363), .Y(G961) );
  NOR3X1 U7706 ( .A(n7364), .B(n7365), .C(n7366), .Y(n7363) );
  NOR3X1 U7707 ( .A(G21571), .B(n7355), .C(n7011), .Y(n7366) );
  NOR2X1 U7708 ( .A(n7367), .B(n7354), .Y(n7365) );
  INVX1 U7709 ( .A(G21571), .Y(n7354) );
  NOR2X1 U7710 ( .A(n6958), .B(n7019), .Y(n7364) );
  NAND2X1 U7711 ( .A(n7020), .B(n6960), .Y(n7362) );
  NAND2X1 U7712 ( .A(n7022), .B(n6961), .Y(n7361) );
  NAND2X1 U7713 ( .A(n7024), .B(n6959), .Y(n7360) );
  NAND4X1 U7714 ( .A(n7368), .B(n7369), .C(n7370), .D(n7371), .Y(G960) );
  NOR3X1 U7715 ( .A(n7372), .B(n7373), .C(n7374), .Y(n7371) );
  NOR2X1 U7716 ( .A(n7367), .B(n7375), .Y(n7374) );
  INVX1 U7717 ( .A(n7359), .Y(n7367) );
  NAND2X1 U7718 ( .A(n7036), .B(n7376), .Y(n7359) );
  NAND2X1 U7719 ( .A(n7242), .B(n7355), .Y(n7376) );
  INVX1 U7720 ( .A(n7377), .Y(n7355) );
  NOR3X1 U7721 ( .A(n7011), .B(n7377), .C(n7378), .Y(n7373) );
  NOR2X1 U7722 ( .A(n7379), .B(n7047), .Y(n7372) );
  NAND2X1 U7723 ( .A(n7054), .B(G21761), .Y(n7370) );
  NAND2X1 U7724 ( .A(n7024), .B(n6969), .Y(n7369) );
  NAND2X1 U7725 ( .A(n7020), .B(n6970), .Y(n7368) );
  NAND4X1 U7726 ( .A(n7380), .B(n7381), .C(n7382), .D(n7383), .Y(G959) );
  NOR3X1 U7727 ( .A(n7384), .B(n7385), .C(n7386), .Y(n7383) );
  NOR2X1 U7728 ( .A(n7387), .B(n7047), .Y(n7386) );
  NOR2X1 U7729 ( .A(n7388), .B(n7011), .Y(n7385) );
  NOR2X1 U7730 ( .A(n7389), .B(n7378), .Y(n7388) );
  NOR2X1 U7731 ( .A(n7390), .B(n7391), .Y(n7389) );
  NOR2X1 U7732 ( .A(n7392), .B(n7052), .Y(n7384) );
  NAND2X1 U7733 ( .A(n7016), .B(G21569), .Y(n7382) );
  NAND2X1 U7734 ( .A(n7020), .B(n6980), .Y(n7381) );
  NAND2X1 U7735 ( .A(n7054), .B(G21760), .Y(n7380) );
  NAND4X1 U7736 ( .A(n7393), .B(n7394), .C(n7395), .D(n7396), .Y(G958) );
  NOR3X1 U7737 ( .A(n7397), .B(n7398), .C(n7399), .Y(n7396) );
  AND3X1 U7738 ( .A(n7400), .B(n7401), .C(n7242), .Y(n7399) );
  INVX1 U7739 ( .A(n7011), .Y(n7242) );
  NOR2X1 U7740 ( .A(n7402), .B(n7400), .Y(n7398) );
  INVX1 U7741 ( .A(G21568), .Y(n7400) );
  NOR2X1 U7742 ( .A(n7403), .B(n7016), .Y(n7402) );
  NOR2X1 U7743 ( .A(n6989), .B(n7019), .Y(n7397) );
  INVX1 U7744 ( .A(n7054), .Y(n7019) );
  NAND2X1 U7745 ( .A(n7020), .B(n6991), .Y(n7395) );
  NAND2X1 U7746 ( .A(n7022), .B(n6992), .Y(n7394) );
  INVX1 U7747 ( .A(n7047), .Y(n7022) );
  NAND2X1 U7748 ( .A(n7024), .B(n6990), .Y(n7393) );
  INVX1 U7749 ( .A(n7052), .Y(n7024) );
  NAND4X1 U7750 ( .A(n7404), .B(n7405), .C(n7406), .D(n7407), .Y(G957) );
  NOR3X1 U7751 ( .A(n7408), .B(n7403), .C(n7409), .Y(n7407) );
  NOR2X1 U7752 ( .A(n7410), .B(n7047), .Y(n7409) );
  NAND2X1 U7753 ( .A(n7411), .B(n7412), .Y(n7047) );
  NAND4X1 U7754 ( .A(n7413), .B(n7414), .C(n7415), .D(n7416), .Y(n7412) );
  INVX1 U7755 ( .A(n7417), .Y(n7416) );
  NOR2X1 U7756 ( .A(n7418), .B(n7419), .Y(n7415) );
  NOR2X1 U7757 ( .A(n7401), .B(n7011), .Y(n7403) );
  NOR2X1 U7758 ( .A(n7421), .B(n7052), .Y(n7408) );
  NAND2X1 U7759 ( .A(n7411), .B(n7422), .Y(n7052) );
  NAND2X1 U7760 ( .A(n7423), .B(n7424), .Y(n7422) );
  NAND2X1 U7761 ( .A(n7016), .B(G21567), .Y(n7406) );
  NAND2X1 U7762 ( .A(n7020), .B(n7002), .Y(n7405) );
  NAND2X1 U7763 ( .A(n7411), .B(n7425), .Y(n7300) );
  NAND4X1 U7764 ( .A(n7426), .B(n7427), .C(n7428), .D(n7429), .Y(n7425) );
  NOR2X1 U7765 ( .A(n7430), .B(n7016), .Y(n7411) );
  NAND2X1 U7766 ( .A(n7054), .B(G21758), .Y(n7404) );
  NOR2X1 U7767 ( .A(G21426), .B(n7016), .Y(n7054) );
  INVX1 U7768 ( .A(n7036), .Y(n7016) );
  NAND2X1 U7769 ( .A(n7431), .B(n7432), .Y(n7036) );
  NAND2X1 U7770 ( .A(n7433), .B(n7434), .Y(n7432) );
  NAND4X1 U7771 ( .A(n7435), .B(n7436), .C(n7437), .D(n7438), .Y(n7434) );
  NAND3X1 U7772 ( .A(n7439), .B(n7440), .C(n7441), .Y(n7438) );
  NAND2X1 U7773 ( .A(n7442), .B(n7443), .Y(n7440) );
  NAND3X1 U7774 ( .A(n7444), .B(n7445), .C(n7446), .Y(n7443) );
  NAND2X1 U7775 ( .A(n7447), .B(n7448), .Y(n7437) );
  NAND2X1 U7776 ( .A(n7449), .B(n7450), .Y(n7448) );
  NAND2X1 U7777 ( .A(n7451), .B(n7452), .Y(n7450) );
  NAND2X1 U7778 ( .A(n7439), .B(n7453), .Y(n7452) );
  NAND2X1 U7779 ( .A(n7454), .B(n7455), .Y(n7453) );
  NAND2X1 U7780 ( .A(n7454), .B(n7456), .Y(n7449) );
  NAND2X1 U7781 ( .A(n7457), .B(n7458), .Y(n7436) );
  NAND3X1 U7782 ( .A(n7459), .B(n7460), .C(n7461), .Y(G956) );
  NAND2X1 U7783 ( .A(n7462), .B(G21565), .Y(n7461) );
  NAND2X1 U7784 ( .A(n7463), .B(n7464), .Y(n7460) );
  NAND2X1 U7785 ( .A(n7465), .B(n6990), .Y(n7459) );
  NAND3X1 U7786 ( .A(n7466), .B(n7467), .C(n7468), .Y(G955) );
  NAND2X1 U7787 ( .A(n7462), .B(G21564), .Y(n7468) );
  NAND2X1 U7788 ( .A(n7469), .B(n7463), .Y(n7467) );
  NAND2X1 U7789 ( .A(n7465), .B(n6979), .Y(n7466) );
  NAND3X1 U7790 ( .A(n7470), .B(n7471), .C(n7472), .Y(G954) );
  NAND2X1 U7791 ( .A(n7462), .B(G21563), .Y(n7472) );
  NAND3X1 U7792 ( .A(n7473), .B(n7430), .C(n7463), .Y(n7471) );
  NAND2X1 U7793 ( .A(n7465), .B(n6969), .Y(n7470) );
  NOR2X1 U7794 ( .A(n7474), .B(n7475), .Y(G953) );
  NAND4X1 U7795 ( .A(n7476), .B(n7477), .C(n7478), .D(n7479), .Y(G952) );
  NOR3X1 U7796 ( .A(n7480), .B(n7481), .C(n7482), .Y(n7479) );
  NOR2X1 U7797 ( .A(n7483), .B(n7484), .Y(n7482) );
  NOR2X1 U7798 ( .A(n7485), .B(n7486), .Y(n7481) );
  NOR2X1 U7799 ( .A(n7487), .B(n7488), .Y(n7480) );
  NAND2X1 U7800 ( .A(G32), .B(n7489), .Y(n7478) );
  NAND2X1 U7801 ( .A(G21556), .B(n7490), .Y(n7477) );
  NAND2X1 U7802 ( .A(G16), .B(n7491), .Y(n7476) );
  NAND4X1 U7803 ( .A(n7492), .B(n7493), .C(n7494), .D(n7495), .Y(G951) );
  NOR3X1 U7804 ( .A(n7496), .B(n7497), .C(n7498), .Y(n7495) );
  NOR2X1 U7805 ( .A(n7499), .B(n7484), .Y(n7498) );
  NOR2X1 U7806 ( .A(n7485), .B(n7500), .Y(n7497) );
  NOR2X1 U7807 ( .A(n7487), .B(n7501), .Y(n7496) );
  NAND2X1 U7808 ( .A(G31), .B(n7489), .Y(n7494) );
  NAND2X1 U7809 ( .A(G21555), .B(n7490), .Y(n7493) );
  NAND2X1 U7810 ( .A(G15), .B(n7491), .Y(n7492) );
  NAND4X1 U7811 ( .A(n7502), .B(n7503), .C(n7504), .D(n7505), .Y(G950) );
  NOR3X1 U7812 ( .A(n7506), .B(n7507), .C(n7508), .Y(n7505) );
  NOR2X1 U7813 ( .A(n7509), .B(n7484), .Y(n7508) );
  NOR2X1 U7814 ( .A(n7485), .B(n7510), .Y(n7507) );
  NOR2X1 U7815 ( .A(n7487), .B(n7511), .Y(n7506) );
  NAND2X1 U7816 ( .A(G30), .B(n7489), .Y(n7504) );
  NAND2X1 U7817 ( .A(G21554), .B(n7490), .Y(n7503) );
  NAND2X1 U7818 ( .A(G14), .B(n7491), .Y(n7502) );
  NAND4X1 U7819 ( .A(n7512), .B(n7513), .C(n7514), .D(n7515), .Y(G949) );
  NOR3X1 U7820 ( .A(n7516), .B(n7517), .C(n7518), .Y(n7515) );
  NOR2X1 U7821 ( .A(n7519), .B(n7484), .Y(n7518) );
  NOR2X1 U7822 ( .A(n7485), .B(n7520), .Y(n7517) );
  NOR2X1 U7823 ( .A(n7487), .B(n7521), .Y(n7516) );
  NAND2X1 U7824 ( .A(G29), .B(n7489), .Y(n7514) );
  NAND2X1 U7825 ( .A(G21553), .B(n7490), .Y(n7513) );
  NAND2X1 U7826 ( .A(G13), .B(n7491), .Y(n7512) );
  NAND4X1 U7827 ( .A(n7522), .B(n7523), .C(n7524), .D(n7525), .Y(G948) );
  NOR3X1 U7828 ( .A(n7526), .B(n7527), .C(n7528), .Y(n7525) );
  NOR2X1 U7829 ( .A(n7529), .B(n7484), .Y(n7528) );
  NOR2X1 U7830 ( .A(n7485), .B(n7530), .Y(n7527) );
  NOR2X1 U7831 ( .A(n7487), .B(n7531), .Y(n7526) );
  NAND2X1 U7832 ( .A(G28), .B(n7489), .Y(n7524) );
  NAND2X1 U7833 ( .A(G21552), .B(n7490), .Y(n7523) );
  NAND2X1 U7834 ( .A(G12), .B(n7491), .Y(n7522) );
  NAND4X1 U7835 ( .A(n7532), .B(n7533), .C(n7534), .D(n7535), .Y(G947) );
  NOR3X1 U7836 ( .A(n7536), .B(n7537), .C(n7538), .Y(n7535) );
  NOR2X1 U7837 ( .A(n7539), .B(n7484), .Y(n7538) );
  NOR2X1 U7838 ( .A(n7485), .B(n7540), .Y(n7537) );
  NOR2X1 U7839 ( .A(n7487), .B(n7541), .Y(n7536) );
  NAND2X1 U7840 ( .A(G27), .B(n7489), .Y(n7534) );
  NAND2X1 U7841 ( .A(G21551), .B(n7490), .Y(n7533) );
  NAND2X1 U7842 ( .A(G11), .B(n7491), .Y(n7532) );
  NAND4X1 U7843 ( .A(n7542), .B(n7543), .C(n7544), .D(n7545), .Y(G946) );
  NOR3X1 U7844 ( .A(n7546), .B(n7547), .C(n7548), .Y(n7545) );
  NOR2X1 U7845 ( .A(n7549), .B(n7484), .Y(n7548) );
  NOR2X1 U7846 ( .A(n7485), .B(n7550), .Y(n7547) );
  NOR2X1 U7847 ( .A(n7487), .B(n7551), .Y(n7546) );
  NAND2X1 U7848 ( .A(G26), .B(n7489), .Y(n7544) );
  NAND2X1 U7849 ( .A(G21550), .B(n7490), .Y(n7543) );
  NAND2X1 U7850 ( .A(G10), .B(n7491), .Y(n7542) );
  NAND4X1 U7851 ( .A(n7552), .B(n7553), .C(n7554), .D(n7555), .Y(G945) );
  NOR3X1 U7852 ( .A(n7556), .B(n7557), .C(n7558), .Y(n7555) );
  NOR2X1 U7853 ( .A(n7559), .B(n7484), .Y(n7558) );
  NOR2X1 U7854 ( .A(n7485), .B(n7560), .Y(n7557) );
  AND2X1 U7855 ( .A(n7561), .B(n7562), .Y(n7485) );
  NAND2X1 U7856 ( .A(n7563), .B(n7564), .Y(n7562) );
  NAND2X1 U7857 ( .A(n7565), .B(G21426), .Y(n7561) );
  NOR2X1 U7858 ( .A(n7487), .B(n7566), .Y(n7556) );
  NAND2X1 U7859 ( .A(G25), .B(n7489), .Y(n7554) );
  NAND2X1 U7860 ( .A(n7567), .B(n7568), .Y(n7489) );
  NAND4X1 U7861 ( .A(n7563), .B(n7569), .C(n7487), .D(n7570), .Y(n7568) );
  INVX1 U7862 ( .A(n7571), .Y(n7563) );
  NAND2X1 U7863 ( .A(n7572), .B(n7573), .Y(n7567) );
  NAND2X1 U7864 ( .A(G21549), .B(n7490), .Y(n7553) );
  NAND2X1 U7865 ( .A(n7574), .B(n7575), .Y(n7490) );
  NAND3X1 U7866 ( .A(n7576), .B(n7577), .C(n7578), .Y(n7575) );
  NAND2X1 U7867 ( .A(n7579), .B(n7565), .Y(n7578) );
  NAND2X1 U7868 ( .A(n7573), .B(n7580), .Y(n7576) );
  INVX1 U7869 ( .A(n7484), .Y(n7573) );
  NAND2X1 U7870 ( .A(n7572), .B(n7484), .Y(n7574) );
  NAND2X1 U7871 ( .A(n7581), .B(n7582), .Y(n7484) );
  AND2X1 U7872 ( .A(n7583), .B(n7571), .Y(n7572) );
  NAND2X1 U7873 ( .A(n7584), .B(n7585), .Y(n7571) );
  NAND2X1 U7874 ( .A(n7586), .B(n7587), .Y(n7583) );
  NAND3X1 U7875 ( .A(n7487), .B(n7570), .C(n7569), .Y(n7587) );
  NAND2X1 U7876 ( .A(G9), .B(n7491), .Y(n7552) );
  AND3X1 U7877 ( .A(n7565), .B(n7487), .C(n7569), .Y(n7491) );
  NAND4X1 U7878 ( .A(n7588), .B(n7589), .C(n7590), .D(n7591), .Y(G944) );
  NOR3X1 U7879 ( .A(n7592), .B(n7593), .C(n7594), .Y(n7591) );
  NOR2X1 U7880 ( .A(n7483), .B(n7595), .Y(n7594) );
  NOR2X1 U7881 ( .A(n7596), .B(n7486), .Y(n7593) );
  NOR2X1 U7882 ( .A(n7597), .B(n7488), .Y(n7592) );
  NAND2X1 U7883 ( .A(G32), .B(n7598), .Y(n7590) );
  NAND2X1 U7884 ( .A(G21548), .B(n7599), .Y(n7589) );
  NAND2X1 U7885 ( .A(n7600), .B(G16), .Y(n7588) );
  NAND4X1 U7886 ( .A(n7601), .B(n7602), .C(n7603), .D(n7604), .Y(G943) );
  NOR3X1 U7887 ( .A(n7605), .B(n7606), .C(n7607), .Y(n7604) );
  NOR2X1 U7888 ( .A(n7499), .B(n7595), .Y(n7607) );
  NOR2X1 U7889 ( .A(n7596), .B(n7500), .Y(n7606) );
  NOR2X1 U7890 ( .A(n7597), .B(n7501), .Y(n7605) );
  NAND2X1 U7891 ( .A(G31), .B(n7598), .Y(n7603) );
  NAND2X1 U7892 ( .A(G21547), .B(n7599), .Y(n7602) );
  NAND2X1 U7893 ( .A(n7600), .B(G15), .Y(n7601) );
  NAND4X1 U7894 ( .A(n7608), .B(n7609), .C(n7610), .D(n7611), .Y(G942) );
  NOR3X1 U7895 ( .A(n7612), .B(n7613), .C(n7614), .Y(n7611) );
  NOR2X1 U7896 ( .A(n7509), .B(n7595), .Y(n7614) );
  NOR2X1 U7897 ( .A(n7596), .B(n7510), .Y(n7613) );
  NOR2X1 U7898 ( .A(n7597), .B(n7511), .Y(n7612) );
  NAND2X1 U7899 ( .A(G30), .B(n7598), .Y(n7610) );
  NAND2X1 U7900 ( .A(G21546), .B(n7599), .Y(n7609) );
  NAND2X1 U7901 ( .A(n7600), .B(G14), .Y(n7608) );
  NAND4X1 U7902 ( .A(n7615), .B(n7616), .C(n7617), .D(n7618), .Y(G941) );
  NOR3X1 U7903 ( .A(n7619), .B(n7620), .C(n7621), .Y(n7618) );
  NOR2X1 U7904 ( .A(n7519), .B(n7595), .Y(n7621) );
  NOR2X1 U7905 ( .A(n7596), .B(n7520), .Y(n7620) );
  NOR2X1 U7906 ( .A(n7597), .B(n7521), .Y(n7619) );
  NAND2X1 U7907 ( .A(G29), .B(n7598), .Y(n7617) );
  NAND2X1 U7908 ( .A(G21545), .B(n7599), .Y(n7616) );
  NAND2X1 U7909 ( .A(n7600), .B(G13), .Y(n7615) );
  NAND4X1 U7910 ( .A(n7622), .B(n7623), .C(n7624), .D(n7625), .Y(G940) );
  NOR3X1 U7911 ( .A(n7626), .B(n7627), .C(n7628), .Y(n7625) );
  NOR2X1 U7912 ( .A(n7529), .B(n7595), .Y(n7628) );
  NOR2X1 U7913 ( .A(n7596), .B(n7530), .Y(n7627) );
  NOR2X1 U7914 ( .A(n7597), .B(n7531), .Y(n7626) );
  NAND2X1 U7915 ( .A(G28), .B(n7598), .Y(n7624) );
  NAND2X1 U7916 ( .A(G21544), .B(n7599), .Y(n7623) );
  NAND2X1 U7917 ( .A(n7600), .B(G12), .Y(n7622) );
  NAND4X1 U7918 ( .A(n7629), .B(n7630), .C(n7631), .D(n7632), .Y(G939) );
  NOR3X1 U7919 ( .A(n7633), .B(n7634), .C(n7635), .Y(n7632) );
  NOR2X1 U7920 ( .A(n7539), .B(n7595), .Y(n7635) );
  NOR2X1 U7921 ( .A(n7596), .B(n7540), .Y(n7634) );
  NOR2X1 U7922 ( .A(n7597), .B(n7541), .Y(n7633) );
  NAND2X1 U7923 ( .A(G27), .B(n7598), .Y(n7631) );
  NAND2X1 U7924 ( .A(G21543), .B(n7599), .Y(n7630) );
  NAND2X1 U7925 ( .A(n7600), .B(G11), .Y(n7629) );
  NAND4X1 U7926 ( .A(n7636), .B(n7637), .C(n7638), .D(n7639), .Y(G938) );
  NOR3X1 U7927 ( .A(n7640), .B(n7641), .C(n7642), .Y(n7639) );
  NOR2X1 U7928 ( .A(n7549), .B(n7595), .Y(n7642) );
  NOR2X1 U7929 ( .A(n7596), .B(n7550), .Y(n7641) );
  NOR2X1 U7930 ( .A(n7597), .B(n7551), .Y(n7640) );
  NAND2X1 U7931 ( .A(G26), .B(n7598), .Y(n7638) );
  NAND2X1 U7932 ( .A(G21542), .B(n7599), .Y(n7637) );
  NAND2X1 U7933 ( .A(n7600), .B(G10), .Y(n7636) );
  NAND4X1 U7934 ( .A(n7643), .B(n7644), .C(n7645), .D(n7646), .Y(G937) );
  NOR3X1 U7935 ( .A(n7647), .B(n7648), .C(n7649), .Y(n7646) );
  NOR2X1 U7936 ( .A(n7559), .B(n7595), .Y(n7649) );
  NOR2X1 U7937 ( .A(n7596), .B(n7560), .Y(n7648) );
  AND2X1 U7938 ( .A(n7650), .B(n7651), .Y(n7596) );
  NAND2X1 U7939 ( .A(n7652), .B(n7564), .Y(n7651) );
  NAND2X1 U7940 ( .A(n7653), .B(G21426), .Y(n7650) );
  NOR2X1 U7941 ( .A(n7597), .B(n7566), .Y(n7647) );
  NAND2X1 U7942 ( .A(G25), .B(n7598), .Y(n7645) );
  NAND2X1 U7943 ( .A(n7654), .B(n7655), .Y(n7598) );
  NAND4X1 U7944 ( .A(n7652), .B(n7569), .C(n7597), .D(n7656), .Y(n7655) );
  INVX1 U7945 ( .A(n7657), .Y(n7652) );
  NAND2X1 U7946 ( .A(n7658), .B(n7659), .Y(n7654) );
  NAND2X1 U7947 ( .A(G21541), .B(n7599), .Y(n7644) );
  NAND2X1 U7948 ( .A(n7660), .B(n7661), .Y(n7599) );
  NAND3X1 U7949 ( .A(n7662), .B(n7577), .C(n7663), .Y(n7661) );
  NAND2X1 U7950 ( .A(n7579), .B(n7653), .Y(n7663) );
  NAND2X1 U7951 ( .A(n7659), .B(n7580), .Y(n7662) );
  INVX1 U7952 ( .A(n7595), .Y(n7659) );
  NAND2X1 U7953 ( .A(n7658), .B(n7595), .Y(n7660) );
  NAND2X1 U7954 ( .A(n7664), .B(n7582), .Y(n7595) );
  AND2X1 U7955 ( .A(n7665), .B(n7657), .Y(n7658) );
  NAND2X1 U7956 ( .A(n7666), .B(n7585), .Y(n7657) );
  NAND2X1 U7957 ( .A(n7586), .B(n7667), .Y(n7665) );
  NAND3X1 U7958 ( .A(n7597), .B(n7656), .C(n7569), .Y(n7667) );
  NAND2X1 U7959 ( .A(n7600), .B(G9), .Y(n7643) );
  AND3X1 U7960 ( .A(n7653), .B(n7597), .C(n7569), .Y(n7600) );
  NAND4X1 U7961 ( .A(n7668), .B(n7669), .C(n7670), .D(n7671), .Y(G936) );
  NOR3X1 U7962 ( .A(n7672), .B(n7673), .C(n7674), .Y(n7671) );
  NOR2X1 U7963 ( .A(n7483), .B(n7675), .Y(n7674) );
  NOR2X1 U7964 ( .A(n7676), .B(n7486), .Y(n7673) );
  NOR2X1 U7965 ( .A(n7677), .B(n7488), .Y(n7672) );
  NAND2X1 U7966 ( .A(G32), .B(n7678), .Y(n7670) );
  NAND2X1 U7967 ( .A(G21540), .B(n7679), .Y(n7669) );
  NAND2X1 U7968 ( .A(n7680), .B(G16), .Y(n7668) );
  NAND4X1 U7969 ( .A(n7681), .B(n7682), .C(n7683), .D(n7684), .Y(G935) );
  NOR3X1 U7970 ( .A(n7685), .B(n7686), .C(n7687), .Y(n7684) );
  NOR2X1 U7971 ( .A(n7499), .B(n7675), .Y(n7687) );
  NOR2X1 U7972 ( .A(n7676), .B(n7500), .Y(n7686) );
  NOR2X1 U7973 ( .A(n7677), .B(n7501), .Y(n7685) );
  NAND2X1 U7974 ( .A(G31), .B(n7678), .Y(n7683) );
  NAND2X1 U7975 ( .A(G21539), .B(n7679), .Y(n7682) );
  NAND2X1 U7976 ( .A(n7680), .B(G15), .Y(n7681) );
  NAND4X1 U7977 ( .A(n7688), .B(n7689), .C(n7690), .D(n7691), .Y(G934) );
  NOR3X1 U7978 ( .A(n7692), .B(n7693), .C(n7694), .Y(n7691) );
  NOR2X1 U7979 ( .A(n7509), .B(n7675), .Y(n7694) );
  NOR2X1 U7980 ( .A(n7676), .B(n7510), .Y(n7693) );
  NOR2X1 U7981 ( .A(n7677), .B(n7511), .Y(n7692) );
  NAND2X1 U7982 ( .A(G30), .B(n7678), .Y(n7690) );
  NAND2X1 U7983 ( .A(G21538), .B(n7679), .Y(n7689) );
  NAND2X1 U7984 ( .A(n7680), .B(G14), .Y(n7688) );
  NAND4X1 U7985 ( .A(n7695), .B(n7696), .C(n7697), .D(n7698), .Y(G933) );
  NOR3X1 U7986 ( .A(n7699), .B(n7700), .C(n7701), .Y(n7698) );
  NOR2X1 U7987 ( .A(n7519), .B(n7675), .Y(n7701) );
  NOR2X1 U7988 ( .A(n7676), .B(n7520), .Y(n7700) );
  NOR2X1 U7989 ( .A(n7677), .B(n7521), .Y(n7699) );
  NAND2X1 U7990 ( .A(G29), .B(n7678), .Y(n7697) );
  NAND2X1 U7991 ( .A(G21537), .B(n7679), .Y(n7696) );
  NAND2X1 U7992 ( .A(n7680), .B(G13), .Y(n7695) );
  NAND4X1 U7993 ( .A(n7702), .B(n7703), .C(n7704), .D(n7705), .Y(G932) );
  NOR3X1 U7994 ( .A(n7706), .B(n7707), .C(n7708), .Y(n7705) );
  NOR2X1 U7995 ( .A(n7529), .B(n7675), .Y(n7708) );
  NOR2X1 U7996 ( .A(n7676), .B(n7530), .Y(n7707) );
  NOR2X1 U7997 ( .A(n7677), .B(n7531), .Y(n7706) );
  NAND2X1 U7998 ( .A(G28), .B(n7678), .Y(n7704) );
  NAND2X1 U7999 ( .A(G21536), .B(n7679), .Y(n7703) );
  NAND2X1 U8000 ( .A(n7680), .B(G12), .Y(n7702) );
  NAND4X1 U8001 ( .A(n7709), .B(n7710), .C(n7711), .D(n7712), .Y(G931) );
  NOR3X1 U8002 ( .A(n7713), .B(n7714), .C(n7715), .Y(n7712) );
  NOR2X1 U8003 ( .A(n7539), .B(n7675), .Y(n7715) );
  NOR2X1 U8004 ( .A(n7676), .B(n7540), .Y(n7714) );
  NOR2X1 U8005 ( .A(n7677), .B(n7541), .Y(n7713) );
  NAND2X1 U8006 ( .A(G27), .B(n7678), .Y(n7711) );
  NAND2X1 U8007 ( .A(G21535), .B(n7679), .Y(n7710) );
  NAND2X1 U8008 ( .A(n7680), .B(G11), .Y(n7709) );
  NAND4X1 U8009 ( .A(n7716), .B(n7717), .C(n7718), .D(n7719), .Y(G930) );
  NOR3X1 U8010 ( .A(n7720), .B(n7721), .C(n7722), .Y(n7719) );
  NOR2X1 U8011 ( .A(n7549), .B(n7675), .Y(n7722) );
  NOR2X1 U8012 ( .A(n7676), .B(n7550), .Y(n7721) );
  NOR2X1 U8013 ( .A(n7677), .B(n7551), .Y(n7720) );
  NAND2X1 U8014 ( .A(G26), .B(n7678), .Y(n7718) );
  NAND2X1 U8015 ( .A(G21534), .B(n7679), .Y(n7717) );
  NAND2X1 U8016 ( .A(n7680), .B(G10), .Y(n7716) );
  NAND4X1 U8017 ( .A(n7723), .B(n7724), .C(n7725), .D(n7726), .Y(G929) );
  NOR3X1 U8018 ( .A(n7727), .B(n7728), .C(n7729), .Y(n7726) );
  NOR2X1 U8019 ( .A(n7559), .B(n7675), .Y(n7729) );
  NOR2X1 U8020 ( .A(n7676), .B(n7560), .Y(n7728) );
  AND2X1 U8021 ( .A(n7730), .B(n7731), .Y(n7676) );
  NAND2X1 U8022 ( .A(n7732), .B(n7564), .Y(n7731) );
  NAND2X1 U8023 ( .A(n7733), .B(G21426), .Y(n7730) );
  NOR2X1 U8024 ( .A(n7677), .B(n7566), .Y(n7727) );
  NAND2X1 U8025 ( .A(G25), .B(n7678), .Y(n7725) );
  NAND2X1 U8026 ( .A(n7734), .B(n7735), .Y(n7678) );
  NAND4X1 U8027 ( .A(n7732), .B(n7569), .C(n7677), .D(n7736), .Y(n7735) );
  INVX1 U8028 ( .A(n7737), .Y(n7732) );
  NAND2X1 U8029 ( .A(n7738), .B(n7739), .Y(n7734) );
  NAND2X1 U8030 ( .A(G21533), .B(n7679), .Y(n7724) );
  NAND2X1 U8031 ( .A(n7740), .B(n7741), .Y(n7679) );
  NAND3X1 U8032 ( .A(n7742), .B(n7577), .C(n7743), .Y(n7741) );
  NAND2X1 U8033 ( .A(n7579), .B(n7733), .Y(n7743) );
  NAND2X1 U8034 ( .A(n7739), .B(n7580), .Y(n7742) );
  INVX1 U8035 ( .A(n7675), .Y(n7739) );
  NAND2X1 U8036 ( .A(n7738), .B(n7675), .Y(n7740) );
  NAND2X1 U8037 ( .A(n7744), .B(n7582), .Y(n7675) );
  AND2X1 U8038 ( .A(n7745), .B(n7737), .Y(n7738) );
  NAND2X1 U8039 ( .A(n7746), .B(n7585), .Y(n7737) );
  NAND2X1 U8040 ( .A(n7586), .B(n7747), .Y(n7745) );
  NAND3X1 U8041 ( .A(n7677), .B(n7736), .C(n7569), .Y(n7747) );
  NAND2X1 U8042 ( .A(n7680), .B(G9), .Y(n7723) );
  AND3X1 U8043 ( .A(n7733), .B(n7677), .C(n7569), .Y(n7680) );
  NAND4X1 U8044 ( .A(n7748), .B(n7749), .C(n7750), .D(n7751), .Y(G928) );
  NOR3X1 U8045 ( .A(n7752), .B(n7753), .C(n7754), .Y(n7751) );
  NOR2X1 U8046 ( .A(n7483), .B(n7755), .Y(n7754) );
  NOR2X1 U8047 ( .A(n7756), .B(n7486), .Y(n7753) );
  NOR2X1 U8048 ( .A(n7757), .B(n7488), .Y(n7752) );
  NAND2X1 U8049 ( .A(G32), .B(n7758), .Y(n7750) );
  NAND2X1 U8050 ( .A(G21532), .B(n7759), .Y(n7749) );
  NAND2X1 U8051 ( .A(n7760), .B(G16), .Y(n7748) );
  NAND4X1 U8052 ( .A(n7761), .B(n7762), .C(n7763), .D(n7764), .Y(G927) );
  NOR3X1 U8053 ( .A(n7765), .B(n7766), .C(n7767), .Y(n7764) );
  NOR2X1 U8054 ( .A(n7499), .B(n7755), .Y(n7767) );
  NOR2X1 U8055 ( .A(n7756), .B(n7500), .Y(n7766) );
  NOR2X1 U8056 ( .A(n7757), .B(n7501), .Y(n7765) );
  NAND2X1 U8057 ( .A(G31), .B(n7758), .Y(n7763) );
  NAND2X1 U8058 ( .A(G21531), .B(n7759), .Y(n7762) );
  NAND2X1 U8059 ( .A(n7760), .B(G15), .Y(n7761) );
  NAND4X1 U8060 ( .A(n7768), .B(n7769), .C(n7770), .D(n7771), .Y(G926) );
  NOR3X1 U8061 ( .A(n7772), .B(n7773), .C(n7774), .Y(n7771) );
  NOR2X1 U8062 ( .A(n7509), .B(n7755), .Y(n7774) );
  NOR2X1 U8063 ( .A(n7756), .B(n7510), .Y(n7773) );
  NOR2X1 U8064 ( .A(n7757), .B(n7511), .Y(n7772) );
  NAND2X1 U8065 ( .A(G30), .B(n7758), .Y(n7770) );
  NAND2X1 U8066 ( .A(G21530), .B(n7759), .Y(n7769) );
  NAND2X1 U8067 ( .A(n7760), .B(G14), .Y(n7768) );
  NAND4X1 U8068 ( .A(n7775), .B(n7776), .C(n7777), .D(n7778), .Y(G925) );
  NOR3X1 U8069 ( .A(n7779), .B(n7780), .C(n7781), .Y(n7778) );
  NOR2X1 U8070 ( .A(n7519), .B(n7755), .Y(n7781) );
  NOR2X1 U8071 ( .A(n7756), .B(n7520), .Y(n7780) );
  NOR2X1 U8072 ( .A(n7757), .B(n7521), .Y(n7779) );
  NAND2X1 U8073 ( .A(G29), .B(n7758), .Y(n7777) );
  NAND2X1 U8074 ( .A(G21529), .B(n7759), .Y(n7776) );
  NAND2X1 U8075 ( .A(n7760), .B(G13), .Y(n7775) );
  NAND4X1 U8076 ( .A(n7782), .B(n7783), .C(n7784), .D(n7785), .Y(G924) );
  NOR3X1 U8077 ( .A(n7786), .B(n7787), .C(n7788), .Y(n7785) );
  NOR2X1 U8078 ( .A(n7529), .B(n7755), .Y(n7788) );
  NOR2X1 U8079 ( .A(n7756), .B(n7530), .Y(n7787) );
  NOR2X1 U8080 ( .A(n7757), .B(n7531), .Y(n7786) );
  NAND2X1 U8081 ( .A(G28), .B(n7758), .Y(n7784) );
  NAND2X1 U8082 ( .A(G21528), .B(n7759), .Y(n7783) );
  NAND2X1 U8083 ( .A(n7760), .B(G12), .Y(n7782) );
  NAND4X1 U8084 ( .A(n7789), .B(n7790), .C(n7791), .D(n7792), .Y(G923) );
  NOR3X1 U8085 ( .A(n7793), .B(n7794), .C(n7795), .Y(n7792) );
  NOR2X1 U8086 ( .A(n7539), .B(n7755), .Y(n7795) );
  NOR2X1 U8087 ( .A(n7756), .B(n7540), .Y(n7794) );
  NOR2X1 U8088 ( .A(n7757), .B(n7541), .Y(n7793) );
  NAND2X1 U8089 ( .A(G27), .B(n7758), .Y(n7791) );
  NAND2X1 U8090 ( .A(G21527), .B(n7759), .Y(n7790) );
  NAND2X1 U8091 ( .A(n7760), .B(G11), .Y(n7789) );
  NAND4X1 U8092 ( .A(n7796), .B(n7797), .C(n7798), .D(n7799), .Y(G922) );
  NOR3X1 U8093 ( .A(n7800), .B(n7801), .C(n7802), .Y(n7799) );
  NOR2X1 U8094 ( .A(n7549), .B(n7755), .Y(n7802) );
  NOR2X1 U8095 ( .A(n7756), .B(n7550), .Y(n7801) );
  NOR2X1 U8096 ( .A(n7757), .B(n7551), .Y(n7800) );
  NAND2X1 U8097 ( .A(G26), .B(n7758), .Y(n7798) );
  NAND2X1 U8098 ( .A(G21526), .B(n7759), .Y(n7797) );
  NAND2X1 U8099 ( .A(n7760), .B(G10), .Y(n7796) );
  NAND4X1 U8100 ( .A(n7803), .B(n7804), .C(n7805), .D(n7806), .Y(G921) );
  NOR3X1 U8101 ( .A(n7807), .B(n7808), .C(n7809), .Y(n7806) );
  NOR2X1 U8102 ( .A(n7559), .B(n7755), .Y(n7809) );
  NOR2X1 U8103 ( .A(n7756), .B(n7560), .Y(n7808) );
  AND2X1 U8104 ( .A(n7810), .B(n7811), .Y(n7756) );
  NAND2X1 U8105 ( .A(n7812), .B(n7564), .Y(n7811) );
  NAND2X1 U8106 ( .A(n7813), .B(G21426), .Y(n7810) );
  NOR2X1 U8107 ( .A(n7757), .B(n7566), .Y(n7807) );
  NAND2X1 U8108 ( .A(G25), .B(n7758), .Y(n7805) );
  NAND2X1 U8109 ( .A(n7814), .B(n7815), .Y(n7758) );
  NAND4X1 U8110 ( .A(n7812), .B(n7569), .C(n7757), .D(n7816), .Y(n7815) );
  INVX1 U8111 ( .A(n7817), .Y(n7812) );
  NAND2X1 U8112 ( .A(n7818), .B(n7819), .Y(n7814) );
  NAND2X1 U8113 ( .A(G21525), .B(n7759), .Y(n7804) );
  NAND2X1 U8114 ( .A(n7820), .B(n7821), .Y(n7759) );
  NAND3X1 U8115 ( .A(n7822), .B(n7577), .C(n7823), .Y(n7821) );
  NAND2X1 U8116 ( .A(n7579), .B(n7813), .Y(n7823) );
  NAND2X1 U8117 ( .A(n7819), .B(n7580), .Y(n7822) );
  INVX1 U8118 ( .A(n7755), .Y(n7819) );
  NAND2X1 U8119 ( .A(n7818), .B(n7755), .Y(n7820) );
  NAND2X1 U8120 ( .A(n7582), .B(n7824), .Y(n7755) );
  NOR2X1 U8121 ( .A(G21564), .B(G21563), .Y(n7582) );
  AND2X1 U8122 ( .A(n7825), .B(n7817), .Y(n7818) );
  NAND2X1 U8123 ( .A(n7826), .B(n7585), .Y(n7817) );
  NOR2X1 U8124 ( .A(n7827), .B(n7828), .Y(n7585) );
  NAND2X1 U8125 ( .A(n7586), .B(n7829), .Y(n7825) );
  NAND3X1 U8126 ( .A(n7757), .B(n7816), .C(n7569), .Y(n7829) );
  NAND2X1 U8127 ( .A(n7760), .B(G9), .Y(n7803) );
  AND3X1 U8128 ( .A(n7813), .B(n7757), .C(n7569), .Y(n7760) );
  NAND4X1 U8129 ( .A(n7830), .B(n7831), .C(n7832), .D(n7833), .Y(G920) );
  NOR3X1 U8130 ( .A(n7834), .B(n7835), .C(n7836), .Y(n7833) );
  NOR2X1 U8131 ( .A(n7483), .B(n7837), .Y(n7836) );
  NOR2X1 U8132 ( .A(n7838), .B(n7486), .Y(n7835) );
  NOR2X1 U8133 ( .A(n7839), .B(n7488), .Y(n7834) );
  NAND2X1 U8134 ( .A(G32), .B(n7840), .Y(n7832) );
  NAND2X1 U8135 ( .A(G21524), .B(n7841), .Y(n7831) );
  NAND2X1 U8136 ( .A(n7842), .B(G16), .Y(n7830) );
  NAND4X1 U8137 ( .A(n7843), .B(n7844), .C(n7845), .D(n7846), .Y(G919) );
  NOR3X1 U8138 ( .A(n7847), .B(n7848), .C(n7849), .Y(n7846) );
  NOR2X1 U8139 ( .A(n7499), .B(n7837), .Y(n7849) );
  NOR2X1 U8140 ( .A(n7838), .B(n7500), .Y(n7848) );
  NOR2X1 U8141 ( .A(n7839), .B(n7501), .Y(n7847) );
  NAND2X1 U8142 ( .A(G31), .B(n7840), .Y(n7845) );
  NAND2X1 U8143 ( .A(G21523), .B(n7841), .Y(n7844) );
  NAND2X1 U8144 ( .A(n7842), .B(G15), .Y(n7843) );
  NAND4X1 U8145 ( .A(n7850), .B(n7851), .C(n7852), .D(n7853), .Y(G918) );
  NOR3X1 U8146 ( .A(n7854), .B(n7855), .C(n7856), .Y(n7853) );
  NOR2X1 U8147 ( .A(n7509), .B(n7837), .Y(n7856) );
  NOR2X1 U8148 ( .A(n7838), .B(n7510), .Y(n7855) );
  NOR2X1 U8149 ( .A(n7839), .B(n7511), .Y(n7854) );
  NAND2X1 U8150 ( .A(G30), .B(n7840), .Y(n7852) );
  NAND2X1 U8151 ( .A(G21522), .B(n7841), .Y(n7851) );
  NAND2X1 U8152 ( .A(n7842), .B(G14), .Y(n7850) );
  NAND4X1 U8153 ( .A(n7857), .B(n7858), .C(n7859), .D(n7860), .Y(G917) );
  NOR3X1 U8154 ( .A(n7861), .B(n7862), .C(n7863), .Y(n7860) );
  NOR2X1 U8155 ( .A(n7519), .B(n7837), .Y(n7863) );
  NOR2X1 U8156 ( .A(n7838), .B(n7520), .Y(n7862) );
  NOR2X1 U8157 ( .A(n7839), .B(n7521), .Y(n7861) );
  NAND2X1 U8158 ( .A(G29), .B(n7840), .Y(n7859) );
  NAND2X1 U8159 ( .A(G21521), .B(n7841), .Y(n7858) );
  NAND2X1 U8160 ( .A(n7842), .B(G13), .Y(n7857) );
  NAND4X1 U8161 ( .A(n7864), .B(n7865), .C(n7866), .D(n7867), .Y(G916) );
  NOR3X1 U8162 ( .A(n7868), .B(n7869), .C(n7870), .Y(n7867) );
  NOR2X1 U8163 ( .A(n7529), .B(n7837), .Y(n7870) );
  NOR2X1 U8164 ( .A(n7838), .B(n7530), .Y(n7869) );
  NOR2X1 U8165 ( .A(n7839), .B(n7531), .Y(n7868) );
  NAND2X1 U8166 ( .A(G28), .B(n7840), .Y(n7866) );
  NAND2X1 U8167 ( .A(G21520), .B(n7841), .Y(n7865) );
  NAND2X1 U8168 ( .A(n7842), .B(G12), .Y(n7864) );
  NAND4X1 U8169 ( .A(n7871), .B(n7872), .C(n7873), .D(n7874), .Y(G915) );
  NOR3X1 U8170 ( .A(n7875), .B(n7876), .C(n7877), .Y(n7874) );
  NOR2X1 U8171 ( .A(n7539), .B(n7837), .Y(n7877) );
  NOR2X1 U8172 ( .A(n7838), .B(n7540), .Y(n7876) );
  NOR2X1 U8173 ( .A(n7839), .B(n7541), .Y(n7875) );
  NAND2X1 U8174 ( .A(G27), .B(n7840), .Y(n7873) );
  NAND2X1 U8175 ( .A(G21519), .B(n7841), .Y(n7872) );
  NAND2X1 U8176 ( .A(n7842), .B(G11), .Y(n7871) );
  NAND4X1 U8177 ( .A(n7878), .B(n7879), .C(n7880), .D(n7881), .Y(G914) );
  NOR3X1 U8178 ( .A(n7882), .B(n7883), .C(n7884), .Y(n7881) );
  NOR2X1 U8179 ( .A(n7549), .B(n7837), .Y(n7884) );
  NOR2X1 U8180 ( .A(n7838), .B(n7550), .Y(n7883) );
  NOR2X1 U8181 ( .A(n7839), .B(n7551), .Y(n7882) );
  NAND2X1 U8182 ( .A(G26), .B(n7840), .Y(n7880) );
  NAND2X1 U8183 ( .A(G21518), .B(n7841), .Y(n7879) );
  NAND2X1 U8184 ( .A(n7842), .B(G10), .Y(n7878) );
  NAND4X1 U8185 ( .A(n7885), .B(n7886), .C(n7887), .D(n7888), .Y(G913) );
  NOR3X1 U8186 ( .A(n7889), .B(n7890), .C(n7891), .Y(n7888) );
  NOR2X1 U8187 ( .A(n7559), .B(n7837), .Y(n7891) );
  NOR2X1 U8188 ( .A(n7838), .B(n7560), .Y(n7890) );
  AND2X1 U8189 ( .A(n7892), .B(n7893), .Y(n7838) );
  NAND2X1 U8190 ( .A(n7894), .B(n7564), .Y(n7893) );
  NAND2X1 U8191 ( .A(n7895), .B(G21426), .Y(n7892) );
  NOR2X1 U8192 ( .A(n7839), .B(n7566), .Y(n7889) );
  NAND2X1 U8193 ( .A(G25), .B(n7840), .Y(n7887) );
  NAND2X1 U8194 ( .A(n7896), .B(n7897), .Y(n7840) );
  NAND4X1 U8195 ( .A(n7894), .B(n7569), .C(n7839), .D(n7898), .Y(n7897) );
  INVX1 U8196 ( .A(n7899), .Y(n7894) );
  NAND2X1 U8197 ( .A(n7900), .B(n7901), .Y(n7896) );
  NAND2X1 U8198 ( .A(G21517), .B(n7841), .Y(n7886) );
  NAND2X1 U8199 ( .A(n7902), .B(n7903), .Y(n7841) );
  NAND3X1 U8200 ( .A(n7904), .B(n7577), .C(n7905), .Y(n7903) );
  NAND2X1 U8201 ( .A(n7579), .B(n7895), .Y(n7905) );
  NAND2X1 U8202 ( .A(n7901), .B(n7580), .Y(n7904) );
  INVX1 U8203 ( .A(n7837), .Y(n7901) );
  NAND2X1 U8204 ( .A(n7900), .B(n7837), .Y(n7902) );
  NAND2X1 U8205 ( .A(n7581), .B(n7906), .Y(n7837) );
  AND2X1 U8206 ( .A(n7907), .B(n7899), .Y(n7900) );
  NAND2X1 U8207 ( .A(n7908), .B(n7584), .Y(n7899) );
  NAND2X1 U8208 ( .A(n7586), .B(n7909), .Y(n7907) );
  NAND3X1 U8209 ( .A(n7839), .B(n7898), .C(n7569), .Y(n7909) );
  NAND2X1 U8210 ( .A(n7842), .B(G9), .Y(n7885) );
  AND3X1 U8211 ( .A(n7895), .B(n7839), .C(n7569), .Y(n7842) );
  NAND4X1 U8212 ( .A(n7910), .B(n7911), .C(n7912), .D(n7913), .Y(G912) );
  NOR3X1 U8213 ( .A(n7914), .B(n7915), .C(n7916), .Y(n7913) );
  NOR2X1 U8214 ( .A(n7483), .B(n7917), .Y(n7916) );
  NOR2X1 U8215 ( .A(n7918), .B(n7486), .Y(n7915) );
  NOR2X1 U8216 ( .A(n7919), .B(n7488), .Y(n7914) );
  NAND2X1 U8217 ( .A(G32), .B(n7920), .Y(n7912) );
  NAND2X1 U8218 ( .A(G21516), .B(n7921), .Y(n7911) );
  NAND2X1 U8219 ( .A(n7922), .B(G16), .Y(n7910) );
  NAND4X1 U8220 ( .A(n7923), .B(n7924), .C(n7925), .D(n7926), .Y(G911) );
  NOR3X1 U8221 ( .A(n7927), .B(n7928), .C(n7929), .Y(n7926) );
  NOR2X1 U8222 ( .A(n7499), .B(n7917), .Y(n7929) );
  NOR2X1 U8223 ( .A(n7918), .B(n7500), .Y(n7928) );
  NOR2X1 U8224 ( .A(n7919), .B(n7501), .Y(n7927) );
  NAND2X1 U8225 ( .A(G31), .B(n7920), .Y(n7925) );
  NAND2X1 U8226 ( .A(G21515), .B(n7921), .Y(n7924) );
  NAND2X1 U8227 ( .A(n7922), .B(G15), .Y(n7923) );
  NAND4X1 U8228 ( .A(n7930), .B(n7931), .C(n7932), .D(n7933), .Y(G910) );
  NOR3X1 U8229 ( .A(n7934), .B(n7935), .C(n7936), .Y(n7933) );
  NOR2X1 U8230 ( .A(n7509), .B(n7917), .Y(n7936) );
  NOR2X1 U8231 ( .A(n7918), .B(n7510), .Y(n7935) );
  NOR2X1 U8232 ( .A(n7919), .B(n7511), .Y(n7934) );
  NAND2X1 U8233 ( .A(G30), .B(n7920), .Y(n7932) );
  NAND2X1 U8234 ( .A(G21514), .B(n7921), .Y(n7931) );
  NAND2X1 U8235 ( .A(n7922), .B(G14), .Y(n7930) );
  NAND4X1 U8236 ( .A(n7937), .B(n7938), .C(n7939), .D(n7940), .Y(G909) );
  NOR3X1 U8237 ( .A(n7941), .B(n7942), .C(n7943), .Y(n7940) );
  NOR2X1 U8238 ( .A(n7519), .B(n7917), .Y(n7943) );
  NOR2X1 U8239 ( .A(n7918), .B(n7520), .Y(n7942) );
  NOR2X1 U8240 ( .A(n7919), .B(n7521), .Y(n7941) );
  NAND2X1 U8241 ( .A(G29), .B(n7920), .Y(n7939) );
  NAND2X1 U8242 ( .A(G21513), .B(n7921), .Y(n7938) );
  NAND2X1 U8243 ( .A(n7922), .B(G13), .Y(n7937) );
  NAND4X1 U8244 ( .A(n7944), .B(n7945), .C(n7946), .D(n7947), .Y(G908) );
  NOR3X1 U8245 ( .A(n7948), .B(n7949), .C(n7950), .Y(n7947) );
  NOR2X1 U8246 ( .A(n7529), .B(n7917), .Y(n7950) );
  NOR2X1 U8247 ( .A(n7918), .B(n7530), .Y(n7949) );
  NOR2X1 U8248 ( .A(n7919), .B(n7531), .Y(n7948) );
  NAND2X1 U8249 ( .A(G28), .B(n7920), .Y(n7946) );
  NAND2X1 U8250 ( .A(G21512), .B(n7921), .Y(n7945) );
  NAND2X1 U8251 ( .A(n7922), .B(G12), .Y(n7944) );
  NAND4X1 U8252 ( .A(n7951), .B(n7952), .C(n7953), .D(n7954), .Y(G907) );
  NOR3X1 U8253 ( .A(n7955), .B(n7956), .C(n7957), .Y(n7954) );
  NOR2X1 U8254 ( .A(n7539), .B(n7917), .Y(n7957) );
  NOR2X1 U8255 ( .A(n7918), .B(n7540), .Y(n7956) );
  NOR2X1 U8256 ( .A(n7919), .B(n7541), .Y(n7955) );
  NAND2X1 U8257 ( .A(G27), .B(n7920), .Y(n7953) );
  NAND2X1 U8258 ( .A(G21511), .B(n7921), .Y(n7952) );
  NAND2X1 U8259 ( .A(n7922), .B(G11), .Y(n7951) );
  NAND4X1 U8260 ( .A(n7958), .B(n7959), .C(n7960), .D(n7961), .Y(G906) );
  NOR3X1 U8261 ( .A(n7962), .B(n7963), .C(n7964), .Y(n7961) );
  NOR2X1 U8262 ( .A(n7549), .B(n7917), .Y(n7964) );
  NOR2X1 U8263 ( .A(n7918), .B(n7550), .Y(n7963) );
  NOR2X1 U8264 ( .A(n7919), .B(n7551), .Y(n7962) );
  NAND2X1 U8265 ( .A(G26), .B(n7920), .Y(n7960) );
  NAND2X1 U8266 ( .A(G21510), .B(n7921), .Y(n7959) );
  NAND2X1 U8267 ( .A(n7922), .B(G10), .Y(n7958) );
  NAND4X1 U8268 ( .A(n7965), .B(n7966), .C(n7967), .D(n7968), .Y(G905) );
  NOR3X1 U8269 ( .A(n7969), .B(n7970), .C(n7971), .Y(n7968) );
  NOR2X1 U8270 ( .A(n7559), .B(n7917), .Y(n7971) );
  NOR2X1 U8271 ( .A(n7918), .B(n7560), .Y(n7970) );
  AND2X1 U8272 ( .A(n7972), .B(n7973), .Y(n7918) );
  NAND2X1 U8273 ( .A(n7974), .B(n7564), .Y(n7973) );
  NAND2X1 U8274 ( .A(n7975), .B(G21426), .Y(n7972) );
  NOR2X1 U8275 ( .A(n7919), .B(n7566), .Y(n7969) );
  NAND2X1 U8276 ( .A(G25), .B(n7920), .Y(n7967) );
  NAND2X1 U8277 ( .A(n7976), .B(n7977), .Y(n7920) );
  NAND4X1 U8278 ( .A(n7974), .B(n7569), .C(n7919), .D(n7978), .Y(n7977) );
  INVX1 U8279 ( .A(n7979), .Y(n7974) );
  NAND2X1 U8280 ( .A(n7980), .B(n7981), .Y(n7976) );
  NAND2X1 U8281 ( .A(G21509), .B(n7921), .Y(n7966) );
  NAND2X1 U8282 ( .A(n7982), .B(n7983), .Y(n7921) );
  NAND3X1 U8283 ( .A(n7984), .B(n7577), .C(n7985), .Y(n7983) );
  NAND2X1 U8284 ( .A(n7579), .B(n7975), .Y(n7985) );
  NAND2X1 U8285 ( .A(n7981), .B(n7580), .Y(n7984) );
  INVX1 U8286 ( .A(n7917), .Y(n7981) );
  NAND2X1 U8287 ( .A(n7980), .B(n7917), .Y(n7982) );
  NAND2X1 U8288 ( .A(n7664), .B(n7906), .Y(n7917) );
  AND2X1 U8289 ( .A(n7986), .B(n7979), .Y(n7980) );
  NAND2X1 U8290 ( .A(n7908), .B(n7666), .Y(n7979) );
  NAND2X1 U8291 ( .A(n7586), .B(n7987), .Y(n7986) );
  NAND3X1 U8292 ( .A(n7919), .B(n7978), .C(n7569), .Y(n7987) );
  NAND2X1 U8293 ( .A(n7922), .B(G9), .Y(n7965) );
  AND3X1 U8294 ( .A(n7975), .B(n7919), .C(n7569), .Y(n7922) );
  NAND4X1 U8295 ( .A(n7988), .B(n7989), .C(n7990), .D(n7991), .Y(G904) );
  NOR3X1 U8296 ( .A(n7992), .B(n7993), .C(n7994), .Y(n7991) );
  NOR2X1 U8297 ( .A(n7483), .B(n7995), .Y(n7994) );
  NOR2X1 U8298 ( .A(n7996), .B(n7486), .Y(n7993) );
  NOR2X1 U8299 ( .A(n7997), .B(n7488), .Y(n7992) );
  NAND2X1 U8300 ( .A(G32), .B(n7998), .Y(n7990) );
  NAND2X1 U8301 ( .A(G21508), .B(n7999), .Y(n7989) );
  NAND2X1 U8302 ( .A(n8000), .B(G16), .Y(n7988) );
  NAND4X1 U8303 ( .A(n8001), .B(n8002), .C(n8003), .D(n8004), .Y(G903) );
  NOR3X1 U8304 ( .A(n8005), .B(n8006), .C(n8007), .Y(n8004) );
  NOR2X1 U8305 ( .A(n7499), .B(n7995), .Y(n8007) );
  NOR2X1 U8306 ( .A(n7996), .B(n7500), .Y(n8006) );
  NOR2X1 U8307 ( .A(n7997), .B(n7501), .Y(n8005) );
  NAND2X1 U8308 ( .A(G31), .B(n7998), .Y(n8003) );
  NAND2X1 U8309 ( .A(G21507), .B(n7999), .Y(n8002) );
  NAND2X1 U8310 ( .A(n8000), .B(G15), .Y(n8001) );
  NAND4X1 U8311 ( .A(n8008), .B(n8009), .C(n8010), .D(n8011), .Y(G902) );
  NOR3X1 U8312 ( .A(n8012), .B(n8013), .C(n8014), .Y(n8011) );
  NOR2X1 U8313 ( .A(n7509), .B(n7995), .Y(n8014) );
  NOR2X1 U8314 ( .A(n7996), .B(n7510), .Y(n8013) );
  NOR2X1 U8315 ( .A(n7997), .B(n7511), .Y(n8012) );
  NAND2X1 U8316 ( .A(G30), .B(n7998), .Y(n8010) );
  NAND2X1 U8317 ( .A(G21506), .B(n7999), .Y(n8009) );
  NAND2X1 U8318 ( .A(n8000), .B(G14), .Y(n8008) );
  NAND4X1 U8319 ( .A(n8015), .B(n8016), .C(n8017), .D(n8018), .Y(G901) );
  NOR3X1 U8320 ( .A(n8019), .B(n8020), .C(n8021), .Y(n8018) );
  NOR2X1 U8321 ( .A(n7519), .B(n7995), .Y(n8021) );
  NOR2X1 U8322 ( .A(n7996), .B(n7520), .Y(n8020) );
  NOR2X1 U8323 ( .A(n7997), .B(n7521), .Y(n8019) );
  NAND2X1 U8324 ( .A(G29), .B(n7998), .Y(n8017) );
  NAND2X1 U8325 ( .A(G21505), .B(n7999), .Y(n8016) );
  NAND2X1 U8326 ( .A(n8000), .B(G13), .Y(n8015) );
  NAND4X1 U8327 ( .A(n8022), .B(n8023), .C(n8024), .D(n8025), .Y(G900) );
  NOR3X1 U8328 ( .A(n8026), .B(n8027), .C(n8028), .Y(n8025) );
  NOR2X1 U8329 ( .A(n7529), .B(n7995), .Y(n8028) );
  NOR2X1 U8330 ( .A(n7996), .B(n7530), .Y(n8027) );
  NOR2X1 U8331 ( .A(n7997), .B(n7531), .Y(n8026) );
  NAND2X1 U8332 ( .A(G28), .B(n7998), .Y(n8024) );
  NAND2X1 U8333 ( .A(G21504), .B(n7999), .Y(n8023) );
  NAND2X1 U8334 ( .A(n8000), .B(G12), .Y(n8022) );
  NAND4X1 U8335 ( .A(n8029), .B(n8030), .C(n8031), .D(n8032), .Y(G899) );
  NOR3X1 U8336 ( .A(n8033), .B(n8034), .C(n8035), .Y(n8032) );
  NOR2X1 U8337 ( .A(n7539), .B(n7995), .Y(n8035) );
  NOR2X1 U8338 ( .A(n7996), .B(n7540), .Y(n8034) );
  NOR2X1 U8339 ( .A(n7997), .B(n7541), .Y(n8033) );
  NAND2X1 U8340 ( .A(G27), .B(n7998), .Y(n8031) );
  NAND2X1 U8341 ( .A(G21503), .B(n7999), .Y(n8030) );
  NAND2X1 U8342 ( .A(n8000), .B(G11), .Y(n8029) );
  NAND4X1 U8343 ( .A(n8036), .B(n8037), .C(n8038), .D(n8039), .Y(G898) );
  NOR3X1 U8344 ( .A(n8040), .B(n8041), .C(n8042), .Y(n8039) );
  NOR2X1 U8345 ( .A(n7549), .B(n7995), .Y(n8042) );
  NOR2X1 U8346 ( .A(n7996), .B(n7550), .Y(n8041) );
  NOR2X1 U8347 ( .A(n7997), .B(n7551), .Y(n8040) );
  NAND2X1 U8348 ( .A(G26), .B(n7998), .Y(n8038) );
  NAND2X1 U8349 ( .A(G21502), .B(n7999), .Y(n8037) );
  NAND2X1 U8350 ( .A(n8000), .B(G10), .Y(n8036) );
  NAND4X1 U8351 ( .A(n8043), .B(n8044), .C(n8045), .D(n8046), .Y(G897) );
  NOR3X1 U8352 ( .A(n8047), .B(n8048), .C(n8049), .Y(n8046) );
  NOR2X1 U8353 ( .A(n7559), .B(n7995), .Y(n8049) );
  NOR2X1 U8354 ( .A(n7996), .B(n7560), .Y(n8048) );
  AND2X1 U8355 ( .A(n8050), .B(n8051), .Y(n7996) );
  NAND2X1 U8356 ( .A(n8052), .B(n7564), .Y(n8051) );
  NAND2X1 U8357 ( .A(n8053), .B(G21426), .Y(n8050) );
  NOR2X1 U8358 ( .A(n7997), .B(n7566), .Y(n8047) );
  NAND2X1 U8359 ( .A(G25), .B(n7998), .Y(n8045) );
  NAND2X1 U8360 ( .A(n8054), .B(n8055), .Y(n7998) );
  NAND4X1 U8361 ( .A(n8052), .B(n7569), .C(n7997), .D(n8056), .Y(n8055) );
  INVX1 U8362 ( .A(n8057), .Y(n8052) );
  NAND2X1 U8363 ( .A(n8058), .B(n8059), .Y(n8054) );
  NAND2X1 U8364 ( .A(G21501), .B(n7999), .Y(n8044) );
  NAND2X1 U8365 ( .A(n8060), .B(n8061), .Y(n7999) );
  NAND3X1 U8366 ( .A(n8062), .B(n7577), .C(n8063), .Y(n8061) );
  NAND2X1 U8367 ( .A(n7579), .B(n8053), .Y(n8063) );
  NAND2X1 U8368 ( .A(n8059), .B(n7580), .Y(n8062) );
  INVX1 U8369 ( .A(n7995), .Y(n8059) );
  NAND2X1 U8370 ( .A(n8058), .B(n7995), .Y(n8060) );
  NAND2X1 U8371 ( .A(n7744), .B(n7906), .Y(n7995) );
  AND2X1 U8372 ( .A(n8064), .B(n8057), .Y(n8058) );
  NAND2X1 U8373 ( .A(n7908), .B(n7746), .Y(n8057) );
  NAND2X1 U8374 ( .A(n7586), .B(n8065), .Y(n8064) );
  NAND3X1 U8375 ( .A(n7997), .B(n8056), .C(n7569), .Y(n8065) );
  NAND2X1 U8376 ( .A(n8000), .B(G9), .Y(n8043) );
  AND3X1 U8377 ( .A(n8053), .B(n7997), .C(n7569), .Y(n8000) );
  NAND4X1 U8378 ( .A(n8066), .B(n8067), .C(n8068), .D(n8069), .Y(G896) );
  NOR3X1 U8379 ( .A(n8070), .B(n8071), .C(n8072), .Y(n8069) );
  NOR2X1 U8380 ( .A(n7483), .B(n8073), .Y(n8072) );
  NOR2X1 U8381 ( .A(n8074), .B(n7486), .Y(n8071) );
  NOR2X1 U8382 ( .A(n8075), .B(n7488), .Y(n8070) );
  NAND2X1 U8383 ( .A(G32), .B(n8076), .Y(n8068) );
  NAND2X1 U8384 ( .A(G21500), .B(n8077), .Y(n8067) );
  NAND2X1 U8385 ( .A(n8078), .B(G16), .Y(n8066) );
  NAND4X1 U8386 ( .A(n8079), .B(n8080), .C(n8081), .D(n8082), .Y(G895) );
  NOR3X1 U8387 ( .A(n8083), .B(n8084), .C(n8085), .Y(n8082) );
  NOR2X1 U8388 ( .A(n7499), .B(n8073), .Y(n8085) );
  NOR2X1 U8389 ( .A(n8074), .B(n7500), .Y(n8084) );
  NOR2X1 U8390 ( .A(n8075), .B(n7501), .Y(n8083) );
  NAND2X1 U8391 ( .A(G31), .B(n8076), .Y(n8081) );
  NAND2X1 U8392 ( .A(G21499), .B(n8077), .Y(n8080) );
  NAND2X1 U8393 ( .A(n8078), .B(G15), .Y(n8079) );
  NAND4X1 U8394 ( .A(n8086), .B(n8087), .C(n8088), .D(n8089), .Y(G894) );
  NOR3X1 U8395 ( .A(n8090), .B(n8091), .C(n8092), .Y(n8089) );
  NOR2X1 U8396 ( .A(n7509), .B(n8073), .Y(n8092) );
  NOR2X1 U8397 ( .A(n8074), .B(n7510), .Y(n8091) );
  NOR2X1 U8398 ( .A(n8075), .B(n7511), .Y(n8090) );
  NAND2X1 U8399 ( .A(G30), .B(n8076), .Y(n8088) );
  NAND2X1 U8400 ( .A(G21498), .B(n8077), .Y(n8087) );
  NAND2X1 U8401 ( .A(n8078), .B(G14), .Y(n8086) );
  NAND4X1 U8402 ( .A(n8093), .B(n8094), .C(n8095), .D(n8096), .Y(G893) );
  NOR3X1 U8403 ( .A(n8097), .B(n8098), .C(n8099), .Y(n8096) );
  NOR2X1 U8404 ( .A(n7519), .B(n8073), .Y(n8099) );
  NOR2X1 U8405 ( .A(n8074), .B(n7520), .Y(n8098) );
  NOR2X1 U8406 ( .A(n8075), .B(n7521), .Y(n8097) );
  NAND2X1 U8407 ( .A(G29), .B(n8076), .Y(n8095) );
  NAND2X1 U8408 ( .A(G21497), .B(n8077), .Y(n8094) );
  NAND2X1 U8409 ( .A(n8078), .B(G13), .Y(n8093) );
  NAND4X1 U8410 ( .A(n8100), .B(n8101), .C(n8102), .D(n8103), .Y(G892) );
  NOR3X1 U8411 ( .A(n8104), .B(n8105), .C(n8106), .Y(n8103) );
  NOR2X1 U8412 ( .A(n7529), .B(n8073), .Y(n8106) );
  NOR2X1 U8413 ( .A(n8074), .B(n7530), .Y(n8105) );
  NOR2X1 U8414 ( .A(n8075), .B(n7531), .Y(n8104) );
  NAND2X1 U8415 ( .A(G28), .B(n8076), .Y(n8102) );
  NAND2X1 U8416 ( .A(G21496), .B(n8077), .Y(n8101) );
  NAND2X1 U8417 ( .A(n8078), .B(G12), .Y(n8100) );
  NAND4X1 U8418 ( .A(n8107), .B(n8108), .C(n8109), .D(n8110), .Y(G891) );
  NOR3X1 U8419 ( .A(n8111), .B(n8112), .C(n8113), .Y(n8110) );
  NOR2X1 U8420 ( .A(n7539), .B(n8073), .Y(n8113) );
  NOR2X1 U8421 ( .A(n8074), .B(n7540), .Y(n8112) );
  NOR2X1 U8422 ( .A(n8075), .B(n7541), .Y(n8111) );
  NAND2X1 U8423 ( .A(G27), .B(n8076), .Y(n8109) );
  NAND2X1 U8424 ( .A(G21495), .B(n8077), .Y(n8108) );
  NAND2X1 U8425 ( .A(n8078), .B(G11), .Y(n8107) );
  NAND4X1 U8426 ( .A(n8114), .B(n8115), .C(n8116), .D(n8117), .Y(G890) );
  NOR3X1 U8427 ( .A(n8118), .B(n8119), .C(n8120), .Y(n8117) );
  NOR2X1 U8428 ( .A(n7549), .B(n8073), .Y(n8120) );
  NOR2X1 U8429 ( .A(n8074), .B(n7550), .Y(n8119) );
  NOR2X1 U8430 ( .A(n8075), .B(n7551), .Y(n8118) );
  NAND2X1 U8431 ( .A(G26), .B(n8076), .Y(n8116) );
  NAND2X1 U8432 ( .A(G21494), .B(n8077), .Y(n8115) );
  NAND2X1 U8433 ( .A(n8078), .B(G10), .Y(n8114) );
  NAND4X1 U8434 ( .A(n8121), .B(n8122), .C(n8123), .D(n8124), .Y(G889) );
  NOR3X1 U8435 ( .A(n8125), .B(n8126), .C(n8127), .Y(n8124) );
  NOR2X1 U8436 ( .A(n7559), .B(n8073), .Y(n8127) );
  NOR2X1 U8437 ( .A(n8074), .B(n7560), .Y(n8126) );
  AND2X1 U8438 ( .A(n8128), .B(n8129), .Y(n8074) );
  NAND2X1 U8439 ( .A(n8130), .B(n7564), .Y(n8129) );
  NAND2X1 U8440 ( .A(n8131), .B(G21426), .Y(n8128) );
  NOR2X1 U8441 ( .A(n8075), .B(n7566), .Y(n8125) );
  NAND2X1 U8442 ( .A(G25), .B(n8076), .Y(n8123) );
  NAND2X1 U8443 ( .A(n8132), .B(n8133), .Y(n8076) );
  NAND4X1 U8444 ( .A(n8130), .B(n7569), .C(n8075), .D(n8134), .Y(n8133) );
  INVX1 U8445 ( .A(n8135), .Y(n8130) );
  NAND2X1 U8446 ( .A(n8136), .B(n8137), .Y(n8132) );
  NAND2X1 U8447 ( .A(G21493), .B(n8077), .Y(n8122) );
  NAND2X1 U8448 ( .A(n8138), .B(n8139), .Y(n8077) );
  NAND3X1 U8449 ( .A(n8140), .B(n7577), .C(n8141), .Y(n8139) );
  NAND2X1 U8450 ( .A(n8137), .B(n7580), .Y(n8141) );
  NAND2X1 U8451 ( .A(n7579), .B(n8131), .Y(n8140) );
  NAND2X1 U8452 ( .A(n8136), .B(n8073), .Y(n8138) );
  AND2X1 U8453 ( .A(n8142), .B(n8135), .Y(n8136) );
  NAND2X1 U8454 ( .A(n7908), .B(n7826), .Y(n8135) );
  NOR2X1 U8455 ( .A(n7827), .B(n8143), .Y(n7908) );
  NAND2X1 U8456 ( .A(n7586), .B(n8144), .Y(n8142) );
  NAND3X1 U8457 ( .A(n8075), .B(n8134), .C(n7569), .Y(n8144) );
  NAND2X1 U8458 ( .A(n8078), .B(G9), .Y(n8121) );
  AND3X1 U8459 ( .A(n8131), .B(n8075), .C(n7569), .Y(n8078) );
  NAND4X1 U8460 ( .A(n8145), .B(n8146), .C(n8147), .D(n8148), .Y(G888) );
  NOR3X1 U8461 ( .A(n8149), .B(n8150), .C(n8151), .Y(n8148) );
  NOR2X1 U8462 ( .A(n7483), .B(n8152), .Y(n8151) );
  NOR2X1 U8463 ( .A(n8153), .B(n7486), .Y(n8150) );
  NOR2X1 U8464 ( .A(n8154), .B(n7488), .Y(n8149) );
  NAND2X1 U8465 ( .A(G32), .B(n8155), .Y(n8147) );
  NAND2X1 U8466 ( .A(G21492), .B(n8156), .Y(n8146) );
  NAND2X1 U8467 ( .A(n8157), .B(G16), .Y(n8145) );
  NAND4X1 U8468 ( .A(n8158), .B(n8159), .C(n8160), .D(n8161), .Y(G887) );
  NOR3X1 U8469 ( .A(n8162), .B(n8163), .C(n8164), .Y(n8161) );
  NOR2X1 U8470 ( .A(n7499), .B(n8152), .Y(n8164) );
  NOR2X1 U8471 ( .A(n8153), .B(n7500), .Y(n8163) );
  NOR2X1 U8472 ( .A(n8154), .B(n7501), .Y(n8162) );
  NAND2X1 U8473 ( .A(G31), .B(n8155), .Y(n8160) );
  NAND2X1 U8474 ( .A(G21491), .B(n8156), .Y(n8159) );
  NAND2X1 U8475 ( .A(n8157), .B(G15), .Y(n8158) );
  NAND4X1 U8476 ( .A(n8165), .B(n8166), .C(n8167), .D(n8168), .Y(G886) );
  NOR3X1 U8477 ( .A(n8169), .B(n8170), .C(n8171), .Y(n8168) );
  NOR2X1 U8478 ( .A(n7509), .B(n8152), .Y(n8171) );
  NOR2X1 U8479 ( .A(n8153), .B(n7510), .Y(n8170) );
  NOR2X1 U8480 ( .A(n8154), .B(n7511), .Y(n8169) );
  NAND2X1 U8481 ( .A(G30), .B(n8155), .Y(n8167) );
  NAND2X1 U8482 ( .A(G21490), .B(n8156), .Y(n8166) );
  NAND2X1 U8483 ( .A(n8157), .B(G14), .Y(n8165) );
  NAND4X1 U8484 ( .A(n8172), .B(n8173), .C(n8174), .D(n8175), .Y(G885) );
  NOR3X1 U8485 ( .A(n8176), .B(n8177), .C(n8178), .Y(n8175) );
  NOR2X1 U8486 ( .A(n7519), .B(n8152), .Y(n8178) );
  NOR2X1 U8487 ( .A(n8153), .B(n7520), .Y(n8177) );
  NOR2X1 U8488 ( .A(n8154), .B(n7521), .Y(n8176) );
  NAND2X1 U8489 ( .A(G29), .B(n8155), .Y(n8174) );
  NAND2X1 U8490 ( .A(G21489), .B(n8156), .Y(n8173) );
  NAND2X1 U8491 ( .A(n8157), .B(G13), .Y(n8172) );
  NAND4X1 U8492 ( .A(n8179), .B(n8180), .C(n8181), .D(n8182), .Y(G884) );
  NOR3X1 U8493 ( .A(n8183), .B(n8184), .C(n8185), .Y(n8182) );
  NOR2X1 U8494 ( .A(n7529), .B(n8152), .Y(n8185) );
  NOR2X1 U8495 ( .A(n8153), .B(n7530), .Y(n8184) );
  NOR2X1 U8496 ( .A(n8154), .B(n7531), .Y(n8183) );
  NAND2X1 U8497 ( .A(G28), .B(n8155), .Y(n8181) );
  NAND2X1 U8498 ( .A(G21488), .B(n8156), .Y(n8180) );
  NAND2X1 U8499 ( .A(n8157), .B(G12), .Y(n8179) );
  NAND4X1 U8500 ( .A(n8186), .B(n8187), .C(n8188), .D(n8189), .Y(G883) );
  NOR3X1 U8501 ( .A(n8190), .B(n8191), .C(n8192), .Y(n8189) );
  NOR2X1 U8502 ( .A(n7539), .B(n8152), .Y(n8192) );
  NOR2X1 U8503 ( .A(n8153), .B(n7540), .Y(n8191) );
  NOR2X1 U8504 ( .A(n8154), .B(n7541), .Y(n8190) );
  NAND2X1 U8505 ( .A(G27), .B(n8155), .Y(n8188) );
  NAND2X1 U8506 ( .A(G21487), .B(n8156), .Y(n8187) );
  NAND2X1 U8507 ( .A(n8157), .B(G11), .Y(n8186) );
  NAND4X1 U8508 ( .A(n8193), .B(n8194), .C(n8195), .D(n8196), .Y(G882) );
  NOR3X1 U8509 ( .A(n8197), .B(n8198), .C(n8199), .Y(n8196) );
  NOR2X1 U8510 ( .A(n7549), .B(n8152), .Y(n8199) );
  NOR2X1 U8511 ( .A(n8153), .B(n7550), .Y(n8198) );
  NOR2X1 U8512 ( .A(n8154), .B(n7551), .Y(n8197) );
  NAND2X1 U8513 ( .A(G26), .B(n8155), .Y(n8195) );
  NAND2X1 U8514 ( .A(G21486), .B(n8156), .Y(n8194) );
  NAND2X1 U8515 ( .A(n8157), .B(G10), .Y(n8193) );
  NAND4X1 U8516 ( .A(n8200), .B(n8201), .C(n8202), .D(n8203), .Y(G881) );
  NOR3X1 U8517 ( .A(n8204), .B(n8205), .C(n8206), .Y(n8203) );
  NOR2X1 U8518 ( .A(n7559), .B(n8152), .Y(n8206) );
  NOR2X1 U8519 ( .A(n8153), .B(n7560), .Y(n8205) );
  AND2X1 U8520 ( .A(n8207), .B(n8208), .Y(n8153) );
  NAND2X1 U8521 ( .A(n8209), .B(n7564), .Y(n8208) );
  NAND2X1 U8522 ( .A(n8210), .B(G21426), .Y(n8207) );
  NOR2X1 U8523 ( .A(n8154), .B(n7566), .Y(n8204) );
  NAND2X1 U8524 ( .A(G25), .B(n8155), .Y(n8202) );
  NAND2X1 U8525 ( .A(n8211), .B(n8212), .Y(n8155) );
  NAND4X1 U8526 ( .A(n8209), .B(n7569), .C(n8154), .D(n8213), .Y(n8212) );
  INVX1 U8527 ( .A(n8214), .Y(n8209) );
  NAND2X1 U8528 ( .A(n8215), .B(n8216), .Y(n8211) );
  NAND2X1 U8529 ( .A(G21485), .B(n8156), .Y(n8201) );
  NAND2X1 U8530 ( .A(n8217), .B(n8218), .Y(n8156) );
  NAND3X1 U8531 ( .A(n8219), .B(n7577), .C(n8220), .Y(n8218) );
  NAND2X1 U8532 ( .A(n7579), .B(n8210), .Y(n8220) );
  NAND2X1 U8533 ( .A(n8216), .B(n7580), .Y(n8219) );
  INVX1 U8534 ( .A(n8152), .Y(n8216) );
  NAND2X1 U8535 ( .A(n8215), .B(n8152), .Y(n8217) );
  NAND2X1 U8536 ( .A(n8221), .B(n7581), .Y(n8152) );
  AND2X1 U8537 ( .A(n8222), .B(n8214), .Y(n8215) );
  NAND2X1 U8538 ( .A(n8223), .B(n7584), .Y(n8214) );
  NAND2X1 U8539 ( .A(n7586), .B(n8224), .Y(n8222) );
  NAND3X1 U8540 ( .A(n8154), .B(n8213), .C(n7569), .Y(n8224) );
  NAND2X1 U8541 ( .A(n8157), .B(G9), .Y(n8200) );
  AND3X1 U8542 ( .A(n8210), .B(n8154), .C(n7569), .Y(n8157) );
  NAND4X1 U8543 ( .A(n8225), .B(n8226), .C(n8227), .D(n8228), .Y(G880) );
  NOR3X1 U8544 ( .A(n8229), .B(n8230), .C(n8231), .Y(n8228) );
  NOR2X1 U8545 ( .A(n7483), .B(n8232), .Y(n8231) );
  NOR2X1 U8546 ( .A(n8233), .B(n7486), .Y(n8230) );
  NOR2X1 U8547 ( .A(n8234), .B(n7488), .Y(n8229) );
  NAND2X1 U8548 ( .A(G32), .B(n8235), .Y(n8227) );
  NAND2X1 U8549 ( .A(G21484), .B(n8236), .Y(n8226) );
  NAND2X1 U8550 ( .A(n8237), .B(G16), .Y(n8225) );
  NAND4X1 U8551 ( .A(n8238), .B(n8239), .C(n8240), .D(n8241), .Y(G879) );
  NOR3X1 U8552 ( .A(n8242), .B(n8243), .C(n8244), .Y(n8241) );
  NOR2X1 U8553 ( .A(n7499), .B(n8232), .Y(n8244) );
  NOR2X1 U8554 ( .A(n8233), .B(n7500), .Y(n8243) );
  NOR2X1 U8555 ( .A(n8234), .B(n7501), .Y(n8242) );
  NAND2X1 U8556 ( .A(G31), .B(n8235), .Y(n8240) );
  NAND2X1 U8557 ( .A(G21483), .B(n8236), .Y(n8239) );
  NAND2X1 U8558 ( .A(n8237), .B(G15), .Y(n8238) );
  NAND4X1 U8559 ( .A(n8245), .B(n8246), .C(n8247), .D(n8248), .Y(G878) );
  NOR3X1 U8560 ( .A(n8249), .B(n8250), .C(n8251), .Y(n8248) );
  NOR2X1 U8561 ( .A(n7509), .B(n8232), .Y(n8251) );
  NOR2X1 U8562 ( .A(n8233), .B(n7510), .Y(n8250) );
  NOR2X1 U8563 ( .A(n8234), .B(n7511), .Y(n8249) );
  NAND2X1 U8564 ( .A(G30), .B(n8235), .Y(n8247) );
  NAND2X1 U8565 ( .A(G21482), .B(n8236), .Y(n8246) );
  NAND2X1 U8566 ( .A(n8237), .B(G14), .Y(n8245) );
  NAND4X1 U8567 ( .A(n8252), .B(n8253), .C(n8254), .D(n8255), .Y(G877) );
  NOR3X1 U8568 ( .A(n8256), .B(n8257), .C(n8258), .Y(n8255) );
  NOR2X1 U8569 ( .A(n7519), .B(n8232), .Y(n8258) );
  NOR2X1 U8570 ( .A(n8233), .B(n7520), .Y(n8257) );
  NOR2X1 U8571 ( .A(n8234), .B(n7521), .Y(n8256) );
  NAND2X1 U8572 ( .A(G29), .B(n8235), .Y(n8254) );
  NAND2X1 U8573 ( .A(G21481), .B(n8236), .Y(n8253) );
  NAND2X1 U8574 ( .A(n8237), .B(G13), .Y(n8252) );
  NAND4X1 U8575 ( .A(n8259), .B(n8260), .C(n8261), .D(n8262), .Y(G876) );
  NOR3X1 U8576 ( .A(n8263), .B(n8264), .C(n8265), .Y(n8262) );
  NOR2X1 U8577 ( .A(n7529), .B(n8232), .Y(n8265) );
  NOR2X1 U8578 ( .A(n8233), .B(n7530), .Y(n8264) );
  NOR2X1 U8579 ( .A(n8234), .B(n7531), .Y(n8263) );
  NAND2X1 U8580 ( .A(G28), .B(n8235), .Y(n8261) );
  NAND2X1 U8581 ( .A(G21480), .B(n8236), .Y(n8260) );
  NAND2X1 U8582 ( .A(n8237), .B(G12), .Y(n8259) );
  NAND4X1 U8583 ( .A(n8266), .B(n8267), .C(n8268), .D(n8269), .Y(G875) );
  NOR3X1 U8584 ( .A(n8270), .B(n8271), .C(n8272), .Y(n8269) );
  NOR2X1 U8585 ( .A(n7539), .B(n8232), .Y(n8272) );
  NOR2X1 U8586 ( .A(n8233), .B(n7540), .Y(n8271) );
  NOR2X1 U8587 ( .A(n8234), .B(n7541), .Y(n8270) );
  NAND2X1 U8588 ( .A(G27), .B(n8235), .Y(n8268) );
  NAND2X1 U8589 ( .A(G21479), .B(n8236), .Y(n8267) );
  NAND2X1 U8590 ( .A(n8237), .B(G11), .Y(n8266) );
  NAND4X1 U8591 ( .A(n8273), .B(n8274), .C(n8275), .D(n8276), .Y(G874) );
  NOR3X1 U8592 ( .A(n8277), .B(n8278), .C(n8279), .Y(n8276) );
  NOR2X1 U8593 ( .A(n7549), .B(n8232), .Y(n8279) );
  NOR2X1 U8594 ( .A(n8233), .B(n7550), .Y(n8278) );
  NOR2X1 U8595 ( .A(n8234), .B(n7551), .Y(n8277) );
  NAND2X1 U8596 ( .A(G26), .B(n8235), .Y(n8275) );
  NAND2X1 U8597 ( .A(G21478), .B(n8236), .Y(n8274) );
  NAND2X1 U8598 ( .A(n8237), .B(G10), .Y(n8273) );
  NAND4X1 U8599 ( .A(n8280), .B(n8281), .C(n8282), .D(n8283), .Y(G873) );
  NOR3X1 U8600 ( .A(n8284), .B(n8285), .C(n8286), .Y(n8283) );
  NOR2X1 U8601 ( .A(n7559), .B(n8232), .Y(n8286) );
  NOR2X1 U8602 ( .A(n8233), .B(n7560), .Y(n8285) );
  AND2X1 U8603 ( .A(n8287), .B(n8288), .Y(n8233) );
  NAND2X1 U8604 ( .A(n8289), .B(n7564), .Y(n8288) );
  NAND2X1 U8605 ( .A(n8290), .B(G21426), .Y(n8287) );
  NOR2X1 U8606 ( .A(n8234), .B(n7566), .Y(n8284) );
  NAND2X1 U8607 ( .A(G25), .B(n8235), .Y(n8282) );
  NAND2X1 U8608 ( .A(n8291), .B(n8292), .Y(n8235) );
  NAND4X1 U8609 ( .A(n8289), .B(n7569), .C(n8234), .D(n8293), .Y(n8292) );
  INVX1 U8610 ( .A(n8294), .Y(n8289) );
  NAND2X1 U8611 ( .A(n8295), .B(n8296), .Y(n8291) );
  NAND2X1 U8612 ( .A(G21477), .B(n8236), .Y(n8281) );
  NAND2X1 U8613 ( .A(n8297), .B(n8298), .Y(n8236) );
  NAND3X1 U8614 ( .A(n8299), .B(n7577), .C(n8300), .Y(n8298) );
  NAND2X1 U8615 ( .A(n7579), .B(n8290), .Y(n8300) );
  NAND2X1 U8616 ( .A(n8296), .B(n7580), .Y(n8299) );
  INVX1 U8617 ( .A(n8232), .Y(n8296) );
  NAND2X1 U8618 ( .A(n8295), .B(n8232), .Y(n8297) );
  NAND2X1 U8619 ( .A(n8221), .B(n7664), .Y(n8232) );
  AND2X1 U8620 ( .A(n8301), .B(n8294), .Y(n8295) );
  NAND2X1 U8621 ( .A(n8223), .B(n7666), .Y(n8294) );
  NAND2X1 U8622 ( .A(n7586), .B(n8302), .Y(n8301) );
  NAND3X1 U8623 ( .A(n8234), .B(n8293), .C(n7569), .Y(n8302) );
  NAND2X1 U8624 ( .A(n8237), .B(G9), .Y(n8280) );
  AND3X1 U8625 ( .A(n8290), .B(n8234), .C(n7569), .Y(n8237) );
  NAND4X1 U8626 ( .A(n8303), .B(n8304), .C(n8305), .D(n8306), .Y(G872) );
  NOR3X1 U8627 ( .A(n8307), .B(n8308), .C(n8309), .Y(n8306) );
  NOR2X1 U8628 ( .A(n7483), .B(n8310), .Y(n8309) );
  NOR2X1 U8629 ( .A(n8311), .B(n7486), .Y(n8308) );
  NOR2X1 U8630 ( .A(n8312), .B(n7488), .Y(n8307) );
  NAND2X1 U8631 ( .A(G32), .B(n8313), .Y(n8305) );
  NAND2X1 U8632 ( .A(G21476), .B(n8314), .Y(n8304) );
  NAND2X1 U8633 ( .A(n8315), .B(G16), .Y(n8303) );
  NAND4X1 U8634 ( .A(n8316), .B(n8317), .C(n8318), .D(n8319), .Y(G871) );
  NOR3X1 U8635 ( .A(n8320), .B(n8321), .C(n8322), .Y(n8319) );
  NOR2X1 U8636 ( .A(n7499), .B(n8310), .Y(n8322) );
  NOR2X1 U8637 ( .A(n8311), .B(n7500), .Y(n8321) );
  NOR2X1 U8638 ( .A(n8312), .B(n7501), .Y(n8320) );
  NAND2X1 U8639 ( .A(G31), .B(n8313), .Y(n8318) );
  NAND2X1 U8640 ( .A(G21475), .B(n8314), .Y(n8317) );
  NAND2X1 U8641 ( .A(n8315), .B(G15), .Y(n8316) );
  NAND4X1 U8642 ( .A(n8323), .B(n8324), .C(n8325), .D(n8326), .Y(G870) );
  NOR3X1 U8643 ( .A(n8327), .B(n8328), .C(n8329), .Y(n8326) );
  NOR2X1 U8644 ( .A(n7509), .B(n8310), .Y(n8329) );
  NOR2X1 U8645 ( .A(n8311), .B(n7510), .Y(n8328) );
  NOR2X1 U8646 ( .A(n8312), .B(n7511), .Y(n8327) );
  NAND2X1 U8647 ( .A(G30), .B(n8313), .Y(n8325) );
  NAND2X1 U8648 ( .A(G21474), .B(n8314), .Y(n8324) );
  NAND2X1 U8649 ( .A(n8315), .B(G14), .Y(n8323) );
  NAND4X1 U8650 ( .A(n8330), .B(n8331), .C(n8332), .D(n8333), .Y(G869) );
  NOR3X1 U8651 ( .A(n8334), .B(n8335), .C(n8336), .Y(n8333) );
  NOR2X1 U8652 ( .A(n7519), .B(n8310), .Y(n8336) );
  NOR2X1 U8653 ( .A(n8311), .B(n7520), .Y(n8335) );
  NOR2X1 U8654 ( .A(n8312), .B(n7521), .Y(n8334) );
  NAND2X1 U8655 ( .A(G29), .B(n8313), .Y(n8332) );
  NAND2X1 U8656 ( .A(G21473), .B(n8314), .Y(n8331) );
  NAND2X1 U8657 ( .A(n8315), .B(G13), .Y(n8330) );
  NAND4X1 U8658 ( .A(n8337), .B(n8338), .C(n8339), .D(n8340), .Y(G868) );
  NOR3X1 U8659 ( .A(n8341), .B(n8342), .C(n8343), .Y(n8340) );
  NOR2X1 U8660 ( .A(n7529), .B(n8310), .Y(n8343) );
  NOR2X1 U8661 ( .A(n8311), .B(n7530), .Y(n8342) );
  NOR2X1 U8662 ( .A(n8312), .B(n7531), .Y(n8341) );
  NAND2X1 U8663 ( .A(G28), .B(n8313), .Y(n8339) );
  NAND2X1 U8664 ( .A(G21472), .B(n8314), .Y(n8338) );
  NAND2X1 U8665 ( .A(n8315), .B(G12), .Y(n8337) );
  NAND4X1 U8666 ( .A(n8344), .B(n8345), .C(n8346), .D(n8347), .Y(G867) );
  NOR3X1 U8667 ( .A(n8348), .B(n8349), .C(n8350), .Y(n8347) );
  NOR2X1 U8668 ( .A(n7539), .B(n8310), .Y(n8350) );
  NOR2X1 U8669 ( .A(n8311), .B(n7540), .Y(n8349) );
  NOR2X1 U8670 ( .A(n8312), .B(n7541), .Y(n8348) );
  NAND2X1 U8671 ( .A(G27), .B(n8313), .Y(n8346) );
  NAND2X1 U8672 ( .A(G21471), .B(n8314), .Y(n8345) );
  NAND2X1 U8673 ( .A(n8315), .B(G11), .Y(n8344) );
  NAND4X1 U8674 ( .A(n8351), .B(n8352), .C(n8353), .D(n8354), .Y(G866) );
  NOR3X1 U8675 ( .A(n8355), .B(n8356), .C(n8357), .Y(n8354) );
  NOR2X1 U8676 ( .A(n7549), .B(n8310), .Y(n8357) );
  NOR2X1 U8677 ( .A(n8311), .B(n7550), .Y(n8356) );
  NOR2X1 U8678 ( .A(n8312), .B(n7551), .Y(n8355) );
  NAND2X1 U8679 ( .A(G26), .B(n8313), .Y(n8353) );
  NAND2X1 U8680 ( .A(G21470), .B(n8314), .Y(n8352) );
  NAND2X1 U8681 ( .A(n8315), .B(G10), .Y(n8351) );
  NAND4X1 U8682 ( .A(n8358), .B(n8359), .C(n8360), .D(n8361), .Y(G865) );
  NOR3X1 U8683 ( .A(n8362), .B(n8363), .C(n8364), .Y(n8361) );
  NOR2X1 U8684 ( .A(n7559), .B(n8310), .Y(n8364) );
  NOR2X1 U8685 ( .A(n8311), .B(n7560), .Y(n8363) );
  AND2X1 U8686 ( .A(n8365), .B(n8366), .Y(n8311) );
  NAND2X1 U8687 ( .A(n8367), .B(n7564), .Y(n8366) );
  NAND2X1 U8688 ( .A(n8368), .B(G21426), .Y(n8365) );
  NOR2X1 U8689 ( .A(n8312), .B(n7566), .Y(n8362) );
  NAND2X1 U8690 ( .A(G25), .B(n8313), .Y(n8360) );
  NAND2X1 U8691 ( .A(n8369), .B(n8370), .Y(n8313) );
  NAND4X1 U8692 ( .A(n8367), .B(n7569), .C(n8312), .D(n8371), .Y(n8370) );
  INVX1 U8693 ( .A(n8372), .Y(n8367) );
  NAND2X1 U8694 ( .A(n8373), .B(n8374), .Y(n8369) );
  NAND2X1 U8695 ( .A(G21469), .B(n8314), .Y(n8359) );
  NAND2X1 U8696 ( .A(n8375), .B(n8376), .Y(n8314) );
  NAND3X1 U8697 ( .A(n8377), .B(n7577), .C(n8378), .Y(n8376) );
  NAND2X1 U8698 ( .A(n7579), .B(n8368), .Y(n8378) );
  NAND2X1 U8699 ( .A(n8374), .B(n7580), .Y(n8377) );
  INVX1 U8700 ( .A(n8310), .Y(n8374) );
  NAND2X1 U8701 ( .A(n8373), .B(n8310), .Y(n8375) );
  NAND2X1 U8702 ( .A(n8221), .B(n7744), .Y(n8310) );
  AND2X1 U8703 ( .A(n8379), .B(n8372), .Y(n8373) );
  NAND2X1 U8704 ( .A(n8223), .B(n7746), .Y(n8372) );
  NAND2X1 U8705 ( .A(n7586), .B(n8380), .Y(n8379) );
  NAND3X1 U8706 ( .A(n8312), .B(n8371), .C(n7569), .Y(n8380) );
  NAND2X1 U8707 ( .A(n8315), .B(G9), .Y(n8358) );
  AND3X1 U8708 ( .A(n8368), .B(n8312), .C(n7569), .Y(n8315) );
  NAND4X1 U8709 ( .A(n8381), .B(n8382), .C(n8383), .D(n8384), .Y(G864) );
  NOR3X1 U8710 ( .A(n8385), .B(n8386), .C(n8387), .Y(n8384) );
  NOR2X1 U8711 ( .A(n7483), .B(n8388), .Y(n8387) );
  NOR2X1 U8712 ( .A(n8389), .B(n7486), .Y(n8386) );
  NOR2X1 U8713 ( .A(n8390), .B(n7488), .Y(n8385) );
  NAND2X1 U8714 ( .A(G32), .B(n8391), .Y(n8383) );
  NAND2X1 U8715 ( .A(G21468), .B(n8392), .Y(n8382) );
  NAND2X1 U8716 ( .A(n8393), .B(G16), .Y(n8381) );
  NAND4X1 U8717 ( .A(n8394), .B(n8395), .C(n8396), .D(n8397), .Y(G863) );
  NOR3X1 U8718 ( .A(n8398), .B(n8399), .C(n8400), .Y(n8397) );
  NOR2X1 U8719 ( .A(n7499), .B(n8388), .Y(n8400) );
  NOR2X1 U8720 ( .A(n8389), .B(n7500), .Y(n8399) );
  NOR2X1 U8721 ( .A(n8390), .B(n7501), .Y(n8398) );
  NAND2X1 U8722 ( .A(G31), .B(n8391), .Y(n8396) );
  NAND2X1 U8723 ( .A(G21467), .B(n8392), .Y(n8395) );
  NAND2X1 U8724 ( .A(n8393), .B(G15), .Y(n8394) );
  NAND4X1 U8725 ( .A(n8401), .B(n8402), .C(n8403), .D(n8404), .Y(G862) );
  NOR3X1 U8726 ( .A(n8405), .B(n8406), .C(n8407), .Y(n8404) );
  NOR2X1 U8727 ( .A(n7509), .B(n8388), .Y(n8407) );
  NOR2X1 U8728 ( .A(n8389), .B(n7510), .Y(n8406) );
  NOR2X1 U8729 ( .A(n8390), .B(n7511), .Y(n8405) );
  NAND2X1 U8730 ( .A(G30), .B(n8391), .Y(n8403) );
  NAND2X1 U8731 ( .A(G21466), .B(n8392), .Y(n8402) );
  NAND2X1 U8732 ( .A(n8393), .B(G14), .Y(n8401) );
  NAND4X1 U8733 ( .A(n8408), .B(n8409), .C(n8410), .D(n8411), .Y(G861) );
  NOR3X1 U8734 ( .A(n8412), .B(n8413), .C(n8414), .Y(n8411) );
  NOR2X1 U8735 ( .A(n7519), .B(n8388), .Y(n8414) );
  NOR2X1 U8736 ( .A(n8389), .B(n7520), .Y(n8413) );
  NOR2X1 U8737 ( .A(n8390), .B(n7521), .Y(n8412) );
  NAND2X1 U8738 ( .A(G29), .B(n8391), .Y(n8410) );
  NAND2X1 U8739 ( .A(G21465), .B(n8392), .Y(n8409) );
  NAND2X1 U8740 ( .A(n8393), .B(G13), .Y(n8408) );
  NAND4X1 U8741 ( .A(n8415), .B(n8416), .C(n8417), .D(n8418), .Y(G860) );
  NOR3X1 U8742 ( .A(n8419), .B(n8420), .C(n8421), .Y(n8418) );
  NOR2X1 U8743 ( .A(n7529), .B(n8388), .Y(n8421) );
  NOR2X1 U8744 ( .A(n8389), .B(n7530), .Y(n8420) );
  NOR2X1 U8745 ( .A(n8390), .B(n7531), .Y(n8419) );
  NAND2X1 U8746 ( .A(G28), .B(n8391), .Y(n8417) );
  NAND2X1 U8747 ( .A(G21464), .B(n8392), .Y(n8416) );
  NAND2X1 U8748 ( .A(n8393), .B(G12), .Y(n8415) );
  NAND4X1 U8749 ( .A(n8422), .B(n8423), .C(n8424), .D(n8425), .Y(G859) );
  NOR3X1 U8750 ( .A(n8426), .B(n8427), .C(n8428), .Y(n8425) );
  NOR2X1 U8751 ( .A(n7539), .B(n8388), .Y(n8428) );
  NOR2X1 U8752 ( .A(n8389), .B(n7540), .Y(n8427) );
  NOR2X1 U8753 ( .A(n8390), .B(n7541), .Y(n8426) );
  NAND2X1 U8754 ( .A(G27), .B(n8391), .Y(n8424) );
  NAND2X1 U8755 ( .A(G21463), .B(n8392), .Y(n8423) );
  NAND2X1 U8756 ( .A(n8393), .B(G11), .Y(n8422) );
  NAND4X1 U8757 ( .A(n8429), .B(n8430), .C(n8431), .D(n8432), .Y(G858) );
  NOR3X1 U8758 ( .A(n8433), .B(n8434), .C(n8435), .Y(n8432) );
  NOR2X1 U8759 ( .A(n7549), .B(n8388), .Y(n8435) );
  NOR2X1 U8760 ( .A(n8389), .B(n7550), .Y(n8434) );
  NOR2X1 U8761 ( .A(n8390), .B(n7551), .Y(n8433) );
  NAND2X1 U8762 ( .A(G26), .B(n8391), .Y(n8431) );
  NAND2X1 U8763 ( .A(G21462), .B(n8392), .Y(n8430) );
  NAND2X1 U8764 ( .A(n8393), .B(G10), .Y(n8429) );
  NAND4X1 U8765 ( .A(n8436), .B(n8437), .C(n8438), .D(n8439), .Y(G857) );
  NOR3X1 U8766 ( .A(n8440), .B(n8441), .C(n8442), .Y(n8439) );
  NOR2X1 U8767 ( .A(n7559), .B(n8388), .Y(n8442) );
  NOR2X1 U8768 ( .A(n8389), .B(n7560), .Y(n8441) );
  AND2X1 U8769 ( .A(n8443), .B(n8444), .Y(n8389) );
  NAND2X1 U8770 ( .A(n8445), .B(n7564), .Y(n8444) );
  NAND2X1 U8771 ( .A(n8446), .B(G21426), .Y(n8443) );
  NOR2X1 U8772 ( .A(n8390), .B(n7566), .Y(n8440) );
  NAND2X1 U8773 ( .A(G25), .B(n8391), .Y(n8438) );
  NAND2X1 U8774 ( .A(n8447), .B(n8448), .Y(n8391) );
  NAND4X1 U8775 ( .A(n8445), .B(n7569), .C(n8390), .D(n8449), .Y(n8448) );
  INVX1 U8776 ( .A(n8450), .Y(n8445) );
  NAND2X1 U8777 ( .A(n8451), .B(n8452), .Y(n8447) );
  NAND2X1 U8778 ( .A(G21461), .B(n8392), .Y(n8437) );
  NAND2X1 U8779 ( .A(n8453), .B(n8454), .Y(n8392) );
  NAND3X1 U8780 ( .A(n8455), .B(n7577), .C(n8456), .Y(n8454) );
  NAND2X1 U8781 ( .A(n7579), .B(n8446), .Y(n8456) );
  NAND2X1 U8782 ( .A(n8452), .B(n7580), .Y(n8455) );
  INVX1 U8783 ( .A(n8388), .Y(n8452) );
  NAND2X1 U8784 ( .A(n8451), .B(n8388), .Y(n8453) );
  NAND2X1 U8785 ( .A(n8221), .B(n7824), .Y(n8388) );
  AND2X1 U8786 ( .A(n8457), .B(n8450), .Y(n8451) );
  NAND2X1 U8787 ( .A(n8223), .B(n7826), .Y(n8450) );
  NOR2X1 U8788 ( .A(n7828), .B(n8458), .Y(n8223) );
  NAND2X1 U8789 ( .A(n7586), .B(n8459), .Y(n8457) );
  NAND3X1 U8790 ( .A(n8390), .B(n8449), .C(n7569), .Y(n8459) );
  NAND2X1 U8791 ( .A(n8393), .B(G9), .Y(n8436) );
  AND3X1 U8792 ( .A(n8446), .B(n8390), .C(n7569), .Y(n8393) );
  NAND4X1 U8793 ( .A(n8460), .B(n8461), .C(n8462), .D(n8463), .Y(G856) );
  NOR3X1 U8794 ( .A(n8464), .B(n8465), .C(n8466), .Y(n8463) );
  NOR2X1 U8795 ( .A(n7483), .B(n8467), .Y(n8466) );
  NOR2X1 U8796 ( .A(n8468), .B(n7486), .Y(n8465) );
  NOR2X1 U8797 ( .A(n8469), .B(n7488), .Y(n8464) );
  NAND2X1 U8798 ( .A(G32), .B(n8470), .Y(n8462) );
  NAND2X1 U8799 ( .A(G21460), .B(n8471), .Y(n8461) );
  NAND2X1 U8800 ( .A(n8472), .B(G16), .Y(n8460) );
  NAND4X1 U8801 ( .A(n8473), .B(n8474), .C(n8475), .D(n8476), .Y(G855) );
  NOR3X1 U8802 ( .A(n8477), .B(n8478), .C(n8479), .Y(n8476) );
  NOR2X1 U8803 ( .A(n7499), .B(n8467), .Y(n8479) );
  NOR2X1 U8804 ( .A(n8468), .B(n7500), .Y(n8478) );
  NOR2X1 U8805 ( .A(n8469), .B(n7501), .Y(n8477) );
  NAND2X1 U8806 ( .A(G31), .B(n8470), .Y(n8475) );
  NAND2X1 U8807 ( .A(G21459), .B(n8471), .Y(n8474) );
  NAND2X1 U8808 ( .A(n8472), .B(G15), .Y(n8473) );
  NAND4X1 U8809 ( .A(n8480), .B(n8481), .C(n8482), .D(n8483), .Y(G854) );
  NOR3X1 U8810 ( .A(n8484), .B(n8485), .C(n8486), .Y(n8483) );
  NOR2X1 U8811 ( .A(n7509), .B(n8467), .Y(n8486) );
  NOR2X1 U8812 ( .A(n8468), .B(n7510), .Y(n8485) );
  NOR2X1 U8813 ( .A(n8469), .B(n7511), .Y(n8484) );
  NAND2X1 U8814 ( .A(G30), .B(n8470), .Y(n8482) );
  NAND2X1 U8815 ( .A(G21458), .B(n8471), .Y(n8481) );
  NAND2X1 U8816 ( .A(n8472), .B(G14), .Y(n8480) );
  NAND4X1 U8817 ( .A(n8487), .B(n8488), .C(n8489), .D(n8490), .Y(G853) );
  NOR3X1 U8818 ( .A(n8491), .B(n8492), .C(n8493), .Y(n8490) );
  NOR2X1 U8819 ( .A(n7519), .B(n8467), .Y(n8493) );
  NOR2X1 U8820 ( .A(n8468), .B(n7520), .Y(n8492) );
  NOR2X1 U8821 ( .A(n8469), .B(n7521), .Y(n8491) );
  NAND2X1 U8822 ( .A(G29), .B(n8470), .Y(n8489) );
  NAND2X1 U8823 ( .A(G21457), .B(n8471), .Y(n8488) );
  NAND2X1 U8824 ( .A(n8472), .B(G13), .Y(n8487) );
  NAND4X1 U8825 ( .A(n8494), .B(n8495), .C(n8496), .D(n8497), .Y(G852) );
  NOR3X1 U8826 ( .A(n8498), .B(n8499), .C(n8500), .Y(n8497) );
  NOR2X1 U8827 ( .A(n7529), .B(n8467), .Y(n8500) );
  NOR2X1 U8828 ( .A(n8468), .B(n7530), .Y(n8499) );
  NOR2X1 U8829 ( .A(n8469), .B(n7531), .Y(n8498) );
  NAND2X1 U8830 ( .A(G28), .B(n8470), .Y(n8496) );
  NAND2X1 U8831 ( .A(G21456), .B(n8471), .Y(n8495) );
  NAND2X1 U8832 ( .A(n8472), .B(G12), .Y(n8494) );
  NAND4X1 U8833 ( .A(n8501), .B(n8502), .C(n8503), .D(n8504), .Y(G851) );
  NOR3X1 U8834 ( .A(n8505), .B(n8506), .C(n8507), .Y(n8504) );
  NOR2X1 U8835 ( .A(n7539), .B(n8467), .Y(n8507) );
  NOR2X1 U8836 ( .A(n8468), .B(n7540), .Y(n8506) );
  NOR2X1 U8837 ( .A(n8469), .B(n7541), .Y(n8505) );
  NAND2X1 U8838 ( .A(G27), .B(n8470), .Y(n8503) );
  NAND2X1 U8839 ( .A(G21455), .B(n8471), .Y(n8502) );
  NAND2X1 U8840 ( .A(n8472), .B(G11), .Y(n8501) );
  NAND4X1 U8841 ( .A(n8508), .B(n8509), .C(n8510), .D(n8511), .Y(G850) );
  NOR3X1 U8842 ( .A(n8512), .B(n8513), .C(n8514), .Y(n8511) );
  NOR2X1 U8843 ( .A(n7549), .B(n8467), .Y(n8514) );
  NOR2X1 U8844 ( .A(n8468), .B(n7550), .Y(n8513) );
  NOR2X1 U8845 ( .A(n8469), .B(n7551), .Y(n8512) );
  NAND2X1 U8846 ( .A(G26), .B(n8470), .Y(n8510) );
  NAND2X1 U8847 ( .A(G21454), .B(n8471), .Y(n8509) );
  NAND2X1 U8848 ( .A(n8472), .B(G10), .Y(n8508) );
  NAND4X1 U8849 ( .A(n8515), .B(n8516), .C(n8517), .D(n8518), .Y(G849) );
  NOR3X1 U8850 ( .A(n8519), .B(n8520), .C(n8521), .Y(n8518) );
  NOR2X1 U8851 ( .A(n7559), .B(n8467), .Y(n8521) );
  NOR2X1 U8852 ( .A(n8468), .B(n7560), .Y(n8520) );
  AND2X1 U8853 ( .A(n8522), .B(n8523), .Y(n8468) );
  NAND2X1 U8854 ( .A(n8524), .B(n7564), .Y(n8523) );
  NAND2X1 U8855 ( .A(n8525), .B(G21426), .Y(n8522) );
  NOR2X1 U8856 ( .A(n8469), .B(n7566), .Y(n8519) );
  NAND2X1 U8857 ( .A(G25), .B(n8470), .Y(n8517) );
  NAND2X1 U8858 ( .A(n8526), .B(n8527), .Y(n8470) );
  NAND4X1 U8859 ( .A(n8524), .B(n7569), .C(n8469), .D(n8528), .Y(n8527) );
  INVX1 U8860 ( .A(n8529), .Y(n8524) );
  NAND2X1 U8861 ( .A(n8530), .B(n8531), .Y(n8526) );
  NAND2X1 U8862 ( .A(G21453), .B(n8471), .Y(n8516) );
  NAND2X1 U8863 ( .A(n8532), .B(n8533), .Y(n8471) );
  NAND3X1 U8864 ( .A(n8534), .B(n7577), .C(n8535), .Y(n8533) );
  NAND2X1 U8865 ( .A(n7579), .B(n8525), .Y(n8535) );
  NAND2X1 U8866 ( .A(n8531), .B(n7580), .Y(n8534) );
  INVX1 U8867 ( .A(n8467), .Y(n8531) );
  NAND2X1 U8868 ( .A(n8530), .B(n8467), .Y(n8532) );
  NAND2X1 U8869 ( .A(n8536), .B(n7581), .Y(n8467) );
  NOR2X1 U8870 ( .A(G21566), .B(G21565), .Y(n7581) );
  AND2X1 U8871 ( .A(n8537), .B(n8529), .Y(n8530) );
  NAND2X1 U8872 ( .A(n8538), .B(n7584), .Y(n8529) );
  NOR2X1 U8873 ( .A(n8539), .B(n8540), .Y(n7584) );
  NAND2X1 U8874 ( .A(n7586), .B(n8541), .Y(n8537) );
  NAND3X1 U8875 ( .A(n8469), .B(n8528), .C(n7569), .Y(n8541) );
  NAND2X1 U8876 ( .A(n8472), .B(G9), .Y(n8515) );
  AND3X1 U8877 ( .A(n8525), .B(n8469), .C(n7569), .Y(n8472) );
  NAND4X1 U8878 ( .A(n8542), .B(n8543), .C(n8544), .D(n8545), .Y(G848) );
  NOR3X1 U8879 ( .A(n8546), .B(n8547), .C(n8548), .Y(n8545) );
  NOR2X1 U8880 ( .A(n7483), .B(n8549), .Y(n8548) );
  NOR2X1 U8881 ( .A(n8550), .B(n7486), .Y(n8547) );
  NOR2X1 U8882 ( .A(n8551), .B(n7488), .Y(n8546) );
  NAND2X1 U8883 ( .A(G32), .B(n8552), .Y(n8544) );
  NAND2X1 U8884 ( .A(G21452), .B(n8553), .Y(n8543) );
  NAND2X1 U8885 ( .A(n8554), .B(G16), .Y(n8542) );
  NAND4X1 U8886 ( .A(n8555), .B(n8556), .C(n8557), .D(n8558), .Y(G847) );
  NOR3X1 U8887 ( .A(n8559), .B(n8560), .C(n8561), .Y(n8558) );
  NOR2X1 U8888 ( .A(n7499), .B(n8549), .Y(n8561) );
  NOR2X1 U8889 ( .A(n8550), .B(n7500), .Y(n8560) );
  NOR2X1 U8890 ( .A(n8551), .B(n7501), .Y(n8559) );
  NAND2X1 U8891 ( .A(G31), .B(n8552), .Y(n8557) );
  NAND2X1 U8892 ( .A(G21451), .B(n8553), .Y(n8556) );
  NAND2X1 U8893 ( .A(n8554), .B(G15), .Y(n8555) );
  NAND4X1 U8894 ( .A(n8562), .B(n8563), .C(n8564), .D(n8565), .Y(G846) );
  NOR3X1 U8895 ( .A(n8566), .B(n8567), .C(n8568), .Y(n8565) );
  NOR2X1 U8896 ( .A(n7509), .B(n8549), .Y(n8568) );
  NOR2X1 U8897 ( .A(n8550), .B(n7510), .Y(n8567) );
  NOR2X1 U8898 ( .A(n8551), .B(n7511), .Y(n8566) );
  NAND2X1 U8899 ( .A(G30), .B(n8552), .Y(n8564) );
  NAND2X1 U8900 ( .A(G21450), .B(n8553), .Y(n8563) );
  NAND2X1 U8901 ( .A(n8554), .B(G14), .Y(n8562) );
  NAND4X1 U8902 ( .A(n8569), .B(n8570), .C(n8571), .D(n8572), .Y(G845) );
  NOR3X1 U8903 ( .A(n8573), .B(n8574), .C(n8575), .Y(n8572) );
  NOR2X1 U8904 ( .A(n7519), .B(n8549), .Y(n8575) );
  NOR2X1 U8905 ( .A(n8550), .B(n7520), .Y(n8574) );
  NOR2X1 U8906 ( .A(n8551), .B(n7521), .Y(n8573) );
  NAND2X1 U8907 ( .A(G29), .B(n8552), .Y(n8571) );
  NAND2X1 U8908 ( .A(G21449), .B(n8553), .Y(n8570) );
  NAND2X1 U8909 ( .A(n8554), .B(G13), .Y(n8569) );
  NAND4X1 U8910 ( .A(n8576), .B(n8577), .C(n8578), .D(n8579), .Y(G844) );
  NOR3X1 U8911 ( .A(n8580), .B(n8581), .C(n8582), .Y(n8579) );
  NOR2X1 U8912 ( .A(n7529), .B(n8549), .Y(n8582) );
  NOR2X1 U8913 ( .A(n8550), .B(n7530), .Y(n8581) );
  NOR2X1 U8914 ( .A(n8551), .B(n7531), .Y(n8580) );
  NAND2X1 U8915 ( .A(G28), .B(n8552), .Y(n8578) );
  NAND2X1 U8916 ( .A(G21448), .B(n8553), .Y(n8577) );
  NAND2X1 U8917 ( .A(n8554), .B(G12), .Y(n8576) );
  NAND4X1 U8918 ( .A(n8583), .B(n8584), .C(n8585), .D(n8586), .Y(G843) );
  NOR3X1 U8919 ( .A(n8587), .B(n8588), .C(n8589), .Y(n8586) );
  NOR2X1 U8920 ( .A(n7539), .B(n8549), .Y(n8589) );
  NOR2X1 U8921 ( .A(n8550), .B(n7540), .Y(n8588) );
  NOR2X1 U8922 ( .A(n8551), .B(n7541), .Y(n8587) );
  NAND2X1 U8923 ( .A(G27), .B(n8552), .Y(n8585) );
  NAND2X1 U8924 ( .A(G21447), .B(n8553), .Y(n8584) );
  NAND2X1 U8925 ( .A(n8554), .B(G11), .Y(n8583) );
  NAND4X1 U8926 ( .A(n8590), .B(n8591), .C(n8592), .D(n8593), .Y(G842) );
  NOR3X1 U8927 ( .A(n8594), .B(n8595), .C(n8596), .Y(n8593) );
  NOR2X1 U8928 ( .A(n7549), .B(n8549), .Y(n8596) );
  NOR2X1 U8929 ( .A(n8550), .B(n7550), .Y(n8595) );
  NOR2X1 U8930 ( .A(n8551), .B(n7551), .Y(n8594) );
  NAND2X1 U8931 ( .A(G26), .B(n8552), .Y(n8592) );
  NAND2X1 U8932 ( .A(G21446), .B(n8553), .Y(n8591) );
  NAND2X1 U8933 ( .A(n8554), .B(G10), .Y(n8590) );
  NAND4X1 U8934 ( .A(n8597), .B(n8598), .C(n8599), .D(n8600), .Y(G841) );
  NOR3X1 U8935 ( .A(n8601), .B(n8602), .C(n8603), .Y(n8600) );
  NOR2X1 U8936 ( .A(n7559), .B(n8549), .Y(n8603) );
  NOR2X1 U8937 ( .A(n8550), .B(n7560), .Y(n8602) );
  AND2X1 U8938 ( .A(n8604), .B(n8605), .Y(n8550) );
  NAND2X1 U8939 ( .A(n8606), .B(n7564), .Y(n8605) );
  NAND2X1 U8940 ( .A(n8607), .B(G21426), .Y(n8604) );
  NOR2X1 U8941 ( .A(n8551), .B(n7566), .Y(n8601) );
  NAND2X1 U8942 ( .A(G25), .B(n8552), .Y(n8599) );
  NAND2X1 U8943 ( .A(n8608), .B(n8609), .Y(n8552) );
  NAND4X1 U8944 ( .A(n8606), .B(n7569), .C(n8551), .D(n8610), .Y(n8609) );
  INVX1 U8945 ( .A(n8611), .Y(n8606) );
  NAND2X1 U8946 ( .A(n8612), .B(n8613), .Y(n8608) );
  NAND2X1 U8947 ( .A(G21445), .B(n8553), .Y(n8598) );
  NAND2X1 U8948 ( .A(n8614), .B(n8615), .Y(n8553) );
  NAND3X1 U8949 ( .A(n8616), .B(n7577), .C(n8617), .Y(n8615) );
  NAND2X1 U8950 ( .A(n7579), .B(n8607), .Y(n8617) );
  NAND2X1 U8951 ( .A(n8613), .B(n7580), .Y(n8616) );
  INVX1 U8952 ( .A(n8549), .Y(n8613) );
  NAND2X1 U8953 ( .A(n8612), .B(n8549), .Y(n8614) );
  NAND2X1 U8954 ( .A(n8536), .B(n7664), .Y(n8549) );
  AND2X1 U8955 ( .A(n8618), .B(n8611), .Y(n8612) );
  NAND2X1 U8956 ( .A(n8538), .B(n7666), .Y(n8611) );
  NOR2X1 U8957 ( .A(n8539), .B(G21566), .Y(n7666) );
  NAND2X1 U8958 ( .A(n7586), .B(n8619), .Y(n8618) );
  NAND3X1 U8959 ( .A(n8551), .B(n8610), .C(n7569), .Y(n8619) );
  NAND2X1 U8960 ( .A(n8554), .B(G9), .Y(n8597) );
  AND3X1 U8961 ( .A(n8607), .B(n8551), .C(n7569), .Y(n8554) );
  NAND4X1 U8962 ( .A(n8620), .B(n8621), .C(n8622), .D(n8623), .Y(G840) );
  NOR3X1 U8963 ( .A(n8624), .B(n8625), .C(n8626), .Y(n8623) );
  NOR2X1 U8964 ( .A(n7483), .B(n8627), .Y(n8626) );
  NOR2X1 U8965 ( .A(n8628), .B(n7486), .Y(n8625) );
  NOR2X1 U8966 ( .A(n8629), .B(n7488), .Y(n8624) );
  NAND2X1 U8967 ( .A(G32), .B(n8630), .Y(n8622) );
  NAND2X1 U8968 ( .A(G21444), .B(n8631), .Y(n8621) );
  NAND2X1 U8969 ( .A(n8632), .B(G16), .Y(n8620) );
  NAND4X1 U8970 ( .A(n8633), .B(n8634), .C(n8635), .D(n8636), .Y(G839) );
  NOR3X1 U8971 ( .A(n8637), .B(n8638), .C(n8639), .Y(n8636) );
  NOR2X1 U8972 ( .A(n7499), .B(n8627), .Y(n8639) );
  NOR2X1 U8973 ( .A(n8628), .B(n7500), .Y(n8638) );
  NOR2X1 U8974 ( .A(n8629), .B(n7501), .Y(n8637) );
  NAND2X1 U8975 ( .A(G31), .B(n8630), .Y(n8635) );
  NAND2X1 U8976 ( .A(G21443), .B(n8631), .Y(n8634) );
  NAND2X1 U8977 ( .A(n8632), .B(G15), .Y(n8633) );
  NAND4X1 U8978 ( .A(n8640), .B(n8641), .C(n8642), .D(n8643), .Y(G838) );
  NOR3X1 U8979 ( .A(n8644), .B(n8645), .C(n8646), .Y(n8643) );
  NOR2X1 U8980 ( .A(n7509), .B(n8627), .Y(n8646) );
  NOR2X1 U8981 ( .A(n8628), .B(n7510), .Y(n8645) );
  NOR2X1 U8982 ( .A(n8629), .B(n7511), .Y(n8644) );
  NAND2X1 U8983 ( .A(G30), .B(n8630), .Y(n8642) );
  NAND2X1 U8984 ( .A(G21442), .B(n8631), .Y(n8641) );
  NAND2X1 U8985 ( .A(n8632), .B(G14), .Y(n8640) );
  NAND4X1 U8986 ( .A(n8647), .B(n8648), .C(n8649), .D(n8650), .Y(G837) );
  NOR3X1 U8987 ( .A(n8651), .B(n8652), .C(n8653), .Y(n8650) );
  NOR2X1 U8988 ( .A(n7519), .B(n8627), .Y(n8653) );
  NOR2X1 U8989 ( .A(n8628), .B(n7520), .Y(n8652) );
  NOR2X1 U8990 ( .A(n8629), .B(n7521), .Y(n8651) );
  NAND2X1 U8991 ( .A(G29), .B(n8630), .Y(n8649) );
  NAND2X1 U8992 ( .A(G21441), .B(n8631), .Y(n8648) );
  NAND2X1 U8993 ( .A(n8632), .B(G13), .Y(n8647) );
  NAND4X1 U8994 ( .A(n8654), .B(n8655), .C(n8656), .D(n8657), .Y(G836) );
  NOR3X1 U8995 ( .A(n8658), .B(n8659), .C(n8660), .Y(n8657) );
  NOR2X1 U8996 ( .A(n7529), .B(n8627), .Y(n8660) );
  NOR2X1 U8997 ( .A(n8628), .B(n7530), .Y(n8659) );
  NOR2X1 U8998 ( .A(n8629), .B(n7531), .Y(n8658) );
  NAND2X1 U8999 ( .A(G28), .B(n8630), .Y(n8656) );
  NAND2X1 U9000 ( .A(G21440), .B(n8631), .Y(n8655) );
  NAND2X1 U9001 ( .A(n8632), .B(G12), .Y(n8654) );
  NAND4X1 U9002 ( .A(n8661), .B(n8662), .C(n8663), .D(n8664), .Y(G835) );
  NOR3X1 U9003 ( .A(n8665), .B(n8666), .C(n8667), .Y(n8664) );
  NOR2X1 U9004 ( .A(n7539), .B(n8627), .Y(n8667) );
  NOR2X1 U9005 ( .A(n8628), .B(n7540), .Y(n8666) );
  NOR2X1 U9006 ( .A(n8629), .B(n7541), .Y(n8665) );
  NAND2X1 U9007 ( .A(G27), .B(n8630), .Y(n8663) );
  NAND2X1 U9008 ( .A(G21439), .B(n8631), .Y(n8662) );
  NAND2X1 U9009 ( .A(n8632), .B(G11), .Y(n8661) );
  NAND4X1 U9010 ( .A(n8668), .B(n8669), .C(n8670), .D(n8671), .Y(G834) );
  NOR3X1 U9011 ( .A(n8672), .B(n8673), .C(n8674), .Y(n8671) );
  NOR2X1 U9012 ( .A(n7549), .B(n8627), .Y(n8674) );
  NOR2X1 U9013 ( .A(n8628), .B(n7550), .Y(n8673) );
  NOR2X1 U9014 ( .A(n8629), .B(n7551), .Y(n8672) );
  NAND2X1 U9015 ( .A(G26), .B(n8630), .Y(n8670) );
  NAND2X1 U9016 ( .A(G21438), .B(n8631), .Y(n8669) );
  NAND2X1 U9017 ( .A(n8632), .B(G10), .Y(n8668) );
  NAND4X1 U9018 ( .A(n8675), .B(n8676), .C(n8677), .D(n8678), .Y(G833) );
  NOR3X1 U9019 ( .A(n8679), .B(n8680), .C(n8681), .Y(n8678) );
  NOR2X1 U9020 ( .A(n7559), .B(n8627), .Y(n8681) );
  NOR2X1 U9021 ( .A(n8628), .B(n7560), .Y(n8680) );
  AND2X1 U9022 ( .A(n8682), .B(n8683), .Y(n8628) );
  NAND2X1 U9023 ( .A(n8684), .B(n7564), .Y(n8683) );
  NAND2X1 U9024 ( .A(n8685), .B(G21426), .Y(n8682) );
  NOR2X1 U9025 ( .A(n8629), .B(n7566), .Y(n8679) );
  NAND2X1 U9026 ( .A(G25), .B(n8630), .Y(n8677) );
  NAND2X1 U9027 ( .A(n8686), .B(n8687), .Y(n8630) );
  NAND4X1 U9028 ( .A(n8684), .B(n7569), .C(n8629), .D(n8688), .Y(n8687) );
  INVX1 U9029 ( .A(n8689), .Y(n8684) );
  NAND2X1 U9030 ( .A(n8690), .B(n8691), .Y(n8686) );
  NAND2X1 U9031 ( .A(G21437), .B(n8631), .Y(n8676) );
  NAND2X1 U9032 ( .A(n8692), .B(n8693), .Y(n8631) );
  NAND3X1 U9033 ( .A(n8694), .B(n7577), .C(n8695), .Y(n8693) );
  NAND2X1 U9034 ( .A(n7579), .B(n8685), .Y(n8695) );
  NAND2X1 U9035 ( .A(n8691), .B(n7580), .Y(n8694) );
  INVX1 U9036 ( .A(n8627), .Y(n8691) );
  NAND2X1 U9037 ( .A(n8690), .B(n8627), .Y(n8692) );
  NAND2X1 U9038 ( .A(n8536), .B(n7744), .Y(n8627) );
  AND2X1 U9039 ( .A(n8696), .B(n8689), .Y(n8690) );
  NAND2X1 U9040 ( .A(n8538), .B(n7746), .Y(n8689) );
  NOR2X1 U9041 ( .A(n8540), .B(n8697), .Y(n7746) );
  NAND2X1 U9042 ( .A(n7586), .B(n8698), .Y(n8696) );
  NAND3X1 U9043 ( .A(n8629), .B(n8688), .C(n7569), .Y(n8698) );
  NAND2X1 U9044 ( .A(n8632), .B(G9), .Y(n8675) );
  AND3X1 U9045 ( .A(n8685), .B(n8629), .C(n7569), .Y(n8632) );
  NAND4X1 U9046 ( .A(n8699), .B(n8700), .C(n8701), .D(n8702), .Y(G832) );
  NOR3X1 U9047 ( .A(n8703), .B(n8704), .C(n8705), .Y(n8702) );
  NOR2X1 U9048 ( .A(n8706), .B(n7488), .Y(n8705) );
  NAND2X1 U9049 ( .A(G8), .B(n7569), .Y(n7488) );
  NOR2X1 U9050 ( .A(n7483), .B(n8707), .Y(n8704) );
  AND2X1 U9051 ( .A(n8708), .B(n8709), .Y(n7483) );
  OR2X1 U9052 ( .A(n7486), .B(n7430), .Y(n8709) );
  NAND2X1 U9053 ( .A(n8710), .B(n8711), .Y(n8708) );
  NOR2X1 U9054 ( .A(n8712), .B(n7486), .Y(n8703) );
  NAND2X1 U9055 ( .A(G32), .B(n7580), .Y(n7486) );
  NAND2X1 U9056 ( .A(G32), .B(n8713), .Y(n8701) );
  NAND2X1 U9057 ( .A(G21436), .B(n8714), .Y(n8700) );
  NAND2X1 U9058 ( .A(n8715), .B(G16), .Y(n8699) );
  NAND4X1 U9059 ( .A(n8716), .B(n8717), .C(n8718), .D(n8719), .Y(G831) );
  NOR3X1 U9060 ( .A(n8720), .B(n8721), .C(n8722), .Y(n8719) );
  NOR2X1 U9061 ( .A(n8706), .B(n7501), .Y(n8722) );
  NAND2X1 U9062 ( .A(G7), .B(n7569), .Y(n7501) );
  NOR2X1 U9063 ( .A(n7499), .B(n8707), .Y(n8721) );
  AND2X1 U9064 ( .A(n8723), .B(n8724), .Y(n7499) );
  OR2X1 U9065 ( .A(n7500), .B(n7430), .Y(n8724) );
  NAND2X1 U9066 ( .A(n8710), .B(n7444), .Y(n8723) );
  NOR2X1 U9067 ( .A(n8712), .B(n7500), .Y(n8720) );
  NAND2X1 U9068 ( .A(G31), .B(n7580), .Y(n7500) );
  NAND2X1 U9069 ( .A(G31), .B(n8713), .Y(n8718) );
  NAND2X1 U9070 ( .A(G21435), .B(n8714), .Y(n8717) );
  NAND2X1 U9071 ( .A(n8715), .B(G15), .Y(n8716) );
  NAND4X1 U9072 ( .A(n8725), .B(n8726), .C(n8727), .D(n8728), .Y(G830) );
  NOR3X1 U9073 ( .A(n8729), .B(n8730), .C(n8731), .Y(n8728) );
  NOR2X1 U9074 ( .A(n8706), .B(n7511), .Y(n8731) );
  NAND2X1 U9075 ( .A(G6), .B(n7569), .Y(n7511) );
  NOR2X1 U9076 ( .A(n7509), .B(n8707), .Y(n8730) );
  AND2X1 U9077 ( .A(n8732), .B(n8733), .Y(n7509) );
  OR2X1 U9078 ( .A(n7510), .B(n7430), .Y(n8733) );
  NAND2X1 U9079 ( .A(n8710), .B(n7456), .Y(n8732) );
  NOR2X1 U9080 ( .A(n8712), .B(n7510), .Y(n8729) );
  NAND2X1 U9081 ( .A(G30), .B(n7580), .Y(n7510) );
  NAND2X1 U9082 ( .A(G30), .B(n8713), .Y(n8727) );
  NAND2X1 U9083 ( .A(G21434), .B(n8714), .Y(n8726) );
  NAND2X1 U9084 ( .A(n8715), .B(G14), .Y(n8725) );
  NAND4X1 U9085 ( .A(n8734), .B(n8735), .C(n8736), .D(n8737), .Y(G829) );
  NOR3X1 U9086 ( .A(n8738), .B(n8739), .C(n8740), .Y(n8737) );
  NOR2X1 U9087 ( .A(n8706), .B(n7521), .Y(n8740) );
  NAND2X1 U9088 ( .A(G5), .B(n7569), .Y(n7521) );
  NOR2X1 U9089 ( .A(n7519), .B(n8707), .Y(n8739) );
  AND2X1 U9090 ( .A(n8741), .B(n8742), .Y(n7519) );
  OR2X1 U9091 ( .A(n7520), .B(n7430), .Y(n8742) );
  NAND2X1 U9092 ( .A(n8710), .B(n8743), .Y(n8741) );
  NOR2X1 U9093 ( .A(n8712), .B(n7520), .Y(n8738) );
  NAND2X1 U9094 ( .A(G29), .B(n7580), .Y(n7520) );
  NAND2X1 U9095 ( .A(G29), .B(n8713), .Y(n8736) );
  NAND2X1 U9096 ( .A(G21433), .B(n8714), .Y(n8735) );
  NAND2X1 U9097 ( .A(n8715), .B(G13), .Y(n8734) );
  NAND4X1 U9098 ( .A(n8744), .B(n8745), .C(n8746), .D(n8747), .Y(G828) );
  NOR3X1 U9099 ( .A(n8748), .B(n8749), .C(n8750), .Y(n8747) );
  NOR2X1 U9100 ( .A(n8706), .B(n7531), .Y(n8750) );
  NAND2X1 U9101 ( .A(G4), .B(n7569), .Y(n7531) );
  NOR2X1 U9102 ( .A(n7529), .B(n8707), .Y(n8749) );
  AND2X1 U9103 ( .A(n8751), .B(n8752), .Y(n7529) );
  OR2X1 U9104 ( .A(n7530), .B(n7430), .Y(n8752) );
  NAND2X1 U9105 ( .A(n8710), .B(n7458), .Y(n8751) );
  NOR2X1 U9106 ( .A(n8712), .B(n7530), .Y(n8748) );
  NAND2X1 U9107 ( .A(G28), .B(n7580), .Y(n7530) );
  NAND2X1 U9108 ( .A(G28), .B(n8713), .Y(n8746) );
  NAND2X1 U9109 ( .A(G21432), .B(n8714), .Y(n8745) );
  NAND2X1 U9110 ( .A(n8715), .B(G12), .Y(n8744) );
  NAND4X1 U9111 ( .A(n8753), .B(n8754), .C(n8755), .D(n8756), .Y(G827) );
  NOR3X1 U9112 ( .A(n8757), .B(n8758), .C(n8759), .Y(n8756) );
  NOR2X1 U9113 ( .A(n8706), .B(n7541), .Y(n8759) );
  NAND2X1 U9114 ( .A(G3), .B(n7569), .Y(n7541) );
  NOR2X1 U9115 ( .A(n7539), .B(n8707), .Y(n8758) );
  AND2X1 U9116 ( .A(n8760), .B(n8761), .Y(n7539) );
  OR2X1 U9117 ( .A(n7540), .B(n7430), .Y(n8761) );
  NAND2X1 U9118 ( .A(n8710), .B(n8762), .Y(n8760) );
  NOR2X1 U9119 ( .A(n8712), .B(n7540), .Y(n8757) );
  NAND2X1 U9120 ( .A(G27), .B(n7580), .Y(n7540) );
  NAND2X1 U9121 ( .A(G27), .B(n8713), .Y(n8755) );
  NAND2X1 U9122 ( .A(G21431), .B(n8714), .Y(n8754) );
  NAND2X1 U9123 ( .A(n8715), .B(G11), .Y(n8753) );
  NAND4X1 U9124 ( .A(n8763), .B(n8764), .C(n8765), .D(n8766), .Y(G826) );
  NOR3X1 U9125 ( .A(n8767), .B(n8768), .C(n8769), .Y(n8766) );
  NOR2X1 U9126 ( .A(n8706), .B(n7551), .Y(n8769) );
  NAND2X1 U9127 ( .A(G2), .B(n7569), .Y(n7551) );
  NOR2X1 U9128 ( .A(n7549), .B(n8707), .Y(n8768) );
  AND2X1 U9129 ( .A(n8770), .B(n8771), .Y(n7549) );
  OR2X1 U9130 ( .A(n7550), .B(n7430), .Y(n8771) );
  NAND2X1 U9131 ( .A(n8710), .B(n8772), .Y(n8770) );
  NOR2X1 U9132 ( .A(n8712), .B(n7550), .Y(n8767) );
  NAND2X1 U9133 ( .A(G26), .B(n7580), .Y(n7550) );
  NAND2X1 U9134 ( .A(G26), .B(n8713), .Y(n8765) );
  NAND2X1 U9135 ( .A(G21430), .B(n8714), .Y(n8764) );
  NAND2X1 U9136 ( .A(n8715), .B(G10), .Y(n8763) );
  NAND4X1 U9137 ( .A(n8773), .B(n8774), .C(n8775), .D(n8776), .Y(G825) );
  NOR3X1 U9138 ( .A(n8777), .B(n8778), .C(n8779), .Y(n8776) );
  NOR2X1 U9139 ( .A(n8706), .B(n7566), .Y(n8779) );
  NAND2X1 U9140 ( .A(G1), .B(n7569), .Y(n7566) );
  NOR2X1 U9141 ( .A(n7559), .B(n8707), .Y(n8778) );
  AND2X1 U9142 ( .A(n8780), .B(n8781), .Y(n7559) );
  NAND2X1 U9143 ( .A(n8710), .B(n8782), .Y(n8781) );
  NOR2X1 U9144 ( .A(n8783), .B(n8784), .Y(n8710) );
  OR2X1 U9145 ( .A(n7560), .B(n7430), .Y(n8780) );
  NOR2X1 U9146 ( .A(n8712), .B(n7560), .Y(n8777) );
  NAND2X1 U9147 ( .A(G25), .B(n7580), .Y(n7560) );
  AND2X1 U9148 ( .A(n8785), .B(n8786), .Y(n8712) );
  NAND2X1 U9149 ( .A(n8787), .B(n7564), .Y(n8786) );
  NAND2X1 U9150 ( .A(n8788), .B(G21426), .Y(n8785) );
  NAND2X1 U9151 ( .A(G25), .B(n8713), .Y(n8775) );
  NAND2X1 U9152 ( .A(n8789), .B(n8790), .Y(n8713) );
  NAND3X1 U9153 ( .A(n7569), .B(n8706), .C(n8787), .Y(n8790) );
  INVX1 U9154 ( .A(n8791), .Y(n8787) );
  NAND2X1 U9155 ( .A(n8792), .B(n8793), .Y(n8789) );
  NAND2X1 U9156 ( .A(G21429), .B(n8714), .Y(n8774) );
  NAND2X1 U9157 ( .A(n8794), .B(n8795), .Y(n8714) );
  NAND3X1 U9158 ( .A(n8796), .B(n7577), .C(n8797), .Y(n8795) );
  NAND2X1 U9159 ( .A(n8793), .B(n7580), .Y(n8797) );
  INVX1 U9160 ( .A(n8707), .Y(n8793) );
  NAND2X1 U9161 ( .A(n7579), .B(n7430), .Y(n7577) );
  NAND2X1 U9162 ( .A(n7579), .B(n8788), .Y(n8796) );
  NOR2X1 U9163 ( .A(n8784), .B(n8798), .Y(n7579) );
  NAND2X1 U9164 ( .A(n8792), .B(n8707), .Y(n8794) );
  NAND2X1 U9165 ( .A(n8536), .B(n7824), .Y(n8707) );
  NOR2X1 U9166 ( .A(n8799), .B(n8800), .Y(n8536) );
  AND2X1 U9167 ( .A(n8801), .B(n8791), .Y(n8792) );
  NAND2X1 U9168 ( .A(n8538), .B(n7826), .Y(n8791) );
  NOR2X1 U9169 ( .A(G21566), .B(n8697), .Y(n7826) );
  NOR2X1 U9170 ( .A(n8143), .B(n8458), .Y(n8538) );
  INVX1 U9171 ( .A(n7828), .Y(n8143) );
  NAND2X1 U9172 ( .A(n7586), .B(n8802), .Y(n8801) );
  NAND3X1 U9173 ( .A(n8706), .B(n8803), .C(n7569), .Y(n8802) );
  NAND2X1 U9174 ( .A(n7564), .B(n7580), .Y(n7586) );
  NAND2X1 U9175 ( .A(n8715), .B(G9), .Y(n8773) );
  AND2X1 U9176 ( .A(n7569), .B(n8788), .Y(n8715) );
  NAND4X1 U9177 ( .A(n8805), .B(n8806), .C(n8807), .D(n8808), .Y(G824) );
  NAND2X1 U9178 ( .A(n8809), .B(G21428), .Y(n8808) );
  NAND2X1 U9179 ( .A(n8810), .B(n8811), .Y(n8807) );
  NAND3X1 U9180 ( .A(n8812), .B(n8813), .C(n8814), .Y(n8810) );
  NAND2X1 U9181 ( .A(n8815), .B(n7457), .Y(n8814) );
  NAND2X1 U9182 ( .A(n8816), .B(n8817), .Y(n8813) );
  NAND3X1 U9183 ( .A(G21425), .B(n7457), .C(n8798), .Y(n8816) );
  NAND2X1 U9184 ( .A(n8818), .B(n8819), .Y(n8812) );
  NAND3X1 U9185 ( .A(n8820), .B(n8821), .C(n8822), .Y(G823) );
  NAND2X1 U9186 ( .A(G21427), .B(n8823), .Y(n8822) );
  NAND2X1 U9187 ( .A(n8811), .B(n8806), .Y(n8823) );
  NAND3X1 U9188 ( .A(G21428), .B(n7430), .C(G35), .Y(n8806) );
  NAND2X1 U9189 ( .A(n8824), .B(n8811), .Y(n8820) );
  NAND2X1 U9190 ( .A(n8825), .B(n8826), .Y(n8824) );
  NAND3X1 U9191 ( .A(G21428), .B(n7445), .C(n8827), .Y(n8826) );
  INVX1 U9192 ( .A(n7433), .Y(n8825) );
  NAND4X1 U9193 ( .A(n8828), .B(n8829), .C(n8830), .D(n8831), .Y(G822) );
  OR2X1 U9194 ( .A(n8804), .B(G21428), .Y(n8831) );
  NAND4X1 U9195 ( .A(n7430), .B(n7445), .C(G21427), .D(G21428), .Y(n8830) );
  NAND3X1 U9196 ( .A(n8832), .B(n8833), .C(n8834), .Y(G821) );
  NAND2X1 U9197 ( .A(n8809), .B(G21425), .Y(n8834) );
  INVX1 U9198 ( .A(n8811), .Y(n8809) );
  NAND4X1 U9199 ( .A(n8835), .B(n8836), .C(n8837), .D(n8838), .Y(n8811) );
  NAND2X1 U9200 ( .A(n8817), .B(n7445), .Y(n8838) );
  NAND2X1 U9201 ( .A(G21428), .B(n8839), .Y(n8837) );
  OR2X1 U9202 ( .A(n8819), .B(G21427), .Y(n8839) );
  NAND4X1 U9203 ( .A(n8840), .B(n7427), .C(n8841), .D(n8842), .Y(n8819) );
  NOR4X1 U9204 ( .A(n8843), .B(n8844), .C(n8845), .D(n8846), .Y(n8842) );
  NOR2X1 U9205 ( .A(n7424), .B(n8847), .Y(n8846) );
  NOR2X1 U9206 ( .A(n8848), .B(n8849), .Y(n8845) );
  NOR2X1 U9207 ( .A(n7441), .B(n7429), .Y(n8844) );
  NOR2X1 U9208 ( .A(n8850), .B(n8851), .Y(n8843) );
  NOR2X1 U9209 ( .A(n8852), .B(n8853), .Y(n8841) );
  NOR2X1 U9210 ( .A(n8854), .B(n7457), .Y(n8853) );
  NOR3X1 U9211 ( .A(n8855), .B(n8856), .C(n8857), .Y(n8854) );
  NOR2X1 U9212 ( .A(n8711), .B(n8858), .Y(n8857) );
  NOR2X1 U9213 ( .A(n8859), .B(n8860), .Y(n8852) );
  NOR2X1 U9214 ( .A(G21795), .B(G21796), .Y(n8859) );
  INVX1 U9215 ( .A(n8861), .Y(n7427) );
  NAND3X1 U9216 ( .A(n8862), .B(n7474), .C(n8863), .Y(n8840) );
  NAND2X1 U9217 ( .A(G21563), .B(n8851), .Y(n8863) );
  NAND3X1 U9218 ( .A(n8864), .B(n8865), .C(n8866), .Y(n8862) );
  OR2X1 U9219 ( .A(n8851), .B(G21563), .Y(n8866) );
  NAND2X1 U9220 ( .A(n8867), .B(n8868), .Y(n8851) );
  NAND2X1 U9221 ( .A(n8869), .B(n8870), .Y(n8868) );
  OR2X1 U9222 ( .A(n8871), .B(n8869), .Y(n8867) );
  NAND3X1 U9223 ( .A(n8872), .B(n8873), .C(n8874), .Y(n8865) );
  NAND2X1 U9224 ( .A(G21564), .B(n8850), .Y(n8874) );
  NAND2X1 U9225 ( .A(n8875), .B(n8849), .Y(n8873) );
  NAND2X1 U9226 ( .A(n8876), .B(n8877), .Y(n8875) );
  NAND2X1 U9227 ( .A(n8878), .B(n8879), .Y(n8877) );
  NAND2X1 U9228 ( .A(n8880), .B(n8881), .Y(n8879) );
  NAND2X1 U9229 ( .A(n8882), .B(G21566), .Y(n8881) );
  INVX1 U9230 ( .A(n8883), .Y(n8878) );
  NAND2X1 U9231 ( .A(n8882), .B(n7824), .Y(n8876) );
  INVX1 U9232 ( .A(n8884), .Y(n8882) );
  NAND2X1 U9233 ( .A(n8869), .B(n8885), .Y(n8872) );
  NAND3X1 U9234 ( .A(n8886), .B(n8887), .C(n8888), .Y(n8885) );
  NAND2X1 U9235 ( .A(G21566), .B(n8889), .Y(n8888) );
  NAND2X1 U9236 ( .A(n7824), .B(n8890), .Y(n8886) );
  OR2X1 U9237 ( .A(n8850), .B(G21564), .Y(n8864) );
  NAND2X1 U9238 ( .A(n8891), .B(n8892), .Y(n8850) );
  NAND2X1 U9239 ( .A(n8869), .B(n8893), .Y(n8892) );
  OR2X1 U9240 ( .A(n8894), .B(n8869), .Y(n8891) );
  INVX1 U9241 ( .A(n8849), .Y(n8869) );
  NAND2X1 U9242 ( .A(n8895), .B(n8856), .Y(n8836) );
  NAND2X1 U9243 ( .A(n8896), .B(n8897), .Y(n8835) );
  INVX1 U9244 ( .A(n8898), .Y(n8833) );
  NOR2X1 U9245 ( .A(n8899), .B(n8900), .Y(G820) );
  NOR2X1 U9246 ( .A(n8899), .B(n8901), .Y(G819) );
  NOR2X1 U9247 ( .A(n8899), .B(n8902), .Y(G818) );
  NOR2X1 U9248 ( .A(n8899), .B(n8903), .Y(G817) );
  NOR2X1 U9249 ( .A(n8899), .B(n8904), .Y(G816) );
  NOR2X1 U9250 ( .A(n8899), .B(n8905), .Y(G815) );
  NOR2X1 U9251 ( .A(n8899), .B(n8906), .Y(G814) );
  NOR2X1 U9252 ( .A(n8899), .B(n8907), .Y(G813) );
  NOR2X1 U9253 ( .A(n8899), .B(n8908), .Y(G812) );
  NOR2X1 U9254 ( .A(n8899), .B(n8909), .Y(G811) );
  NOR2X1 U9255 ( .A(n8899), .B(n8910), .Y(G810) );
  NOR2X1 U9256 ( .A(n8899), .B(n8911), .Y(G809) );
  NOR2X1 U9257 ( .A(n8899), .B(n8912), .Y(G808) );
  NOR2X1 U9258 ( .A(n8899), .B(n8913), .Y(G807) );
  NOR2X1 U9259 ( .A(n8899), .B(n8914), .Y(G806) );
  NOR2X1 U9260 ( .A(n8899), .B(n8915), .Y(G805) );
  AND2X1 U9261 ( .A(n8916), .B(G21408), .Y(G804) );
  AND2X1 U9262 ( .A(n8916), .B(G21407), .Y(G803) );
  AND2X1 U9263 ( .A(n8916), .B(G21406), .Y(G802) );
  AND2X1 U9264 ( .A(n8916), .B(G21405), .Y(G801) );
  AND2X1 U9265 ( .A(n8916), .B(G21404), .Y(G800) );
  AND2X1 U9266 ( .A(n8916), .B(G21403), .Y(G799) );
  AND2X1 U9267 ( .A(n8916), .B(G21402), .Y(G798) );
  AND2X1 U9268 ( .A(n8916), .B(G21401), .Y(G797) );
  NOR2X1 U9269 ( .A(n8899), .B(n8917), .Y(G796) );
  NOR2X1 U9270 ( .A(n8899), .B(n8918), .Y(G795) );
  NOR2X1 U9271 ( .A(n8899), .B(n8919), .Y(G794) );
  NOR2X1 U9272 ( .A(n8899), .B(n8920), .Y(G793) );
  AND2X1 U9273 ( .A(n8916), .B(G21396), .Y(G792) );
  AND2X1 U9274 ( .A(n8916), .B(G21395), .Y(G791) );
  NAND3X1 U9275 ( .A(n8921), .B(n8922), .C(n8923), .Y(G790) );
  NOR3X1 U9276 ( .A(n8924), .B(n8925), .C(n8926), .Y(n8923) );
  NOR3X1 U9277 ( .A(n8927), .B(G21392), .C(G21391), .Y(n8926) );
  NOR2X1 U9278 ( .A(G21798), .B(n8928), .Y(n8924) );
  NAND2X1 U9279 ( .A(n8929), .B(n8930), .Y(n8922) );
  NAND2X1 U9280 ( .A(n8931), .B(n8932), .Y(n8921) );
  NAND4X1 U9281 ( .A(n8933), .B(n8934), .C(n8935), .D(n8936), .Y(G789) );
  NAND2X1 U9282 ( .A(n8937), .B(n8938), .Y(n8936) );
  NAND2X1 U9283 ( .A(n8939), .B(n8940), .Y(n8937) );
  NAND3X1 U9284 ( .A(G21392), .B(n8941), .C(G21798), .Y(n8940) );
  NAND4X1 U9285 ( .A(n8942), .B(n8939), .C(n8943), .D(G21391), .Y(n8935) );
  NAND2X1 U9286 ( .A(n8944), .B(n8945), .Y(n8943) );
  NAND2X1 U9287 ( .A(n8931), .B(n7445), .Y(n8942) );
  INVX1 U9288 ( .A(n8941), .Y(n8931) );
  NAND2X1 U9289 ( .A(G36), .B(G21390), .Y(n8941) );
  INVX1 U9290 ( .A(n8946), .Y(n8934) );
  NAND2X1 U9291 ( .A(n8947), .B(G35), .Y(n8933) );
  NAND4X1 U9292 ( .A(n8948), .B(n8949), .C(n8950), .D(n8951), .Y(G787) );
  INVX1 U9293 ( .A(n8928), .Y(n8951) );
  NAND3X1 U9294 ( .A(G21392), .B(n8952), .C(G36), .Y(n8950) );
  NAND3X1 U9295 ( .A(n8953), .B(n8954), .C(n8955), .Y(n8952) );
  NAND2X1 U9296 ( .A(n8938), .B(n8945), .Y(n8954) );
  NAND3X1 U9297 ( .A(G35), .B(n8927), .C(G21391), .Y(n8953) );
  NAND3X1 U9298 ( .A(G21390), .B(n8930), .C(G21391), .Y(n8949) );
  INVX1 U9299 ( .A(n8944), .Y(n8930) );
  NOR2X1 U9300 ( .A(G36), .B(G35), .Y(n8944) );
  NAND2X1 U9301 ( .A(n8956), .B(n8927), .Y(n8948) );
  INVX1 U9302 ( .A(G33), .Y(n8927) );
  NAND2X1 U9303 ( .A(n8939), .B(n8957), .Y(n8956) );
  OR3X1 U9304 ( .A(n8945), .B(n7445), .C(n8958), .Y(n8957) );
  NAND2X1 U9305 ( .A(G21390), .B(n8959), .Y(n8939) );
  NAND3X1 U9306 ( .A(n8960), .B(n8961), .C(n8962), .Y(G786) );
  NAND2X1 U9307 ( .A(G21389), .B(n8932), .Y(n8962) );
  NAND2X1 U9308 ( .A(n8928), .B(G21759), .Y(n8961) );
  NAND2X1 U9309 ( .A(n8946), .B(G21760), .Y(n8960) );
  NAND3X1 U9310 ( .A(n8963), .B(n8964), .C(n8965), .Y(G785) );
  NAND2X1 U9311 ( .A(G21388), .B(n8932), .Y(n8965) );
  NAND2X1 U9312 ( .A(n8928), .B(G21760), .Y(n8964) );
  NAND2X1 U9313 ( .A(n8946), .B(G21761), .Y(n8963) );
  NAND3X1 U9314 ( .A(n8966), .B(n8967), .C(n8968), .Y(G784) );
  NAND2X1 U9315 ( .A(G21387), .B(n8932), .Y(n8968) );
  NAND2X1 U9316 ( .A(n8928), .B(G21761), .Y(n8967) );
  NAND2X1 U9317 ( .A(n8946), .B(G21762), .Y(n8966) );
  NAND3X1 U9318 ( .A(n8969), .B(n8970), .C(n8971), .Y(G783) );
  NAND2X1 U9319 ( .A(G21386), .B(n8932), .Y(n8971) );
  NAND2X1 U9320 ( .A(n8928), .B(G21762), .Y(n8970) );
  NAND2X1 U9321 ( .A(n8946), .B(G21763), .Y(n8969) );
  NAND3X1 U9322 ( .A(n8972), .B(n8973), .C(n8974), .Y(G782) );
  NAND2X1 U9323 ( .A(G21385), .B(n8932), .Y(n8974) );
  NAND2X1 U9324 ( .A(n8928), .B(G21763), .Y(n8973) );
  NAND2X1 U9325 ( .A(n8946), .B(G21764), .Y(n8972) );
  NAND3X1 U9326 ( .A(n8975), .B(n8976), .C(n8977), .Y(G781) );
  NAND2X1 U9327 ( .A(G21384), .B(n8932), .Y(n8977) );
  NAND2X1 U9328 ( .A(n8928), .B(G21764), .Y(n8976) );
  NAND2X1 U9329 ( .A(n8946), .B(G21765), .Y(n8975) );
  NAND3X1 U9330 ( .A(n8978), .B(n8979), .C(n8980), .Y(G780) );
  NAND2X1 U9331 ( .A(G21383), .B(n8932), .Y(n8980) );
  NAND2X1 U9332 ( .A(n8928), .B(G21765), .Y(n8979) );
  NAND2X1 U9333 ( .A(n8946), .B(G21766), .Y(n8978) );
  NAND3X1 U9334 ( .A(n8981), .B(n8982), .C(n8983), .Y(G779) );
  NAND2X1 U9335 ( .A(G21382), .B(n8932), .Y(n8983) );
  NAND2X1 U9336 ( .A(n8928), .B(G21766), .Y(n8982) );
  NAND2X1 U9337 ( .A(n8946), .B(G21767), .Y(n8981) );
  NAND3X1 U9338 ( .A(n8984), .B(n8985), .C(n8986), .Y(G778) );
  NAND2X1 U9339 ( .A(G21381), .B(n8932), .Y(n8986) );
  NAND2X1 U9340 ( .A(n8928), .B(G21767), .Y(n8985) );
  NAND2X1 U9341 ( .A(n8946), .B(G21768), .Y(n8984) );
  NAND3X1 U9342 ( .A(n8987), .B(n8988), .C(n8989), .Y(G777) );
  NAND2X1 U9343 ( .A(G21380), .B(n8932), .Y(n8989) );
  NAND2X1 U9344 ( .A(n8928), .B(G21768), .Y(n8988) );
  NAND2X1 U9345 ( .A(n8946), .B(G21769), .Y(n8987) );
  NAND3X1 U9346 ( .A(n8990), .B(n8991), .C(n8992), .Y(G776) );
  NAND2X1 U9347 ( .A(G21379), .B(n8932), .Y(n8992) );
  NAND2X1 U9348 ( .A(n8928), .B(G21769), .Y(n8991) );
  NAND2X1 U9349 ( .A(n8946), .B(G21770), .Y(n8990) );
  NAND3X1 U9350 ( .A(n8993), .B(n8994), .C(n8995), .Y(G775) );
  NAND2X1 U9351 ( .A(G21378), .B(n8932), .Y(n8995) );
  NAND2X1 U9352 ( .A(n8928), .B(G21770), .Y(n8994) );
  NAND2X1 U9353 ( .A(n8946), .B(G21771), .Y(n8993) );
  NAND3X1 U9354 ( .A(n8996), .B(n8997), .C(n8998), .Y(G774) );
  NAND2X1 U9355 ( .A(G21377), .B(n8932), .Y(n8998) );
  NAND2X1 U9356 ( .A(n8928), .B(G21771), .Y(n8997) );
  NAND2X1 U9357 ( .A(n8946), .B(G21772), .Y(n8996) );
  NAND3X1 U9358 ( .A(n8999), .B(n9000), .C(n9001), .Y(G773) );
  NAND2X1 U9359 ( .A(G21376), .B(n8932), .Y(n9001) );
  NAND2X1 U9360 ( .A(n8928), .B(G21772), .Y(n9000) );
  NAND2X1 U9361 ( .A(n8946), .B(G21773), .Y(n8999) );
  NAND3X1 U9362 ( .A(n9002), .B(n9003), .C(n9004), .Y(G772) );
  NAND2X1 U9363 ( .A(G21375), .B(n8932), .Y(n9004) );
  NAND2X1 U9364 ( .A(n8928), .B(G21773), .Y(n9003) );
  NAND2X1 U9365 ( .A(n8946), .B(G21774), .Y(n9002) );
  NAND3X1 U9366 ( .A(n9005), .B(n9006), .C(n9007), .Y(G771) );
  NAND2X1 U9367 ( .A(G21374), .B(n8932), .Y(n9007) );
  NAND2X1 U9368 ( .A(n8928), .B(G21774), .Y(n9006) );
  NAND2X1 U9369 ( .A(n8946), .B(G21775), .Y(n9005) );
  NAND3X1 U9370 ( .A(n9008), .B(n9009), .C(n9010), .Y(G770) );
  NAND2X1 U9371 ( .A(G21373), .B(n8932), .Y(n9010) );
  NAND2X1 U9372 ( .A(n8928), .B(G21775), .Y(n9009) );
  NAND2X1 U9373 ( .A(n8946), .B(G21776), .Y(n9008) );
  NAND3X1 U9374 ( .A(n9011), .B(n9012), .C(n9013), .Y(G769) );
  NAND2X1 U9375 ( .A(G21372), .B(n8932), .Y(n9013) );
  NAND2X1 U9376 ( .A(n8928), .B(G21776), .Y(n9012) );
  NAND2X1 U9377 ( .A(n8946), .B(G21777), .Y(n9011) );
  NAND3X1 U9378 ( .A(n9014), .B(n9015), .C(n9016), .Y(G768) );
  NAND2X1 U9379 ( .A(G21371), .B(n8932), .Y(n9016) );
  NAND2X1 U9380 ( .A(n8928), .B(G21777), .Y(n9015) );
  NAND2X1 U9381 ( .A(n8946), .B(G21778), .Y(n9014) );
  NAND3X1 U9382 ( .A(n9017), .B(n9018), .C(n9019), .Y(G767) );
  NAND2X1 U9383 ( .A(G21370), .B(n8932), .Y(n9019) );
  NAND2X1 U9384 ( .A(n8928), .B(G21778), .Y(n9018) );
  NAND2X1 U9385 ( .A(n8946), .B(G21779), .Y(n9017) );
  NAND3X1 U9386 ( .A(n9020), .B(n9021), .C(n9022), .Y(G766) );
  NAND2X1 U9387 ( .A(G21369), .B(n8932), .Y(n9022) );
  NAND2X1 U9388 ( .A(n8928), .B(G21779), .Y(n9021) );
  NAND2X1 U9389 ( .A(n8946), .B(G21780), .Y(n9020) );
  NAND3X1 U9390 ( .A(n9023), .B(n9024), .C(n9025), .Y(G765) );
  NAND2X1 U9391 ( .A(G21368), .B(n8932), .Y(n9025) );
  NAND2X1 U9392 ( .A(n8928), .B(G21780), .Y(n9024) );
  NAND2X1 U9393 ( .A(n8946), .B(G21781), .Y(n9023) );
  NAND3X1 U9394 ( .A(n9026), .B(n9027), .C(n9028), .Y(G764) );
  NAND2X1 U9395 ( .A(G21367), .B(n8932), .Y(n9028) );
  NAND2X1 U9396 ( .A(n8928), .B(G21781), .Y(n9027) );
  NAND2X1 U9397 ( .A(n8946), .B(G21782), .Y(n9026) );
  NAND3X1 U9398 ( .A(n9029), .B(n9030), .C(n9031), .Y(G763) );
  NAND2X1 U9399 ( .A(G21366), .B(n8932), .Y(n9031) );
  NAND2X1 U9400 ( .A(n8928), .B(G21782), .Y(n9030) );
  NAND2X1 U9401 ( .A(n8946), .B(G21783), .Y(n9029) );
  NAND3X1 U9402 ( .A(n9032), .B(n9033), .C(n9034), .Y(G762) );
  NAND2X1 U9403 ( .A(G21365), .B(n8932), .Y(n9034) );
  NAND2X1 U9404 ( .A(n8928), .B(G21783), .Y(n9033) );
  NAND2X1 U9405 ( .A(n8946), .B(G21784), .Y(n9032) );
  NAND3X1 U9406 ( .A(n9035), .B(n9036), .C(n9037), .Y(G761) );
  NAND2X1 U9407 ( .A(G21364), .B(n8932), .Y(n9037) );
  NAND2X1 U9408 ( .A(n8928), .B(G21784), .Y(n9036) );
  NAND2X1 U9409 ( .A(n8946), .B(G21785), .Y(n9035) );
  NAND3X1 U9410 ( .A(n9038), .B(n9039), .C(n9040), .Y(G760) );
  NAND2X1 U9411 ( .A(G21363), .B(n8932), .Y(n9040) );
  NAND2X1 U9412 ( .A(n8928), .B(G21785), .Y(n9039) );
  NAND2X1 U9413 ( .A(n8946), .B(G21786), .Y(n9038) );
  NAND3X1 U9414 ( .A(n9041), .B(n9042), .C(n9043), .Y(G759) );
  NAND2X1 U9415 ( .A(G21362), .B(n8932), .Y(n9043) );
  NAND2X1 U9416 ( .A(n8928), .B(G21786), .Y(n9042) );
  NAND2X1 U9417 ( .A(n8946), .B(G21787), .Y(n9041) );
  NAND3X1 U9418 ( .A(n9044), .B(n9045), .C(n9046), .Y(G758) );
  NAND2X1 U9419 ( .A(G21361), .B(n8932), .Y(n9046) );
  NAND2X1 U9420 ( .A(n8928), .B(G21787), .Y(n9045) );
  NAND2X1 U9421 ( .A(n8946), .B(G21788), .Y(n9044) );
  NAND3X1 U9422 ( .A(n9047), .B(n9048), .C(n9049), .Y(G757) );
  NAND2X1 U9423 ( .A(G21360), .B(n8932), .Y(n9049) );
  NAND2X1 U9424 ( .A(n8928), .B(G21788), .Y(n9048) );
  NAND2X1 U9425 ( .A(n8946), .B(G21789), .Y(n9047) );
  NAND2X1 U9426 ( .A(n9050), .B(n9051), .Y(G1751) );
  NAND2X1 U9427 ( .A(G21804), .B(n9052), .Y(n9051) );
  OR2X1 U9428 ( .A(n9052), .B(n9053), .Y(n9050) );
  NAND2X1 U9429 ( .A(n9054), .B(n9055), .Y(G1750) );
  NAND2X1 U9430 ( .A(n9052), .B(G21803), .Y(n9055) );
  OR2X1 U9431 ( .A(n9056), .B(n9052), .Y(n9054) );
  NOR2X1 U9432 ( .A(n9057), .B(n9058), .Y(n9052) );
  NOR3X1 U9433 ( .A(n9059), .B(n9060), .C(n7430), .Y(n9056) );
  NAND2X1 U9434 ( .A(n9061), .B(n9062), .Y(G1749) );
  NAND2X1 U9435 ( .A(G21800), .B(n8932), .Y(n9062) );
  NAND2X1 U9436 ( .A(G21804), .B(n8947), .Y(n9061) );
  NAND2X1 U9437 ( .A(n9063), .B(n9064), .Y(G1748) );
  OR2X1 U9438 ( .A(n9065), .B(n8945), .Y(n9064) );
  INVX1 U9439 ( .A(G21798), .Y(n8945) );
  NAND2X1 U9440 ( .A(n9066), .B(n9065), .Y(n9063) );
  NAND3X1 U9441 ( .A(n9067), .B(n9068), .C(n9069), .Y(n9065) );
  NAND3X1 U9442 ( .A(n8897), .B(n9070), .C(n8896), .Y(n9068) );
  NAND2X1 U9443 ( .A(G21428), .B(G21426), .Y(n8896) );
  NAND3X1 U9444 ( .A(G21427), .B(n7445), .C(n9071), .Y(n9067) );
  NAND2X1 U9445 ( .A(n8783), .B(n9072), .Y(n9066) );
  NAND2X1 U9446 ( .A(G21428), .B(n9073), .Y(n9072) );
  NAND4X1 U9447 ( .A(G21426), .B(n9074), .C(n9075), .D(n7445), .Y(n9073) );
  OR3X1 U9448 ( .A(n9076), .B(G21797), .C(n7444), .Y(n9075) );
  OR2X1 U9449 ( .A(n7454), .B(n9077), .Y(n9074) );
  NAND2X1 U9450 ( .A(n9078), .B(n9079), .Y(G1747) );
  OR2X1 U9451 ( .A(n8932), .B(G21803), .Y(n9079) );
  NAND2X1 U9452 ( .A(G21794), .B(n8932), .Y(n9078) );
  NAND4X1 U9453 ( .A(n9080), .B(n9081), .C(n9082), .D(n9083), .Y(G1746) );
  NAND3X1 U9454 ( .A(G21428), .B(n7457), .C(n7475), .Y(n9083) );
  NAND2X1 U9455 ( .A(n7462), .B(G21566), .Y(n9082) );
  NAND3X1 U9456 ( .A(n9084), .B(n7430), .C(n7463), .Y(n9081) );
  NOR2X1 U9457 ( .A(n9085), .B(n7462), .Y(n7463) );
  INVX1 U9458 ( .A(n7475), .Y(n7462) );
  NAND2X1 U9459 ( .A(n7465), .B(n7001), .Y(n9080) );
  AND2X1 U9460 ( .A(n9086), .B(n7475), .Y(n7465) );
  NAND3X1 U9461 ( .A(n9087), .B(n9088), .C(n8784), .Y(n7475) );
  INVX1 U9462 ( .A(n7580), .Y(n8784) );
  NAND3X1 U9463 ( .A(n9089), .B(n9090), .C(n9091), .Y(n7580) );
  OR2X1 U9464 ( .A(n8832), .B(n9092), .Y(n9091) );
  NAND2X1 U9465 ( .A(n9071), .B(n9093), .Y(n9090) );
  NAND3X1 U9466 ( .A(n7430), .B(n8817), .C(G21427), .Y(n9089) );
  NAND2X1 U9467 ( .A(n8898), .B(n9092), .Y(n9087) );
  NAND2X1 U9468 ( .A(n8829), .B(n9094), .Y(n9086) );
  NAND2X1 U9469 ( .A(n9085), .B(n7430), .Y(n9094) );
  NAND2X1 U9470 ( .A(n9095), .B(n9096), .Y(G1745) );
  NAND2X1 U9471 ( .A(n9097), .B(G21561), .Y(n9096) );
  NAND2X1 U9472 ( .A(n9098), .B(n9099), .Y(n9095) );
  NAND3X1 U9473 ( .A(n9100), .B(n9101), .C(n9102), .Y(n9098) );
  NAND2X1 U9474 ( .A(n8818), .B(n8884), .Y(n9102) );
  NAND3X1 U9475 ( .A(n9103), .B(n9104), .C(n9105), .Y(n8884) );
  NOR3X1 U9476 ( .A(n9106), .B(n9107), .C(n9108), .Y(n9105) );
  NOR2X1 U9477 ( .A(n9109), .B(n9110), .Y(n9108) );
  AND2X1 U9478 ( .A(n8890), .B(n8855), .Y(n9107) );
  NOR2X1 U9479 ( .A(n9111), .B(n9112), .Y(n9106) );
  NAND2X1 U9480 ( .A(n7001), .B(n9113), .Y(n9104) );
  NAND2X1 U9481 ( .A(n7003), .B(n9114), .Y(n9103) );
  NAND2X1 U9482 ( .A(G21427), .B(n9115), .Y(n9101) );
  NAND2X1 U9483 ( .A(G21567), .B(n9112), .Y(n9115) );
  NAND2X1 U9484 ( .A(n9116), .B(n7003), .Y(n9100) );
  NAND2X1 U9485 ( .A(n9117), .B(n9118), .Y(G1744) );
  NAND2X1 U9486 ( .A(n9097), .B(G21560), .Y(n9118) );
  NAND2X1 U9487 ( .A(n9119), .B(n9099), .Y(n9117) );
  NAND3X1 U9488 ( .A(n9120), .B(n9121), .C(n9122), .Y(n9119) );
  NAND2X1 U9489 ( .A(n9123), .B(n9124), .Y(n9122) );
  NAND2X1 U9490 ( .A(n9116), .B(n6992), .Y(n9121) );
  NAND2X1 U9491 ( .A(n8818), .B(n8883), .Y(n9120) );
  NAND4X1 U9492 ( .A(n9125), .B(n9126), .C(n9127), .D(n9128), .Y(n8883) );
  NOR3X1 U9493 ( .A(n9129), .B(n9130), .C(n9131), .Y(n9128) );
  NOR2X1 U9494 ( .A(n9109), .B(n9132), .Y(n9131) );
  NOR2X1 U9495 ( .A(n9133), .B(n9134), .Y(n9130) );
  NOR2X1 U9496 ( .A(n9135), .B(n9136), .Y(n9133) );
  NOR2X1 U9497 ( .A(n9111), .B(n9137), .Y(n9129) );
  NAND2X1 U9498 ( .A(n9138), .B(n9139), .Y(n9127) );
  NAND2X1 U9499 ( .A(n6990), .B(n9113), .Y(n9126) );
  NAND2X1 U9500 ( .A(n6992), .B(n9114), .Y(n9125) );
  NAND2X1 U9501 ( .A(n9140), .B(n9141), .Y(G1743) );
  NAND2X1 U9502 ( .A(n9097), .B(G21559), .Y(n9141) );
  NAND2X1 U9503 ( .A(n9142), .B(n9099), .Y(n9140) );
  NAND3X1 U9504 ( .A(n9143), .B(n9144), .C(n9145), .Y(n9142) );
  NAND2X1 U9505 ( .A(n9123), .B(n9146), .Y(n9145) );
  NAND2X1 U9506 ( .A(n9116), .B(n6981), .Y(n9144) );
  NAND2X1 U9507 ( .A(n8818), .B(n8894), .Y(n9143) );
  NAND4X1 U9508 ( .A(n9147), .B(n9148), .C(n9149), .D(n9150), .Y(n8894) );
  NOR3X1 U9509 ( .A(n9151), .B(n9152), .C(n9153), .Y(n9150) );
  NOR2X1 U9510 ( .A(n9111), .B(n9154), .Y(n9153) );
  NOR2X1 U9511 ( .A(n9109), .B(n9155), .Y(n9152) );
  NOR2X1 U9512 ( .A(n9156), .B(n7392), .Y(n9151) );
  NAND2X1 U9513 ( .A(n9138), .B(n9157), .Y(n9149) );
  NAND2X1 U9514 ( .A(n9114), .B(n6981), .Y(n9148) );
  NAND2X1 U9515 ( .A(n9158), .B(n7420), .Y(n9147) );
  NAND2X1 U9516 ( .A(n9159), .B(n9160), .Y(G1742) );
  NAND2X1 U9517 ( .A(n9097), .B(G21558), .Y(n9160) );
  NAND2X1 U9518 ( .A(n9161), .B(n9099), .Y(n9159) );
  NAND2X1 U9519 ( .A(n9162), .B(n9163), .Y(n9161) );
  NAND2X1 U9520 ( .A(n9116), .B(n6971), .Y(n9163) );
  NOR2X1 U9521 ( .A(n9092), .B(G21426), .Y(n9116) );
  NAND2X1 U9522 ( .A(n8818), .B(n8871), .Y(n9162) );
  NAND4X1 U9523 ( .A(n9164), .B(n9165), .C(n9166), .D(n9167), .Y(n8871) );
  NOR3X1 U9524 ( .A(n9168), .B(n9169), .C(n9170), .Y(n9167) );
  NOR2X1 U9525 ( .A(n9111), .B(n9171), .Y(n9170) );
  AND2X1 U9526 ( .A(n9172), .B(n7429), .Y(n9111) );
  NOR2X1 U9527 ( .A(n9109), .B(n9173), .Y(n9169) );
  NOR2X1 U9528 ( .A(n9174), .B(n9175), .Y(n9109) );
  NOR2X1 U9529 ( .A(n9156), .B(n9176), .Y(n9168) );
  INVX1 U9530 ( .A(n9113), .Y(n9156) );
  NAND3X1 U9531 ( .A(n7413), .B(n7414), .C(n9177), .Y(n9113) );
  NOR3X1 U9532 ( .A(n9178), .B(n7418), .C(n7419), .Y(n9177) );
  NOR4X1 U9533 ( .A(n8782), .B(n7456), .C(n7444), .D(n9076), .Y(n7419) );
  NOR2X1 U9534 ( .A(n7451), .B(n9179), .Y(n9178) );
  AND4X1 U9535 ( .A(n9180), .B(n9181), .C(n9182), .D(n9183), .Y(n7414) );
  NAND2X1 U9536 ( .A(n9184), .B(n8782), .Y(n9183) );
  NAND2X1 U9537 ( .A(n9185), .B(n7458), .Y(n9182) );
  NAND3X1 U9538 ( .A(n7444), .B(n8711), .C(n7456), .Y(n9181) );
  INVX1 U9539 ( .A(n9186), .Y(n9180) );
  AND3X1 U9540 ( .A(n9187), .B(n9188), .C(n9189), .Y(n7413) );
  NAND2X1 U9541 ( .A(n7446), .B(n9190), .Y(n9189) );
  NAND2X1 U9542 ( .A(n9191), .B(n9192), .Y(n9190) );
  OR2X1 U9543 ( .A(n9193), .B(n9194), .Y(n9191) );
  NAND2X1 U9544 ( .A(n9076), .B(n9195), .Y(n9188) );
  NAND2X1 U9545 ( .A(n9196), .B(n9138), .Y(n9166) );
  NAND2X1 U9546 ( .A(n6971), .B(n9114), .Y(n9165) );
  NAND4X1 U9547 ( .A(n9197), .B(n9198), .C(n7426), .D(n7424), .Y(n9114) );
  NAND2X1 U9548 ( .A(n9199), .B(n7458), .Y(n9198) );
  NAND2X1 U9549 ( .A(n9200), .B(n9201), .Y(n9199) );
  NAND2X1 U9550 ( .A(n9202), .B(n9203), .Y(n9201) );
  NAND2X1 U9551 ( .A(n7420), .B(n9204), .Y(n9164) );
  INVX1 U9552 ( .A(n9134), .Y(n7420) );
  NAND2X1 U9553 ( .A(n9205), .B(n9206), .Y(G1740) );
  NAND4X1 U9554 ( .A(n6961), .B(n9207), .C(n8818), .D(n9099), .Y(n9206) );
  NAND2X1 U9555 ( .A(n9097), .B(G21557), .Y(n9205) );
  INVX1 U9556 ( .A(n9099), .Y(n9097) );
  NAND3X1 U9557 ( .A(n8832), .B(n9088), .C(n9208), .Y(n9099) );
  NAND2X1 U9558 ( .A(n7433), .B(n8849), .Y(n9208) );
  NAND4X1 U9559 ( .A(n7435), .B(n9209), .C(n9210), .D(n9211), .Y(n8849) );
  NAND3X1 U9560 ( .A(n7441), .B(n7445), .C(n9212), .Y(n9211) );
  NAND2X1 U9561 ( .A(n7447), .B(n9213), .Y(n9210) );
  NAND2X1 U9562 ( .A(n7424), .B(n9214), .Y(n9213) );
  NAND2X1 U9563 ( .A(n7454), .B(n9215), .Y(n9214) );
  NAND2X1 U9564 ( .A(n9187), .B(n9216), .Y(n9215) );
  NAND2X1 U9565 ( .A(n7457), .B(n8855), .Y(n9209) );
  NAND2X1 U9566 ( .A(n7428), .B(n9134), .Y(n8855) );
  AND4X1 U9567 ( .A(n9217), .B(n9218), .C(n9219), .D(n9220), .Y(n7435) );
  NOR2X1 U9568 ( .A(n9221), .B(n9222), .Y(n9220) );
  ADDHXL U9569 ( .A(n8762), .B(n9223), .S(n9222) );
  NAND2X1 U9570 ( .A(n9224), .B(n7446), .Y(n9217) );
  NAND2X1 U9571 ( .A(n8898), .B(G21795), .Y(n9088) );
  NOR2X1 U9572 ( .A(n8897), .B(n8817), .Y(n8898) );
  NAND2X1 U9573 ( .A(G21425), .B(n8817), .Y(n8832) );
  NAND2X1 U9574 ( .A(n9225), .B(n9226), .Y(G1738) );
  NAND2X1 U9575 ( .A(G21394), .B(n8916), .Y(n9226) );
  NAND2X1 U9576 ( .A(n9227), .B(n8899), .Y(n9225) );
  NAND2X1 U9577 ( .A(n9228), .B(n9229), .Y(n9227) );
  NAND2X1 U9578 ( .A(n9230), .B(n9231), .Y(G1737) );
  NAND3X1 U9579 ( .A(n9229), .B(n9228), .C(n8899), .Y(n9231) );
  INVX1 U9580 ( .A(G34), .Y(n9228) );
  INVX1 U9581 ( .A(n8925), .Y(n9229) );
  NAND2X1 U9582 ( .A(G21393), .B(n8916), .Y(n9230) );
  NAND2X1 U9583 ( .A(n9232), .B(n9233), .Y(G1735) );
  NAND2X1 U9584 ( .A(G21359), .B(n8932), .Y(n9233) );
  NAND2X1 U9585 ( .A(G21793), .B(n8947), .Y(n9232) );
  NAND2X1 U9586 ( .A(n9234), .B(n9235), .Y(G1734) );
  NAND2X1 U9587 ( .A(G21358), .B(n8932), .Y(n9235) );
  NAND2X1 U9588 ( .A(G21792), .B(n8947), .Y(n9234) );
  NAND2X1 U9589 ( .A(n9236), .B(n9237), .Y(G1733) );
  NAND2X1 U9590 ( .A(G21357), .B(n8932), .Y(n9237) );
  NAND2X1 U9591 ( .A(G21791), .B(n8947), .Y(n9236) );
  NAND2X1 U9592 ( .A(n9238), .B(n9239), .Y(G1732) );
  NAND2X1 U9593 ( .A(G21356), .B(n8932), .Y(n9239) );
  NAND2X1 U9594 ( .A(G21790), .B(n8947), .Y(n9238) );
  NAND2X1 U9595 ( .A(n8916), .B(n9240), .Y(G1189) );
  NAND2X1 U9596 ( .A(G21802), .B(G21392), .Y(n9240) );
  NAND2X1 U9597 ( .A(n9241), .B(n9242), .Y(G1188) );
  NAND2X1 U9598 ( .A(G21801), .B(n9243), .Y(n9242) );
  NAND2X1 U9599 ( .A(n9244), .B(n7433), .Y(n9243) );
  NAND2X1 U9600 ( .A(n9058), .B(G21428), .Y(n9241) );
  NAND3X1 U9601 ( .A(n9245), .B(n9246), .C(n9247), .Y(G1187) );
  OR2X1 U9602 ( .A(n8932), .B(G21801), .Y(n9246) );
  NAND2X1 U9603 ( .A(G21799), .B(n8932), .Y(n9245) );
  NOR2X1 U9604 ( .A(n8938), .B(G21392), .Y(n8947) );
  NAND3X1 U9605 ( .A(n9248), .B(n9249), .C(n9247), .Y(G1186) );
  NAND2X1 U9606 ( .A(n8925), .B(n8938), .Y(n9247) );
  NOR2X1 U9607 ( .A(G21392), .B(G21390), .Y(n8925) );
  NAND2X1 U9608 ( .A(G34), .B(n8899), .Y(n9249) );
  NAND2X1 U9609 ( .A(n8916), .B(G21797), .Y(n9248) );
  INVX1 U9610 ( .A(n8899), .Y(n8916) );
  NAND2X1 U9611 ( .A(n9250), .B(n8958), .Y(n8899) );
  NAND2X1 U9612 ( .A(G21392), .B(n8929), .Y(n8958) );
  NAND2X1 U9613 ( .A(n8959), .B(n8938), .Y(n9250) );
  INVX1 U9614 ( .A(G21392), .Y(n8959) );
  NAND2X1 U9615 ( .A(n9251), .B(n9252), .Y(G1185) );
  NAND2X1 U9616 ( .A(n9253), .B(n8860), .Y(n9252) );
  NAND2X1 U9617 ( .A(n9254), .B(n9255), .Y(n9253) );
  NAND2X1 U9618 ( .A(n9256), .B(n9257), .Y(n9255) );
  NAND2X1 U9619 ( .A(n9258), .B(n9259), .Y(n9256) );
  NAND2X1 U9620 ( .A(n8818), .B(n9260), .Y(n9259) );
  NAND2X1 U9621 ( .A(n9092), .B(n9261), .Y(n9254) );
  NAND3X1 U9622 ( .A(n9262), .B(n9263), .C(n9264), .Y(n9261) );
  NAND2X1 U9623 ( .A(n7433), .B(n8856), .Y(n9264) );
  NAND2X1 U9624 ( .A(n8818), .B(n9265), .Y(n9262) );
  NAND2X1 U9625 ( .A(n9266), .B(n9267), .Y(n9265) );
  NAND2X1 U9626 ( .A(G21796), .B(n9268), .Y(n9251) );
  NAND2X1 U9627 ( .A(n9269), .B(n9270), .Y(G1184) );
  NAND2X1 U9628 ( .A(G21795), .B(n9268), .Y(n9270) );
  NAND2X1 U9629 ( .A(n7433), .B(n8860), .Y(n9268) );
  NAND2X1 U9630 ( .A(n9244), .B(n9271), .Y(n8860) );
  NAND2X1 U9631 ( .A(n9272), .B(n7445), .Y(n9271) );
  NAND2X1 U9632 ( .A(n9273), .B(n9274), .Y(n9272) );
  ADDHXL U9633 ( .A(n7451), .B(n7456), .S(n9273) );
  AND4X1 U9634 ( .A(n9275), .B(n9276), .C(n9277), .D(n9278), .Y(n9244) );
  NAND2X1 U9635 ( .A(n7439), .B(n9279), .Y(n9277) );
  NAND3X1 U9636 ( .A(n7455), .B(n9280), .C(n9281), .Y(n9279) );
  NAND2X1 U9637 ( .A(n7444), .B(n9257), .Y(n9280) );
  NAND2X1 U9638 ( .A(n9092), .B(n9282), .Y(n9276) );
  NAND2X1 U9639 ( .A(n7439), .B(n7444), .Y(n9282) );
  INVX1 U9640 ( .A(n9221), .Y(n9275) );
  NAND3X1 U9641 ( .A(n9193), .B(n8782), .C(n9283), .Y(n9221) );
  NAND2X1 U9642 ( .A(n7456), .B(n9284), .Y(n9283) );
  NAND2X1 U9643 ( .A(n9285), .B(n9076), .Y(n9284) );
  NAND3X1 U9644 ( .A(n9286), .B(n9287), .C(n9288), .Y(G1183) );
  NAND2X1 U9645 ( .A(G21793), .B(n9289), .Y(n9287) );
  OR2X1 U9646 ( .A(n9289), .B(n7000), .Y(n9286) );
  NAND3X1 U9647 ( .A(n9288), .B(n9290), .C(n9291), .Y(G1182) );
  NAND2X1 U9648 ( .A(G21792), .B(n9289), .Y(n9291) );
  INVX1 U9649 ( .A(n9292), .Y(n9288) );
  NAND3X1 U9650 ( .A(n9293), .B(n9294), .C(n9295), .Y(G1181) );
  NAND2X1 U9651 ( .A(G21791), .B(n9289), .Y(n9295) );
  NAND3X1 U9652 ( .A(n9296), .B(n6989), .C(n9297), .Y(n9294) );
  NAND2X1 U9653 ( .A(G21393), .B(G21758), .Y(n9296) );
  NAND2X1 U9654 ( .A(n9292), .B(G21758), .Y(n9293) );
  NOR2X1 U9655 ( .A(n9289), .B(n6989), .Y(n9292) );
  NAND3X1 U9656 ( .A(n9298), .B(n9290), .C(n9299), .Y(G1180) );
  NAND2X1 U9657 ( .A(G21790), .B(n9289), .Y(n9299) );
  NAND3X1 U9658 ( .A(n9300), .B(n7000), .C(n9297), .Y(n9290) );
  INVX1 U9659 ( .A(G21758), .Y(n7000) );
  INVX1 U9660 ( .A(G21393), .Y(n9300) );
  NAND2X1 U9661 ( .A(n9297), .B(n6989), .Y(n9298) );
  NOR2X1 U9662 ( .A(n9289), .B(G21394), .Y(n9297) );
  NAND4X1 U9663 ( .A(n9301), .B(n9302), .C(n9303), .D(n9304), .Y(n9289) );
  NOR4X1 U9664 ( .A(n9305), .B(n9306), .C(n9307), .D(n9308), .Y(n9304) );
  NAND4X1 U9665 ( .A(n8915), .B(n8914), .C(n8913), .D(n8912), .Y(n9308) );
  INVX1 U9666 ( .A(G21412), .Y(n8912) );
  INVX1 U9667 ( .A(G21411), .Y(n8913) );
  INVX1 U9668 ( .A(G21410), .Y(n8914) );
  INVX1 U9669 ( .A(G21409), .Y(n8915) );
  NAND4X1 U9670 ( .A(n8911), .B(n8910), .C(n8909), .D(n8908), .Y(n9307) );
  INVX1 U9671 ( .A(G21416), .Y(n8908) );
  INVX1 U9672 ( .A(G21415), .Y(n8909) );
  INVX1 U9673 ( .A(G21414), .Y(n8910) );
  INVX1 U9674 ( .A(G21413), .Y(n8911) );
  NAND4X1 U9675 ( .A(n8907), .B(n8906), .C(n8905), .D(n8904), .Y(n9306) );
  INVX1 U9676 ( .A(G21420), .Y(n8904) );
  INVX1 U9677 ( .A(G21419), .Y(n8905) );
  INVX1 U9678 ( .A(G21418), .Y(n8906) );
  INVX1 U9679 ( .A(G21417), .Y(n8907) );
  NAND4X1 U9680 ( .A(n8903), .B(n8902), .C(n8901), .D(n8900), .Y(n9305) );
  INVX1 U9681 ( .A(G21424), .Y(n8900) );
  INVX1 U9682 ( .A(G21423), .Y(n8901) );
  INVX1 U9683 ( .A(G21422), .Y(n8902) );
  INVX1 U9684 ( .A(G21421), .Y(n8903) );
  NOR4X1 U9685 ( .A(n9309), .B(n9310), .C(G21396), .D(G21395), .Y(n9303) );
  AND2X1 U9686 ( .A(G21394), .B(G21393), .Y(n9310) );
  NAND4X1 U9687 ( .A(n8920), .B(n8919), .C(n8918), .D(n8917), .Y(n9309) );
  INVX1 U9688 ( .A(G21400), .Y(n8917) );
  INVX1 U9689 ( .A(G21399), .Y(n8918) );
  INVX1 U9690 ( .A(G21398), .Y(n8919) );
  INVX1 U9691 ( .A(G21397), .Y(n8920) );
  NOR4X1 U9692 ( .A(G21408), .B(G21407), .C(G21406), .D(G21405), .Y(n9302) );
  NOR4X1 U9693 ( .A(G21404), .B(G21403), .C(G21402), .D(G21401), .Y(n9301) );
  NAND4X1 U9694 ( .A(n9311), .B(n9312), .C(n9313), .D(n9314), .Y(G1179) );
  NOR3X1 U9695 ( .A(n9315), .B(n9316), .C(n9317), .Y(n9314) );
  NOR2X1 U9696 ( .A(n9318), .B(n9319), .Y(n9317) );
  NOR2X1 U9697 ( .A(n9320), .B(n9321), .Y(n9316) );
  NOR2X1 U9698 ( .A(n9322), .B(n9323), .Y(n9315) );
  NAND2X1 U9699 ( .A(n9324), .B(G21789), .Y(n9313) );
  NAND2X1 U9700 ( .A(n7025), .B(n9325), .Y(n9312) );
  NAND2X1 U9701 ( .A(n9326), .B(n7021), .Y(n9311) );
  NAND4X1 U9702 ( .A(n9327), .B(n9328), .C(n9329), .D(n9330), .Y(G1178) );
  NOR3X1 U9703 ( .A(n9331), .B(n9332), .C(n9333), .Y(n9330) );
  NOR2X1 U9704 ( .A(n9334), .B(n9319), .Y(n9333) );
  NOR2X1 U9705 ( .A(n9335), .B(n9321), .Y(n9332) );
  INVX1 U9706 ( .A(G21756), .Y(n9335) );
  NOR2X1 U9707 ( .A(n9322), .B(n9336), .Y(n9331) );
  NAND2X1 U9708 ( .A(n9324), .B(G21788), .Y(n9329) );
  NAND2X1 U9709 ( .A(n7039), .B(n9325), .Y(n9328) );
  NAND2X1 U9710 ( .A(n9326), .B(n7037), .Y(n9327) );
  NAND4X1 U9711 ( .A(n9337), .B(n9338), .C(n9339), .D(n9340), .Y(G1177) );
  NOR3X1 U9712 ( .A(n9341), .B(n9342), .C(n9343), .Y(n9340) );
  NOR2X1 U9713 ( .A(n9344), .B(n9319), .Y(n9343) );
  NOR2X1 U9714 ( .A(n9345), .B(n9321), .Y(n9342) );
  NOR2X1 U9715 ( .A(n9322), .B(n7048), .Y(n9341) );
  NAND2X1 U9716 ( .A(n9324), .B(G21787), .Y(n9339) );
  NAND2X1 U9717 ( .A(n9346), .B(n9325), .Y(n9338) );
  NAND2X1 U9718 ( .A(n9326), .B(n7053), .Y(n9337) );
  NAND4X1 U9719 ( .A(n9347), .B(n9348), .C(n9349), .D(n9350), .Y(G1176) );
  NOR3X1 U9720 ( .A(n9351), .B(n9352), .C(n9353), .Y(n9350) );
  NOR2X1 U9721 ( .A(n9354), .B(n9319), .Y(n9353) );
  NOR2X1 U9722 ( .A(n9355), .B(n9321), .Y(n9352) );
  INVX1 U9723 ( .A(G21754), .Y(n9355) );
  NOR2X1 U9724 ( .A(n9322), .B(n9356), .Y(n9351) );
  NAND2X1 U9725 ( .A(n9324), .B(G21786), .Y(n9349) );
  NAND2X1 U9726 ( .A(n7067), .B(n9325), .Y(n9348) );
  NAND2X1 U9727 ( .A(n9326), .B(n7065), .Y(n9347) );
  NAND4X1 U9728 ( .A(n9357), .B(n9358), .C(n9359), .D(n9360), .Y(G1175) );
  NOR3X1 U9729 ( .A(n9361), .B(n9362), .C(n9363), .Y(n9360) );
  NOR2X1 U9730 ( .A(n9364), .B(n9319), .Y(n9363) );
  NOR2X1 U9731 ( .A(n9365), .B(n9321), .Y(n9362) );
  INVX1 U9732 ( .A(G21753), .Y(n9365) );
  NOR2X1 U9733 ( .A(n9322), .B(n7075), .Y(n9361) );
  NAND2X1 U9734 ( .A(n9324), .B(G21785), .Y(n9359) );
  NAND2X1 U9735 ( .A(n9366), .B(n9325), .Y(n9358) );
  NAND2X1 U9736 ( .A(n9326), .B(n7079), .Y(n9357) );
  NAND4X1 U9737 ( .A(n9367), .B(n9368), .C(n9369), .D(n9370), .Y(G1174) );
  NOR3X1 U9738 ( .A(n9371), .B(n9372), .C(n9373), .Y(n9370) );
  NOR2X1 U9739 ( .A(n9374), .B(n9319), .Y(n9373) );
  NOR2X1 U9740 ( .A(n9375), .B(n9321), .Y(n9372) );
  INVX1 U9741 ( .A(G21752), .Y(n9375) );
  NOR2X1 U9742 ( .A(n9322), .B(n7087), .Y(n9371) );
  NAND2X1 U9743 ( .A(n9324), .B(G21784), .Y(n9369) );
  NAND2X1 U9744 ( .A(n9376), .B(n9325), .Y(n9368) );
  NAND2X1 U9745 ( .A(n9326), .B(n7091), .Y(n9367) );
  NAND4X1 U9746 ( .A(n9377), .B(n9378), .C(n9379), .D(n9380), .Y(G1173) );
  NOR3X1 U9747 ( .A(n9381), .B(n9382), .C(n9383), .Y(n9380) );
  NOR2X1 U9748 ( .A(n9384), .B(n9319), .Y(n9383) );
  NOR2X1 U9749 ( .A(n9385), .B(n9321), .Y(n9382) );
  INVX1 U9750 ( .A(G21751), .Y(n9385) );
  NOR2X1 U9751 ( .A(n9322), .B(n9386), .Y(n9381) );
  NAND2X1 U9752 ( .A(n9324), .B(G21783), .Y(n9379) );
  NAND2X1 U9753 ( .A(n7104), .B(n9325), .Y(n9378) );
  NAND2X1 U9754 ( .A(n9326), .B(n7102), .Y(n9377) );
  NAND4X1 U9755 ( .A(n9387), .B(n9388), .C(n9389), .D(n9390), .Y(G1172) );
  NOR3X1 U9756 ( .A(n9391), .B(n9392), .C(n9393), .Y(n9390) );
  NOR2X1 U9757 ( .A(n9394), .B(n9319), .Y(n9393) );
  NOR2X1 U9758 ( .A(n9395), .B(n9321), .Y(n9392) );
  INVX1 U9759 ( .A(G21750), .Y(n9395) );
  NOR2X1 U9760 ( .A(n9322), .B(n7112), .Y(n9391) );
  NAND2X1 U9761 ( .A(n9324), .B(G21782), .Y(n9389) );
  NAND2X1 U9762 ( .A(n9396), .B(n9325), .Y(n9388) );
  NAND2X1 U9763 ( .A(n9326), .B(n7115), .Y(n9387) );
  NAND4X1 U9764 ( .A(n9397), .B(n9398), .C(n9399), .D(n9400), .Y(G1171) );
  NOR3X1 U9765 ( .A(n9401), .B(n9402), .C(n9403), .Y(n9400) );
  NOR2X1 U9766 ( .A(n9404), .B(n9319), .Y(n9403) );
  NOR2X1 U9767 ( .A(n9405), .B(n9321), .Y(n9402) );
  INVX1 U9768 ( .A(G21749), .Y(n9405) );
  NOR2X1 U9769 ( .A(n9322), .B(n9406), .Y(n9401) );
  NAND2X1 U9770 ( .A(n9324), .B(G21781), .Y(n9399) );
  NAND2X1 U9771 ( .A(n7127), .B(n9325), .Y(n9398) );
  NAND2X1 U9772 ( .A(n9326), .B(n7125), .Y(n9397) );
  NAND4X1 U9773 ( .A(n9407), .B(n9408), .C(n9409), .D(n9410), .Y(G1170) );
  NOR3X1 U9774 ( .A(n9411), .B(n9412), .C(n9413), .Y(n9410) );
  NOR2X1 U9775 ( .A(n9414), .B(n9319), .Y(n9413) );
  NOR2X1 U9776 ( .A(n9415), .B(n9321), .Y(n9412) );
  INVX1 U9777 ( .A(G21748), .Y(n9415) );
  NOR2X1 U9778 ( .A(n9322), .B(n9416), .Y(n9411) );
  NAND2X1 U9779 ( .A(n9324), .B(G21780), .Y(n9409) );
  NAND2X1 U9780 ( .A(n7140), .B(n9325), .Y(n9408) );
  NAND2X1 U9781 ( .A(n9326), .B(n7138), .Y(n9407) );
  NAND4X1 U9782 ( .A(n9417), .B(n9418), .C(n9419), .D(n9420), .Y(G1169) );
  NOR3X1 U9783 ( .A(n9421), .B(n9422), .C(n9423), .Y(n9420) );
  NOR2X1 U9784 ( .A(n9424), .B(n9319), .Y(n9423) );
  NOR2X1 U9785 ( .A(n9425), .B(n9321), .Y(n9422) );
  INVX1 U9786 ( .A(G21747), .Y(n9425) );
  NOR2X1 U9787 ( .A(n9322), .B(n9426), .Y(n9421) );
  NAND2X1 U9788 ( .A(n9324), .B(G21779), .Y(n9419) );
  NAND2X1 U9789 ( .A(n7153), .B(n9325), .Y(n9418) );
  NAND2X1 U9790 ( .A(n9326), .B(n7151), .Y(n9417) );
  NAND4X1 U9791 ( .A(n9427), .B(n9428), .C(n9429), .D(n9430), .Y(G1168) );
  NOR3X1 U9792 ( .A(n9431), .B(n9432), .C(n9433), .Y(n9430) );
  NOR2X1 U9793 ( .A(n9434), .B(n9319), .Y(n9433) );
  NOR2X1 U9794 ( .A(n9435), .B(n9321), .Y(n9432) );
  INVX1 U9795 ( .A(G21746), .Y(n9435) );
  NOR2X1 U9796 ( .A(n9322), .B(n9436), .Y(n9431) );
  NAND2X1 U9797 ( .A(n9324), .B(G21778), .Y(n9429) );
  NAND2X1 U9798 ( .A(n7165), .B(n9325), .Y(n9428) );
  NAND2X1 U9799 ( .A(n9326), .B(n7163), .Y(n9427) );
  NAND4X1 U9800 ( .A(n9437), .B(n9438), .C(n9439), .D(n9440), .Y(G1167) );
  NOR4X1 U9801 ( .A(n9441), .B(n9442), .C(n9443), .D(n9444), .Y(n9440) );
  NOR2X1 U9802 ( .A(n9322), .B(n9445), .Y(n9444) );
  NOR2X1 U9803 ( .A(n9446), .B(n9319), .Y(n9443) );
  NOR2X1 U9804 ( .A(n9447), .B(n9321), .Y(n9442) );
  INVX1 U9805 ( .A(G21745), .Y(n9447) );
  NAND2X1 U9806 ( .A(n9324), .B(G21777), .Y(n9439) );
  NAND2X1 U9807 ( .A(n7178), .B(n9325), .Y(n9438) );
  NAND2X1 U9808 ( .A(n9326), .B(n7176), .Y(n9437) );
  NAND4X1 U9809 ( .A(n9448), .B(n9449), .C(n9450), .D(n9451), .Y(G1166) );
  NOR4X1 U9810 ( .A(n9441), .B(n9452), .C(n9453), .D(n9454), .Y(n9451) );
  NOR2X1 U9811 ( .A(n9322), .B(n9455), .Y(n9454) );
  NOR2X1 U9812 ( .A(n9456), .B(n9319), .Y(n9453) );
  NOR2X1 U9813 ( .A(n9457), .B(n9321), .Y(n9452) );
  INVX1 U9814 ( .A(G21744), .Y(n9457) );
  NAND2X1 U9815 ( .A(n9324), .B(G21776), .Y(n9450) );
  NAND2X1 U9816 ( .A(n7190), .B(n9325), .Y(n9449) );
  NAND2X1 U9817 ( .A(n9326), .B(n7188), .Y(n9448) );
  NAND4X1 U9818 ( .A(n9458), .B(n9459), .C(n9460), .D(n9461), .Y(G1165) );
  NOR4X1 U9819 ( .A(n9441), .B(n9462), .C(n9463), .D(n9464), .Y(n9461) );
  NOR2X1 U9820 ( .A(n9322), .B(n9465), .Y(n9464) );
  NOR2X1 U9821 ( .A(n9466), .B(n9319), .Y(n9463) );
  NOR2X1 U9822 ( .A(n9467), .B(n9321), .Y(n9462) );
  INVX1 U9823 ( .A(G21743), .Y(n9467) );
  NAND2X1 U9824 ( .A(n9324), .B(G21775), .Y(n9460) );
  NAND2X1 U9825 ( .A(n7203), .B(n9325), .Y(n9459) );
  NAND2X1 U9826 ( .A(n9326), .B(n7201), .Y(n9458) );
  NAND4X1 U9827 ( .A(n9468), .B(n9469), .C(n9470), .D(n9471), .Y(G1164) );
  NOR4X1 U9828 ( .A(n9441), .B(n9472), .C(n9473), .D(n9474), .Y(n9471) );
  NOR2X1 U9829 ( .A(n9322), .B(n9475), .Y(n9474) );
  NOR2X1 U9830 ( .A(n9476), .B(n9319), .Y(n9473) );
  NOR2X1 U9831 ( .A(n9477), .B(n9321), .Y(n9472) );
  INVX1 U9832 ( .A(G21742), .Y(n9477) );
  NAND2X1 U9833 ( .A(n9324), .B(G21774), .Y(n9470) );
  NAND2X1 U9834 ( .A(n7216), .B(n9325), .Y(n9469) );
  NAND2X1 U9835 ( .A(n9326), .B(n7214), .Y(n9468) );
  NAND4X1 U9836 ( .A(n9478), .B(n9479), .C(n9480), .D(n9481), .Y(G1163) );
  NOR4X1 U9837 ( .A(n9441), .B(n9482), .C(n9483), .D(n9484), .Y(n9481) );
  NOR2X1 U9838 ( .A(n9322), .B(n9485), .Y(n9484) );
  NOR2X1 U9839 ( .A(n9486), .B(n9319), .Y(n9483) );
  NOR2X1 U9840 ( .A(n9487), .B(n9321), .Y(n9482) );
  INVX1 U9841 ( .A(G21741), .Y(n9487) );
  NAND2X1 U9842 ( .A(n9324), .B(G21773), .Y(n9480) );
  NAND2X1 U9843 ( .A(n7233), .B(n9325), .Y(n9479) );
  NAND2X1 U9844 ( .A(n9326), .B(n7231), .Y(n9478) );
  NAND4X1 U9845 ( .A(n9488), .B(n9489), .C(n9490), .D(n9491), .Y(G1162) );
  NOR4X1 U9846 ( .A(n9441), .B(n9492), .C(n9493), .D(n9494), .Y(n9491) );
  NOR2X1 U9847 ( .A(n9322), .B(n9495), .Y(n9494) );
  NOR2X1 U9848 ( .A(n9496), .B(n9319), .Y(n9493) );
  NOR2X1 U9849 ( .A(n9497), .B(n9321), .Y(n9492) );
  INVX1 U9850 ( .A(G21740), .Y(n9497) );
  NAND2X1 U9851 ( .A(n9324), .B(G21772), .Y(n9490) );
  NAND2X1 U9852 ( .A(n7246), .B(n9325), .Y(n9489) );
  NAND2X1 U9853 ( .A(n9326), .B(n7244), .Y(n9488) );
  NAND4X1 U9854 ( .A(n9498), .B(n9499), .C(n9500), .D(n9501), .Y(G1161) );
  NOR4X1 U9855 ( .A(n9441), .B(n9502), .C(n9503), .D(n9504), .Y(n9501) );
  NOR2X1 U9856 ( .A(n9322), .B(n9505), .Y(n9504) );
  NOR2X1 U9857 ( .A(n9506), .B(n9319), .Y(n9503) );
  NOR2X1 U9858 ( .A(n9507), .B(n9321), .Y(n9502) );
  INVX1 U9859 ( .A(G21739), .Y(n9507) );
  NAND2X1 U9860 ( .A(n9324), .B(G21771), .Y(n9500) );
  NAND2X1 U9861 ( .A(n7263), .B(n9325), .Y(n9499) );
  NAND2X1 U9862 ( .A(n9326), .B(n7261), .Y(n9498) );
  NAND4X1 U9863 ( .A(n9508), .B(n9509), .C(n9510), .D(n9511), .Y(G1160) );
  NOR4X1 U9864 ( .A(n9441), .B(n9512), .C(n9513), .D(n9514), .Y(n9511) );
  NOR2X1 U9865 ( .A(n9322), .B(n9515), .Y(n9514) );
  NOR2X1 U9866 ( .A(n9516), .B(n9319), .Y(n9513) );
  NOR2X1 U9867 ( .A(n9517), .B(n9321), .Y(n9512) );
  INVX1 U9868 ( .A(G21738), .Y(n9517) );
  NAND2X1 U9869 ( .A(n9324), .B(G21770), .Y(n9510) );
  NAND2X1 U9870 ( .A(n7275), .B(n9325), .Y(n9509) );
  NAND2X1 U9871 ( .A(n9326), .B(n7273), .Y(n9508) );
  NAND4X1 U9872 ( .A(n9518), .B(n9519), .C(n9520), .D(n9521), .Y(G1159) );
  NOR4X1 U9873 ( .A(n9441), .B(n9522), .C(n9523), .D(n9524), .Y(n9521) );
  NOR2X1 U9874 ( .A(n9322), .B(n9525), .Y(n9524) );
  NOR2X1 U9875 ( .A(n9526), .B(n9319), .Y(n9523) );
  NOR2X1 U9876 ( .A(n9527), .B(n9321), .Y(n9522) );
  INVX1 U9877 ( .A(G21737), .Y(n9527) );
  NAND2X1 U9878 ( .A(n9324), .B(G21769), .Y(n9520) );
  NAND2X1 U9879 ( .A(n7291), .B(n9325), .Y(n9519) );
  NAND2X1 U9880 ( .A(n9326), .B(n7289), .Y(n9518) );
  NAND4X1 U9881 ( .A(n9528), .B(n9529), .C(n9530), .D(n9531), .Y(G1158) );
  NOR4X1 U9882 ( .A(n9441), .B(n9532), .C(n9533), .D(n9534), .Y(n9531) );
  NOR2X1 U9883 ( .A(n9322), .B(n6886), .Y(n9534) );
  NOR2X1 U9884 ( .A(n6892), .B(n9319), .Y(n9533) );
  INVX1 U9885 ( .A(G21609), .Y(n6892) );
  NOR2X1 U9886 ( .A(n9535), .B(n9321), .Y(n9532) );
  INVX1 U9887 ( .A(G21736), .Y(n9535) );
  NAND2X1 U9888 ( .A(n9324), .B(G21768), .Y(n9530) );
  NAND2X1 U9889 ( .A(n9325), .B(n6883), .Y(n9529) );
  NAND2X1 U9890 ( .A(n9326), .B(n9536), .Y(n9528) );
  NAND4X1 U9891 ( .A(n9537), .B(n9538), .C(n9539), .D(n9540), .Y(G1157) );
  NOR2X1 U9892 ( .A(n9322), .B(n7310), .Y(n9543) );
  NOR2X1 U9893 ( .A(n6899), .B(n9319), .Y(n9542) );
  NOR2X1 U9894 ( .A(n9544), .B(n9321), .Y(n9541) );
  INVX1 U9895 ( .A(G21735), .Y(n9544) );
  NAND2X1 U9896 ( .A(n9324), .B(G21767), .Y(n9539) );
  NAND2X1 U9897 ( .A(n6902), .B(n9325), .Y(n9538) );
  NAND2X1 U9898 ( .A(n9326), .B(n6904), .Y(n9537) );
  NAND4X1 U9899 ( .A(n9545), .B(n9546), .C(n9547), .D(n9548), .Y(G1156) );
  NOR2X1 U9900 ( .A(n9322), .B(n9552), .Y(n9551) );
  NOR2X1 U9901 ( .A(n6913), .B(n9319), .Y(n9550) );
  INVX1 U9902 ( .A(G21607), .Y(n6913) );
  NOR2X1 U9903 ( .A(n9553), .B(n9321), .Y(n9549) );
  INVX1 U9904 ( .A(G21734), .Y(n9553) );
  NAND2X1 U9905 ( .A(n9324), .B(G21766), .Y(n9547) );
  NAND2X1 U9906 ( .A(n6915), .B(n9325), .Y(n9546) );
  NAND2X1 U9907 ( .A(n9326), .B(n6916), .Y(n9545) );
  NAND4X1 U9908 ( .A(n9554), .B(n9555), .C(n9556), .D(n9557), .Y(G1155) );
  NOR2X1 U9909 ( .A(n9322), .B(n9561), .Y(n9560) );
  INVX1 U9910 ( .A(n6928), .Y(n9561) );
  NOR2X1 U9911 ( .A(n6924), .B(n9319), .Y(n9559) );
  INVX1 U9912 ( .A(G21606), .Y(n6924) );
  NOR2X1 U9913 ( .A(n9562), .B(n9321), .Y(n9558) );
  INVX1 U9914 ( .A(G21733), .Y(n9562) );
  NAND2X1 U9915 ( .A(n9324), .B(G21765), .Y(n9556) );
  NAND2X1 U9916 ( .A(n6926), .B(n9325), .Y(n9555) );
  NAND2X1 U9917 ( .A(n9326), .B(n6927), .Y(n9554) );
  NAND4X1 U9918 ( .A(n9563), .B(n9564), .C(n9565), .D(n9566), .Y(G1154) );
  NOR4X1 U9919 ( .A(n9441), .B(n9567), .C(n9568), .D(n9569), .Y(n9566) );
  NOR2X1 U9920 ( .A(n9322), .B(n9570), .Y(n9569) );
  NOR2X1 U9921 ( .A(n6935), .B(n9319), .Y(n9568) );
  INVX1 U9922 ( .A(G21605), .Y(n6935) );
  NOR2X1 U9923 ( .A(n9571), .B(n9321), .Y(n9567) );
  INVX1 U9924 ( .A(G21732), .Y(n9571) );
  NAND2X1 U9925 ( .A(n9324), .B(G21764), .Y(n9565) );
  NAND2X1 U9926 ( .A(n6937), .B(n9325), .Y(n9564) );
  NAND2X1 U9927 ( .A(n9326), .B(n6938), .Y(n9563) );
  NAND4X1 U9928 ( .A(n9572), .B(n9573), .C(n9574), .D(n9575), .Y(G1153) );
  NOR4X1 U9929 ( .A(n9441), .B(n9576), .C(n9577), .D(n9578), .Y(n9575) );
  NOR2X1 U9930 ( .A(n9579), .B(n9580), .Y(n9578) );
  INVX1 U9931 ( .A(n6950), .Y(n9580) );
  NOR2X1 U9932 ( .A(n6946), .B(n9319), .Y(n9577) );
  INVX1 U9933 ( .A(G21604), .Y(n6946) );
  NOR2X1 U9934 ( .A(n9581), .B(n9321), .Y(n9576) );
  INVX1 U9935 ( .A(G21731), .Y(n9581) );
  NAND2X1 U9936 ( .A(n9324), .B(G21763), .Y(n9574) );
  NAND2X1 U9937 ( .A(n6948), .B(n9325), .Y(n9573) );
  NAND2X1 U9938 ( .A(n6949), .B(n9582), .Y(n9572) );
  NAND4X1 U9939 ( .A(n9583), .B(n9584), .C(n9585), .D(n9586), .Y(G1152) );
  NOR4X1 U9940 ( .A(n9441), .B(n9587), .C(n9588), .D(n9589), .Y(n9586) );
  NOR2X1 U9941 ( .A(n9579), .B(n8847), .Y(n9589) );
  INVX1 U9942 ( .A(n6961), .Y(n8847) );
  NOR2X1 U9943 ( .A(n6957), .B(n9319), .Y(n9588) );
  NOR2X1 U9944 ( .A(n9590), .B(n9321), .Y(n9587) );
  INVX1 U9945 ( .A(G21730), .Y(n9590) );
  NOR3X1 U9946 ( .A(G21427), .B(G21428), .C(n9324), .Y(n9441) );
  NAND2X1 U9947 ( .A(n9324), .B(G21762), .Y(n9585) );
  NAND2X1 U9948 ( .A(n6959), .B(n9325), .Y(n9584) );
  NAND2X1 U9949 ( .A(n6960), .B(n9582), .Y(n9583) );
  NAND4X1 U9950 ( .A(n9591), .B(n9592), .C(n9593), .D(n9594), .Y(G1151) );
  NOR3X1 U9951 ( .A(n9595), .B(n9596), .C(n9597), .Y(n9594) );
  NOR2X1 U9952 ( .A(n6968), .B(n9319), .Y(n9597) );
  NOR2X1 U9953 ( .A(n9598), .B(n9321), .Y(n9596) );
  NOR2X1 U9954 ( .A(n9579), .B(n7379), .Y(n9595) );
  NAND2X1 U9955 ( .A(n9324), .B(G21761), .Y(n9593) );
  NAND2X1 U9956 ( .A(n6969), .B(n9325), .Y(n9592) );
  NAND2X1 U9957 ( .A(n6970), .B(n9582), .Y(n9591) );
  NAND4X1 U9958 ( .A(n9599), .B(n9600), .C(n9601), .D(n9602), .Y(G1150) );
  NOR3X1 U9959 ( .A(n9603), .B(n9604), .C(n9605), .Y(n9602) );
  NOR2X1 U9960 ( .A(n6978), .B(n9319), .Y(n9605) );
  NOR2X1 U9961 ( .A(n9606), .B(n9321), .Y(n9604) );
  NOR2X1 U9962 ( .A(n7387), .B(n9579), .Y(n9603) );
  NAND2X1 U9963 ( .A(n9324), .B(G21760), .Y(n9601) );
  NAND2X1 U9964 ( .A(n6979), .B(n9325), .Y(n9600) );
  NAND2X1 U9965 ( .A(n6980), .B(n9582), .Y(n9599) );
  NAND4X1 U9966 ( .A(n9607), .B(n9608), .C(n9609), .D(n9610), .Y(G1149) );
  NOR3X1 U9967 ( .A(n9611), .B(n9612), .C(n9613), .Y(n9610) );
  NOR2X1 U9968 ( .A(n6988), .B(n9319), .Y(n9613) );
  NOR2X1 U9969 ( .A(n9614), .B(n9321), .Y(n9612) );
  NOR2X1 U9970 ( .A(n9579), .B(n9615), .Y(n9611) );
  NAND2X1 U9971 ( .A(n9324), .B(G21759), .Y(n9609) );
  NAND2X1 U9972 ( .A(n6990), .B(n9325), .Y(n9608) );
  NAND2X1 U9973 ( .A(n6991), .B(n9582), .Y(n9607) );
  NAND4X1 U9974 ( .A(n9616), .B(n9617), .C(n9618), .D(n9619), .Y(G1148) );
  NOR3X1 U9975 ( .A(n9620), .B(n9621), .C(n9622), .Y(n9619) );
  NOR2X1 U9976 ( .A(n6999), .B(n9319), .Y(n9622) );
  NOR2X1 U9977 ( .A(n9624), .B(n9321), .Y(n9621) );
  NAND2X1 U9978 ( .A(n9627), .B(n9628), .Y(n9626) );
  NAND3X1 U9979 ( .A(n9629), .B(n9630), .C(n9631), .Y(n9628) );
  OR2X1 U9980 ( .A(n9632), .B(n8895), .Y(n9627) );
  NOR2X1 U9981 ( .A(n9579), .B(n7410), .Y(n9620) );
  AND2X1 U9982 ( .A(n9322), .B(n9633), .Y(n9579) );
  NAND3X1 U9983 ( .A(n8772), .B(n7444), .C(n9625), .Y(n9633) );
  AND2X1 U9984 ( .A(n9634), .B(n9635), .Y(n9322) );
  NAND3X1 U9985 ( .A(n9636), .B(n9631), .C(n9625), .Y(n9635) );
  NAND3X1 U9986 ( .A(G21427), .B(n9623), .C(n7025), .Y(n9634) );
  NAND2X1 U9987 ( .A(n9324), .B(G21758), .Y(n9618) );
  NAND2X1 U9988 ( .A(n7001), .B(n9325), .Y(n9617) );
  NAND4X1 U9989 ( .A(n9625), .B(n9631), .C(n9639), .D(n9630), .Y(n9638) );
  INVX1 U9990 ( .A(n9629), .Y(n9639) );
  NAND3X1 U9991 ( .A(n9640), .B(n9623), .C(G21427), .Y(n9637) );
  NAND2X1 U9992 ( .A(n7002), .B(n9582), .Y(n9616) );
  OR2X1 U9993 ( .A(n9326), .B(n9641), .Y(n9582) );
  NOR3X1 U9994 ( .A(n9324), .B(n7442), .C(n9642), .Y(n9641) );
  AND3X1 U9995 ( .A(n8895), .B(n9203), .C(n9625), .Y(n9326) );
  NOR2X1 U9996 ( .A(n7430), .B(n9324), .Y(n9625) );
  NAND4X1 U9997 ( .A(n9069), .B(n7431), .C(n8821), .D(n8805), .Y(n9623) );
  NAND3X1 U9998 ( .A(G21425), .B(G21428), .C(n8798), .Y(n8805) );
  NAND3X1 U9999 ( .A(n7430), .B(n8817), .C(n7564), .Y(n8821) );
  NAND2X1 U10000 ( .A(n9058), .B(n8817), .Y(n7431) );
  NOR2X1 U10001 ( .A(n8783), .B(G21425), .Y(n9058) );
  INVX1 U10002 ( .A(n9057), .Y(n9069) );
  NAND3X1 U10003 ( .A(n9643), .B(n9644), .C(n9645), .Y(n9057) );
  OR2X1 U10004 ( .A(n9263), .B(n9092), .Y(n9645) );
  NAND3X1 U10005 ( .A(n9053), .B(n9646), .C(n9647), .Y(n9263) );
  NAND3X1 U10006 ( .A(n9260), .B(n7441), .C(n8818), .Y(n9643) );
  NOR2X1 U10007 ( .A(n9630), .B(n9274), .Y(n8895) );
  INVX1 U10008 ( .A(n7454), .Y(n9274) );
  INVX1 U10009 ( .A(n9636), .Y(n9630) );
  NOR2X1 U10010 ( .A(G35), .B(G21797), .Y(n9636) );
  NAND2X1 U10011 ( .A(n9648), .B(n9649), .Y(G1147) );
  NAND2X1 U10012 ( .A(n9650), .B(n7025), .Y(n9649) );
  NAND2X1 U10013 ( .A(G21757), .B(n9651), .Y(n9648) );
  NAND3X1 U10014 ( .A(n9652), .B(n9653), .C(n9654), .Y(G1146) );
  NAND2X1 U10015 ( .A(G21756), .B(n9651), .Y(n9654) );
  NAND2X1 U10016 ( .A(n9650), .B(n7039), .Y(n9653) );
  NAND2X1 U10017 ( .A(n9655), .B(n7038), .Y(n9652) );
  NAND3X1 U10018 ( .A(n9656), .B(n9657), .C(n9658), .Y(G1145) );
  NAND2X1 U10019 ( .A(G21755), .B(n9651), .Y(n9658) );
  NAND2X1 U10020 ( .A(n9650), .B(n9346), .Y(n9657) );
  NAND2X1 U10021 ( .A(n9655), .B(n9659), .Y(n9656) );
  NAND3X1 U10022 ( .A(n9660), .B(n9661), .C(n9662), .Y(G1144) );
  NAND2X1 U10023 ( .A(G21754), .B(n9651), .Y(n9662) );
  NAND2X1 U10024 ( .A(n9650), .B(n7067), .Y(n9661) );
  NAND2X1 U10025 ( .A(n9655), .B(n7066), .Y(n9660) );
  NAND3X1 U10026 ( .A(n9663), .B(n9664), .C(n9665), .Y(G1143) );
  NAND2X1 U10027 ( .A(G21753), .B(n9651), .Y(n9665) );
  NAND2X1 U10028 ( .A(n9650), .B(n9366), .Y(n9664) );
  NAND2X1 U10029 ( .A(n9655), .B(n9666), .Y(n9663) );
  NAND3X1 U10030 ( .A(n9667), .B(n9668), .C(n9669), .Y(G1142) );
  NAND2X1 U10031 ( .A(G21752), .B(n9651), .Y(n9669) );
  NAND2X1 U10032 ( .A(n9650), .B(n9376), .Y(n9668) );
  NAND2X1 U10033 ( .A(n9655), .B(n9670), .Y(n9667) );
  NAND3X1 U10034 ( .A(n9671), .B(n9672), .C(n9673), .Y(G1141) );
  NAND2X1 U10035 ( .A(G21751), .B(n9651), .Y(n9673) );
  NAND2X1 U10036 ( .A(n9650), .B(n7104), .Y(n9672) );
  NAND2X1 U10037 ( .A(n9655), .B(n7103), .Y(n9671) );
  NAND3X1 U10038 ( .A(n9674), .B(n9675), .C(n9676), .Y(G1140) );
  NAND2X1 U10039 ( .A(G21750), .B(n9651), .Y(n9676) );
  NAND2X1 U10040 ( .A(n9650), .B(n9396), .Y(n9675) );
  NAND2X1 U10041 ( .A(n9655), .B(n9677), .Y(n9674) );
  NAND3X1 U10042 ( .A(n9678), .B(n9679), .C(n9680), .Y(G1139) );
  NAND2X1 U10043 ( .A(G21749), .B(n9651), .Y(n9680) );
  NAND2X1 U10044 ( .A(n9650), .B(n7127), .Y(n9679) );
  NAND2X1 U10045 ( .A(n9655), .B(n7126), .Y(n9678) );
  NAND3X1 U10046 ( .A(n9681), .B(n9682), .C(n9683), .Y(G1138) );
  NAND2X1 U10047 ( .A(G21748), .B(n9651), .Y(n9683) );
  NAND2X1 U10048 ( .A(n9650), .B(n7140), .Y(n9682) );
  NAND2X1 U10049 ( .A(n9655), .B(n7139), .Y(n9681) );
  NAND3X1 U10050 ( .A(n9684), .B(n9685), .C(n9686), .Y(G1137) );
  NAND2X1 U10051 ( .A(G21747), .B(n9651), .Y(n9686) );
  NAND2X1 U10052 ( .A(n9650), .B(n7153), .Y(n9685) );
  NAND2X1 U10053 ( .A(n9655), .B(n7152), .Y(n9684) );
  NAND3X1 U10054 ( .A(n9687), .B(n9688), .C(n9689), .Y(G1136) );
  NAND2X1 U10055 ( .A(G21746), .B(n9651), .Y(n9689) );
  NAND2X1 U10056 ( .A(n9650), .B(n7165), .Y(n9688) );
  NAND2X1 U10057 ( .A(n9655), .B(n7164), .Y(n9687) );
  NAND3X1 U10058 ( .A(n9690), .B(n9691), .C(n9692), .Y(G1135) );
  NAND2X1 U10059 ( .A(G21745), .B(n9651), .Y(n9692) );
  NAND2X1 U10060 ( .A(n9650), .B(n7178), .Y(n9691) );
  NAND2X1 U10061 ( .A(n9655), .B(n7177), .Y(n9690) );
  NAND3X1 U10062 ( .A(n9693), .B(n9694), .C(n9695), .Y(G1134) );
  NAND2X1 U10063 ( .A(G21744), .B(n9651), .Y(n9695) );
  NAND2X1 U10064 ( .A(n9650), .B(n7190), .Y(n9694) );
  NAND2X1 U10065 ( .A(n9655), .B(n7189), .Y(n9693) );
  NAND3X1 U10066 ( .A(n9696), .B(n9697), .C(n9698), .Y(G1133) );
  NAND2X1 U10067 ( .A(G21743), .B(n9651), .Y(n9698) );
  NAND2X1 U10068 ( .A(n9650), .B(n7203), .Y(n9697) );
  NAND2X1 U10069 ( .A(n9655), .B(n7202), .Y(n9696) );
  NAND3X1 U10070 ( .A(n9699), .B(n9700), .C(n9701), .Y(G1132) );
  NAND2X1 U10071 ( .A(G21742), .B(n9651), .Y(n9701) );
  NAND2X1 U10072 ( .A(n9650), .B(n7216), .Y(n9700) );
  NAND2X1 U10073 ( .A(n9655), .B(n7215), .Y(n9699) );
  NAND3X1 U10074 ( .A(n9702), .B(n9703), .C(n9704), .Y(G1131) );
  NAND2X1 U10075 ( .A(G21741), .B(n9651), .Y(n9704) );
  NAND2X1 U10076 ( .A(n9650), .B(n7233), .Y(n9703) );
  NAND2X1 U10077 ( .A(n9655), .B(n7232), .Y(n9702) );
  NAND3X1 U10078 ( .A(n9705), .B(n9706), .C(n9707), .Y(G1130) );
  NAND2X1 U10079 ( .A(G21740), .B(n9651), .Y(n9707) );
  NAND2X1 U10080 ( .A(n9650), .B(n7246), .Y(n9706) );
  NAND2X1 U10081 ( .A(n9655), .B(n7245), .Y(n9705) );
  NAND3X1 U10082 ( .A(n9708), .B(n9709), .C(n9710), .Y(G1129) );
  NAND2X1 U10083 ( .A(G21739), .B(n9651), .Y(n9710) );
  NAND2X1 U10084 ( .A(n9650), .B(n7263), .Y(n9709) );
  NAND2X1 U10085 ( .A(n9655), .B(n7262), .Y(n9708) );
  NAND3X1 U10086 ( .A(n9711), .B(n9712), .C(n9713), .Y(G1128) );
  NAND2X1 U10087 ( .A(G21738), .B(n9651), .Y(n9713) );
  NAND2X1 U10088 ( .A(n9650), .B(n7275), .Y(n9712) );
  NAND2X1 U10089 ( .A(n9655), .B(n7274), .Y(n9711) );
  NAND3X1 U10090 ( .A(n9714), .B(n9715), .C(n9716), .Y(G1127) );
  NAND2X1 U10091 ( .A(G21737), .B(n9651), .Y(n9716) );
  NAND2X1 U10092 ( .A(n9650), .B(n7291), .Y(n9715) );
  NAND2X1 U10093 ( .A(n9655), .B(n7290), .Y(n9714) );
  NAND3X1 U10094 ( .A(n9717), .B(n9718), .C(n9719), .Y(G1126) );
  NAND2X1 U10095 ( .A(G21736), .B(n9651), .Y(n9719) );
  NAND2X1 U10096 ( .A(n9650), .B(n6883), .Y(n9718) );
  NAND2X1 U10097 ( .A(n9655), .B(n9720), .Y(n9717) );
  NAND3X1 U10098 ( .A(n9721), .B(n9722), .C(n9723), .Y(G1125) );
  NAND2X1 U10099 ( .A(G21735), .B(n9651), .Y(n9723) );
  NAND2X1 U10100 ( .A(n9650), .B(n6902), .Y(n9722) );
  NAND2X1 U10101 ( .A(n9655), .B(n6906), .Y(n9721) );
  NAND3X1 U10102 ( .A(n9724), .B(n9725), .C(n9726), .Y(G1124) );
  NAND2X1 U10103 ( .A(G21734), .B(n9651), .Y(n9726) );
  NAND2X1 U10104 ( .A(n9650), .B(n6915), .Y(n9725) );
  NAND2X1 U10105 ( .A(n9655), .B(n6917), .Y(n9724) );
  NAND3X1 U10106 ( .A(n9727), .B(n9728), .C(n9729), .Y(G1123) );
  NAND2X1 U10107 ( .A(G21733), .B(n9651), .Y(n9729) );
  NAND2X1 U10108 ( .A(n9650), .B(n6926), .Y(n9728) );
  NAND2X1 U10109 ( .A(n9655), .B(n6928), .Y(n9727) );
  NAND3X1 U10110 ( .A(n9730), .B(n9731), .C(n9732), .Y(G1122) );
  NAND2X1 U10111 ( .A(G21732), .B(n9651), .Y(n9732) );
  NAND2X1 U10112 ( .A(n9650), .B(n6937), .Y(n9731) );
  NAND2X1 U10113 ( .A(n9655), .B(n6939), .Y(n9730) );
  NAND3X1 U10114 ( .A(n9733), .B(n9734), .C(n9735), .Y(G1121) );
  NAND2X1 U10115 ( .A(G21731), .B(n9651), .Y(n9735) );
  NAND2X1 U10116 ( .A(n9650), .B(n6948), .Y(n9734) );
  NAND2X1 U10117 ( .A(n9655), .B(n6950), .Y(n9733) );
  NAND3X1 U10118 ( .A(n9736), .B(n9737), .C(n9738), .Y(G1120) );
  NAND2X1 U10119 ( .A(G21730), .B(n9651), .Y(n9738) );
  NAND2X1 U10120 ( .A(n9650), .B(n6959), .Y(n9737) );
  NAND2X1 U10121 ( .A(n9655), .B(n6961), .Y(n9736) );
  NAND3X1 U10122 ( .A(n9739), .B(n9740), .C(n9741), .Y(G1119) );
  NAND2X1 U10123 ( .A(G21729), .B(n9651), .Y(n9741) );
  NAND2X1 U10124 ( .A(n9650), .B(n6969), .Y(n9740) );
  NAND2X1 U10125 ( .A(n9655), .B(n6971), .Y(n9739) );
  NAND3X1 U10126 ( .A(n9742), .B(n9743), .C(n9744), .Y(G1118) );
  NAND2X1 U10127 ( .A(G21728), .B(n9651), .Y(n9744) );
  NAND2X1 U10128 ( .A(n9650), .B(n6979), .Y(n9743) );
  NAND2X1 U10129 ( .A(n9655), .B(n6981), .Y(n9742) );
  NAND3X1 U10130 ( .A(n9745), .B(n9746), .C(n9747), .Y(G1117) );
  NAND2X1 U10131 ( .A(G21727), .B(n9651), .Y(n9747) );
  NAND2X1 U10132 ( .A(n9650), .B(n6990), .Y(n9746) );
  NAND2X1 U10133 ( .A(n9655), .B(n6992), .Y(n9745) );
  NAND3X1 U10134 ( .A(n9748), .B(n9749), .C(n9750), .Y(G1116) );
  NAND2X1 U10135 ( .A(G21726), .B(n9651), .Y(n9750) );
  NAND2X1 U10136 ( .A(n9650), .B(n7001), .Y(n9749) );
  NAND2X1 U10137 ( .A(n9655), .B(n7003), .Y(n9748) );
  NAND2X1 U10138 ( .A(n9753), .B(n9754), .Y(n9752) );
  NAND2X1 U10139 ( .A(n9755), .B(n7457), .Y(n9754) );
  NAND3X1 U10140 ( .A(n9756), .B(n9757), .C(n9758), .Y(G1115) );
  NAND2X1 U10141 ( .A(G21725), .B(n9759), .Y(n9758) );
  NAND2X1 U10142 ( .A(n9760), .B(G1), .Y(n9757) );
  NAND2X1 U10143 ( .A(n9761), .B(n7025), .Y(n9756) );
  NAND3X1 U10144 ( .A(n9762), .B(n9763), .C(n9764), .Y(G1114) );
  NOR3X1 U10145 ( .A(n9765), .B(n9766), .C(n9767), .Y(n9764) );
  AND2X1 U10146 ( .A(G2), .B(n9760), .Y(n9767) );
  NOR2X1 U10147 ( .A(n9768), .B(n9769), .Y(n9766) );
  INVX1 U10148 ( .A(G18), .Y(n9769) );
  NOR2X1 U10149 ( .A(n9770), .B(n9771), .Y(n9765) );
  NAND2X1 U10150 ( .A(n9772), .B(n7037), .Y(n9763) );
  NAND2X1 U10151 ( .A(G21724), .B(n9759), .Y(n9762) );
  NAND3X1 U10152 ( .A(n9773), .B(n9774), .C(n9775), .Y(G1113) );
  NOR3X1 U10153 ( .A(n9776), .B(n9777), .C(n9778), .Y(n9775) );
  AND2X1 U10154 ( .A(G3), .B(n9760), .Y(n9778) );
  NOR2X1 U10155 ( .A(n9768), .B(n9779), .Y(n9777) );
  INVX1 U10156 ( .A(G19), .Y(n9779) );
  NOR2X1 U10157 ( .A(n7051), .B(n9771), .Y(n9776) );
  INVX1 U10158 ( .A(n9346), .Y(n7051) );
  NAND2X1 U10159 ( .A(n9772), .B(n7053), .Y(n9774) );
  NAND2X1 U10160 ( .A(G21723), .B(n9759), .Y(n9773) );
  NAND3X1 U10161 ( .A(n9780), .B(n9781), .C(n9782), .Y(G1112) );
  NOR3X1 U10162 ( .A(n9783), .B(n9784), .C(n9785), .Y(n9782) );
  AND2X1 U10163 ( .A(G4), .B(n9760), .Y(n9785) );
  NOR2X1 U10164 ( .A(n9768), .B(n9786), .Y(n9784) );
  INVX1 U10165 ( .A(G20), .Y(n9786) );
  NOR2X1 U10166 ( .A(n9787), .B(n9771), .Y(n9783) );
  NAND2X1 U10167 ( .A(n9772), .B(n7065), .Y(n9781) );
  NAND2X1 U10168 ( .A(G21722), .B(n9759), .Y(n9780) );
  NAND3X1 U10169 ( .A(n9788), .B(n9789), .C(n9790), .Y(G1111) );
  NOR3X1 U10170 ( .A(n9791), .B(n9792), .C(n9793), .Y(n9790) );
  AND2X1 U10171 ( .A(G5), .B(n9760), .Y(n9793) );
  NOR2X1 U10172 ( .A(n9768), .B(n9794), .Y(n9792) );
  INVX1 U10173 ( .A(G21), .Y(n9794) );
  NOR2X1 U10174 ( .A(n7078), .B(n9771), .Y(n9791) );
  INVX1 U10175 ( .A(n9366), .Y(n7078) );
  NAND2X1 U10176 ( .A(n9772), .B(n7079), .Y(n9789) );
  NAND2X1 U10177 ( .A(G21721), .B(n9759), .Y(n9788) );
  NAND3X1 U10178 ( .A(n9795), .B(n9796), .C(n9797), .Y(G1110) );
  NOR3X1 U10179 ( .A(n9798), .B(n9799), .C(n9800), .Y(n9797) );
  AND2X1 U10180 ( .A(G6), .B(n9760), .Y(n9800) );
  NOR2X1 U10181 ( .A(n9768), .B(n9801), .Y(n9799) );
  INVX1 U10182 ( .A(G22), .Y(n9801) );
  NOR2X1 U10183 ( .A(n7090), .B(n9771), .Y(n9798) );
  NAND2X1 U10184 ( .A(n9772), .B(n7091), .Y(n9796) );
  NAND2X1 U10185 ( .A(G21720), .B(n9759), .Y(n9795) );
  NAND3X1 U10186 ( .A(n9802), .B(n9803), .C(n9804), .Y(G1109) );
  NOR3X1 U10187 ( .A(n9805), .B(n9806), .C(n9807), .Y(n9804) );
  AND2X1 U10188 ( .A(G7), .B(n9760), .Y(n9807) );
  NOR2X1 U10189 ( .A(n9768), .B(n9808), .Y(n9806) );
  INVX1 U10190 ( .A(G23), .Y(n9808) );
  AND2X1 U10191 ( .A(n7104), .B(n9761), .Y(n9805) );
  NAND2X1 U10192 ( .A(n9772), .B(n7102), .Y(n9803) );
  NAND2X1 U10193 ( .A(G21719), .B(n9759), .Y(n9802) );
  NAND3X1 U10194 ( .A(n9809), .B(n9810), .C(n9811), .Y(G1108) );
  NOR3X1 U10195 ( .A(n9812), .B(n9813), .C(n9814), .Y(n9811) );
  AND2X1 U10196 ( .A(G8), .B(n9760), .Y(n9814) );
  NOR2X1 U10197 ( .A(n9768), .B(n9815), .Y(n9813) );
  INVX1 U10198 ( .A(G24), .Y(n9815) );
  NOR2X1 U10199 ( .A(n7114), .B(n9771), .Y(n9812) );
  NAND2X1 U10200 ( .A(n9772), .B(n7115), .Y(n9810) );
  NAND2X1 U10201 ( .A(G21718), .B(n9759), .Y(n9809) );
  NAND3X1 U10202 ( .A(n9816), .B(n9817), .C(n9818), .Y(G1107) );
  NOR3X1 U10203 ( .A(n9819), .B(n9820), .C(n9821), .Y(n9818) );
  AND2X1 U10204 ( .A(G9), .B(n9760), .Y(n9821) );
  NOR2X1 U10205 ( .A(n9822), .B(n9768), .Y(n9820) );
  INVX1 U10206 ( .A(G25), .Y(n9822) );
  NOR2X1 U10207 ( .A(n9823), .B(n9771), .Y(n9819) );
  NAND2X1 U10208 ( .A(n9772), .B(n7125), .Y(n9817) );
  NAND2X1 U10209 ( .A(G21717), .B(n9759), .Y(n9816) );
  NAND3X1 U10210 ( .A(n9824), .B(n9825), .C(n9826), .Y(G1106) );
  NOR3X1 U10211 ( .A(n9827), .B(n9828), .C(n9829), .Y(n9826) );
  AND2X1 U10212 ( .A(G10), .B(n9760), .Y(n9829) );
  NOR2X1 U10213 ( .A(n9830), .B(n9768), .Y(n9828) );
  INVX1 U10214 ( .A(G26), .Y(n9830) );
  NOR2X1 U10215 ( .A(n9831), .B(n9771), .Y(n9827) );
  NAND2X1 U10216 ( .A(n9772), .B(n7138), .Y(n9825) );
  NAND2X1 U10217 ( .A(G21716), .B(n9759), .Y(n9824) );
  NAND3X1 U10218 ( .A(n9832), .B(n9833), .C(n9834), .Y(G1105) );
  NOR3X1 U10219 ( .A(n9835), .B(n9836), .C(n9837), .Y(n9834) );
  AND2X1 U10220 ( .A(G11), .B(n9760), .Y(n9837) );
  NOR2X1 U10221 ( .A(n9838), .B(n9768), .Y(n9836) );
  INVX1 U10222 ( .A(G27), .Y(n9838) );
  NOR2X1 U10223 ( .A(n9839), .B(n9771), .Y(n9835) );
  NAND2X1 U10224 ( .A(n9772), .B(n7151), .Y(n9833) );
  NAND2X1 U10225 ( .A(G21715), .B(n9759), .Y(n9832) );
  NAND3X1 U10226 ( .A(n9840), .B(n9841), .C(n9842), .Y(G1104) );
  NOR3X1 U10227 ( .A(n9843), .B(n9844), .C(n9845), .Y(n9842) );
  AND2X1 U10228 ( .A(G12), .B(n9760), .Y(n9845) );
  NOR2X1 U10229 ( .A(n9846), .B(n9768), .Y(n9844) );
  INVX1 U10230 ( .A(G28), .Y(n9846) );
  NOR2X1 U10231 ( .A(n9847), .B(n9771), .Y(n9843) );
  NAND2X1 U10232 ( .A(n9772), .B(n7163), .Y(n9841) );
  NAND2X1 U10233 ( .A(G21714), .B(n9759), .Y(n9840) );
  NAND3X1 U10234 ( .A(n9848), .B(n9849), .C(n9850), .Y(G1103) );
  NOR3X1 U10235 ( .A(n9851), .B(n9852), .C(n9853), .Y(n9850) );
  AND2X1 U10236 ( .A(G13), .B(n9760), .Y(n9853) );
  NOR2X1 U10237 ( .A(n9854), .B(n9768), .Y(n9852) );
  INVX1 U10238 ( .A(G29), .Y(n9854) );
  AND2X1 U10239 ( .A(n7178), .B(n9761), .Y(n9851) );
  NAND2X1 U10240 ( .A(n9772), .B(n7176), .Y(n9849) );
  NAND2X1 U10241 ( .A(G21713), .B(n9759), .Y(n9848) );
  NAND3X1 U10242 ( .A(n9855), .B(n9856), .C(n9857), .Y(G1102) );
  NOR3X1 U10243 ( .A(n9858), .B(n9859), .C(n9860), .Y(n9857) );
  AND2X1 U10244 ( .A(G14), .B(n9760), .Y(n9860) );
  NOR2X1 U10245 ( .A(n9861), .B(n9768), .Y(n9859) );
  INVX1 U10246 ( .A(G30), .Y(n9861) );
  NOR2X1 U10247 ( .A(n9862), .B(n9771), .Y(n9858) );
  NAND2X1 U10248 ( .A(n9772), .B(n7188), .Y(n9856) );
  NAND2X1 U10249 ( .A(G21712), .B(n9759), .Y(n9855) );
  NAND3X1 U10250 ( .A(n9863), .B(n9864), .C(n9865), .Y(G1101) );
  NOR3X1 U10251 ( .A(n9866), .B(n9867), .C(n9868), .Y(n9865) );
  AND2X1 U10252 ( .A(G15), .B(n9760), .Y(n9868) );
  NOR2X1 U10253 ( .A(n9869), .B(n9768), .Y(n9867) );
  INVX1 U10254 ( .A(G31), .Y(n9869) );
  NOR2X1 U10255 ( .A(n9870), .B(n9771), .Y(n9866) );
  NAND2X1 U10256 ( .A(n9772), .B(n7201), .Y(n9864) );
  NAND2X1 U10257 ( .A(G21711), .B(n9759), .Y(n9863) );
  NAND3X1 U10258 ( .A(n9871), .B(n9872), .C(n9873), .Y(G1100) );
  NOR3X1 U10259 ( .A(n9874), .B(n9875), .C(n9876), .Y(n9873) );
  AND2X1 U10260 ( .A(G16), .B(n9760), .Y(n9876) );
  NOR2X1 U10261 ( .A(n9759), .B(n7439), .Y(n9760) );
  NOR2X1 U10262 ( .A(n9877), .B(n9768), .Y(n9875) );
  OR2X1 U10263 ( .A(n9759), .B(n9076), .Y(n9768) );
  INVX1 U10264 ( .A(G32), .Y(n9877) );
  NOR2X1 U10265 ( .A(n9878), .B(n9771), .Y(n9874) );
  INVX1 U10266 ( .A(n9761), .Y(n9771) );
  NAND2X1 U10267 ( .A(n9772), .B(n7214), .Y(n9872) );
  NAND2X1 U10268 ( .A(G21710), .B(n9759), .Y(n9871) );
  NAND4X1 U10269 ( .A(n9879), .B(n9880), .C(n9881), .D(n9882), .Y(G1099) );
  NAND2X1 U10270 ( .A(n9761), .B(n7233), .Y(n9882) );
  NAND2X1 U10271 ( .A(n9772), .B(n7231), .Y(n9881) );
  NAND2X1 U10272 ( .A(G17), .B(n9883), .Y(n9880) );
  NAND2X1 U10273 ( .A(G21709), .B(n9759), .Y(n9879) );
  NAND4X1 U10274 ( .A(n9884), .B(n9885), .C(n9886), .D(n9887), .Y(G1098) );
  NAND2X1 U10275 ( .A(n9761), .B(n7246), .Y(n9887) );
  NAND2X1 U10276 ( .A(n9772), .B(n7244), .Y(n9886) );
  NAND2X1 U10277 ( .A(n9883), .B(G18), .Y(n9885) );
  NAND2X1 U10278 ( .A(G21708), .B(n9759), .Y(n9884) );
  NAND4X1 U10279 ( .A(n9888), .B(n9889), .C(n9890), .D(n9891), .Y(G1097) );
  NAND2X1 U10280 ( .A(n9761), .B(n7263), .Y(n9891) );
  NAND2X1 U10281 ( .A(n9772), .B(n7261), .Y(n9890) );
  NAND2X1 U10282 ( .A(n9883), .B(G19), .Y(n9889) );
  NAND2X1 U10283 ( .A(G21707), .B(n9759), .Y(n9888) );
  NAND4X1 U10284 ( .A(n9892), .B(n9893), .C(n9894), .D(n9895), .Y(G1096) );
  NAND2X1 U10285 ( .A(n9761), .B(n7275), .Y(n9895) );
  NAND2X1 U10286 ( .A(n9772), .B(n7273), .Y(n9894) );
  NAND2X1 U10287 ( .A(n9883), .B(G20), .Y(n9893) );
  NAND2X1 U10288 ( .A(G21706), .B(n9759), .Y(n9892) );
  NAND4X1 U10289 ( .A(n9896), .B(n9897), .C(n9898), .D(n9899), .Y(G1095) );
  NAND2X1 U10290 ( .A(n9761), .B(n7291), .Y(n9899) );
  NAND2X1 U10291 ( .A(n9772), .B(n7289), .Y(n9898) );
  NAND2X1 U10292 ( .A(n9883), .B(G21), .Y(n9897) );
  NAND2X1 U10293 ( .A(G21705), .B(n9759), .Y(n9896) );
  NAND4X1 U10294 ( .A(n9900), .B(n9901), .C(n9902), .D(n9903), .Y(G1094) );
  NAND2X1 U10295 ( .A(n9772), .B(n9536), .Y(n9903) );
  INVX1 U10296 ( .A(n6888), .Y(n9536) );
  NAND3X1 U10297 ( .A(n9904), .B(n9905), .C(n9906), .Y(n6888) );
  NAND2X1 U10298 ( .A(n9907), .B(n9908), .Y(n9906) );
  NAND2X1 U10299 ( .A(n9909), .B(n9910), .Y(n9907) );
  OR2X1 U10300 ( .A(n9911), .B(n9912), .Y(n9910) );
  NAND2X1 U10301 ( .A(n9913), .B(n9911), .Y(n9905) );
  OR2X1 U10302 ( .A(n9909), .B(n9911), .Y(n9904) );
  NAND2X1 U10303 ( .A(n9761), .B(n6883), .Y(n9902) );
  NAND2X1 U10304 ( .A(n9883), .B(G22), .Y(n9901) );
  NAND2X1 U10305 ( .A(G21704), .B(n9759), .Y(n9900) );
  NAND4X1 U10306 ( .A(n9914), .B(n9915), .C(n9916), .D(n9917), .Y(G1093) );
  NAND2X1 U10307 ( .A(n9772), .B(n6904), .Y(n9917) );
  NAND3X1 U10308 ( .A(n9918), .B(n9919), .C(n9920), .Y(n6904) );
  INVX1 U10309 ( .A(n9913), .Y(n9920) );
  NOR3X1 U10310 ( .A(n9921), .B(n9908), .C(n9922), .Y(n9913) );
  NAND2X1 U10311 ( .A(n9923), .B(n9908), .Y(n9919) );
  ADDHXL U10312 ( .A(n9924), .B(n9925), .S(n9923) );
  NAND2X1 U10313 ( .A(n9912), .B(n9926), .Y(n9918) );
  NAND2X1 U10314 ( .A(n9761), .B(n6902), .Y(n9916) );
  NAND2X1 U10315 ( .A(n9883), .B(G23), .Y(n9915) );
  NAND2X1 U10316 ( .A(G21703), .B(n9759), .Y(n9914) );
  NAND4X1 U10317 ( .A(n9927), .B(n9928), .C(n9929), .D(n9930), .Y(G1092) );
  NAND2X1 U10318 ( .A(n9772), .B(n6916), .Y(n9930) );
  ADDFXL U10319 ( .A(n9926), .B(n9931), .CI(n9932), .S(n6916) );
  NAND2X1 U10320 ( .A(n9761), .B(n6915), .Y(n9929) );
  NAND2X1 U10321 ( .A(n9883), .B(G24), .Y(n9928) );
  NAND2X1 U10322 ( .A(G21702), .B(n9759), .Y(n9927) );
  NAND4X1 U10323 ( .A(n9933), .B(n9934), .C(n9935), .D(n9936), .Y(G1091) );
  NAND2X1 U10324 ( .A(n9772), .B(n6927), .Y(n9936) );
  ADDHXL U10325 ( .A(n9937), .B(n9938), .S(n6927) );
  AND2X1 U10326 ( .A(n9939), .B(n9940), .Y(n9938) );
  NAND2X1 U10327 ( .A(n9761), .B(n6926), .Y(n9935) );
  NAND2X1 U10328 ( .A(n9883), .B(G25), .Y(n9934) );
  NAND2X1 U10329 ( .A(G21701), .B(n9759), .Y(n9933) );
  NAND4X1 U10330 ( .A(n9941), .B(n9942), .C(n9943), .D(n9944), .Y(G1090) );
  NAND2X1 U10331 ( .A(n9772), .B(n6938), .Y(n9944) );
  AND2X1 U10332 ( .A(n9945), .B(n9946), .Y(n6938) );
  NAND2X1 U10333 ( .A(n9947), .B(n9948), .Y(n9946) );
  INVX1 U10334 ( .A(n9949), .Y(n9947) );
  NAND3X1 U10335 ( .A(n9950), .B(n9951), .C(n9952), .Y(n9945) );
  NAND2X1 U10336 ( .A(n9948), .B(n9953), .Y(n9950) );
  NAND2X1 U10337 ( .A(n9761), .B(n6937), .Y(n9943) );
  NAND2X1 U10338 ( .A(n9883), .B(G26), .Y(n9942) );
  NAND2X1 U10339 ( .A(G21700), .B(n9759), .Y(n9941) );
  NAND4X1 U10340 ( .A(n9954), .B(n9955), .C(n9956), .D(n9957), .Y(G1089) );
  NAND2X1 U10341 ( .A(n9772), .B(n6949), .Y(n9957) );
  ADDHXL U10342 ( .A(n9958), .B(n9959), .S(n6949) );
  AND2X1 U10343 ( .A(n9951), .B(n9960), .Y(n9959) );
  NAND2X1 U10344 ( .A(n9761), .B(n6948), .Y(n9956) );
  NAND2X1 U10345 ( .A(n9883), .B(G27), .Y(n9955) );
  NAND2X1 U10346 ( .A(G21699), .B(n9759), .Y(n9954) );
  NAND4X1 U10347 ( .A(n9961), .B(n9962), .C(n9963), .D(n9964), .Y(G1088) );
  NAND2X1 U10348 ( .A(n9772), .B(n6960), .Y(n9964) );
  ADDHXL U10349 ( .A(n9965), .B(n9966), .S(n6960) );
  AND2X1 U10350 ( .A(n9967), .B(n9968), .Y(n9966) );
  NAND2X1 U10351 ( .A(n9761), .B(n6959), .Y(n9963) );
  NAND2X1 U10352 ( .A(n9883), .B(G28), .Y(n9962) );
  NAND2X1 U10353 ( .A(G21698), .B(n9759), .Y(n9961) );
  NAND4X1 U10354 ( .A(n9969), .B(n9970), .C(n9971), .D(n9972), .Y(G1087) );
  NAND2X1 U10355 ( .A(n9772), .B(n6970), .Y(n9972) );
  AND2X1 U10356 ( .A(n9973), .B(n9974), .Y(n6970) );
  NAND2X1 U10357 ( .A(n9975), .B(n9976), .Y(n9974) );
  NAND2X1 U10358 ( .A(n9977), .B(n9978), .Y(n9976) );
  INVX1 U10359 ( .A(n9979), .Y(n9975) );
  NAND3X1 U10360 ( .A(n9977), .B(n9978), .C(n9979), .Y(n9973) );
  NAND2X1 U10361 ( .A(n9761), .B(n6969), .Y(n9971) );
  NAND2X1 U10362 ( .A(n9883), .B(G29), .Y(n9970) );
  NAND2X1 U10363 ( .A(G21697), .B(n9759), .Y(n9969) );
  NAND4X1 U10364 ( .A(n9980), .B(n9981), .C(n9982), .D(n9983), .Y(G1086) );
  NAND2X1 U10365 ( .A(n9772), .B(n6980), .Y(n9983) );
  AND2X1 U10366 ( .A(n9984), .B(n9985), .Y(n6980) );
  NAND3X1 U10367 ( .A(n9986), .B(n9987), .C(n9988), .Y(n9985) );
  NAND2X1 U10368 ( .A(n9989), .B(n9990), .Y(n9986) );
  NAND2X1 U10369 ( .A(n9991), .B(n9989), .Y(n9984) );
  INVX1 U10370 ( .A(n9992), .Y(n9991) );
  NAND2X1 U10371 ( .A(n9761), .B(n6979), .Y(n9982) );
  NAND2X1 U10372 ( .A(n9883), .B(G30), .Y(n9981) );
  NAND2X1 U10373 ( .A(G21696), .B(n9759), .Y(n9980) );
  NAND4X1 U10374 ( .A(n9993), .B(n9994), .C(n9995), .D(n9996), .Y(G1085) );
  NAND2X1 U10375 ( .A(n9772), .B(n6991), .Y(n9996) );
  ADDHXL U10376 ( .A(n9997), .B(n9998), .S(n6991) );
  AND2X1 U10377 ( .A(n9987), .B(n9999), .Y(n9998) );
  NAND2X1 U10378 ( .A(n9761), .B(n6990), .Y(n9995) );
  NAND2X1 U10379 ( .A(n9883), .B(G31), .Y(n9994) );
  NAND2X1 U10380 ( .A(G21695), .B(n9759), .Y(n9993) );
  NAND4X1 U10381 ( .A(n10000), .B(n10001), .C(n10002), .D(n10003), .Y(G1084)
         );
  NAND2X1 U10382 ( .A(n9761), .B(n7001), .Y(n10003) );
  NOR2X1 U10383 ( .A(n9759), .B(n9193), .Y(n9761) );
  NAND2X1 U10384 ( .A(n9772), .B(n7002), .Y(n10002) );
  ADDHXL U10385 ( .A(n9926), .B(n10004), .S(n7002) );
  NOR2X1 U10386 ( .A(n10005), .B(n10006), .Y(n10004) );
  INVX1 U10387 ( .A(n10007), .Y(n10005) );
  NAND2X1 U10388 ( .A(n9883), .B(G32), .Y(n10001) );
  NOR2X1 U10389 ( .A(n9759), .B(n9224), .Y(n9883) );
  NAND2X1 U10390 ( .A(G21694), .B(n9759), .Y(n10000) );
  NAND3X1 U10391 ( .A(n7441), .B(n7445), .C(n9260), .Y(n10011) );
  NAND2X1 U10392 ( .A(n10013), .B(n7447), .Y(n10010) );
  NOR2X1 U10393 ( .A(n9092), .B(G35), .Y(n7447) );
  NAND2X1 U10394 ( .A(n10014), .B(n7457), .Y(n10009) );
  AND2X1 U10395 ( .A(G21693), .B(n10015), .Y(G1083) );
  NAND3X1 U10396 ( .A(n10016), .B(n10017), .C(n10018), .Y(G1082) );
  NAND2X1 U10397 ( .A(G21692), .B(n10015), .Y(n10018) );
  NAND2X1 U10398 ( .A(n10019), .B(G21724), .Y(n10017) );
  NAND2X1 U10399 ( .A(G21647), .B(n10020), .Y(n10016) );
  NAND3X1 U10400 ( .A(n10021), .B(n10022), .C(n10023), .Y(G1081) );
  NAND2X1 U10401 ( .A(G21691), .B(n10015), .Y(n10023) );
  NAND2X1 U10402 ( .A(n10019), .B(G21723), .Y(n10022) );
  NAND2X1 U10403 ( .A(G21648), .B(n10020), .Y(n10021) );
  NAND3X1 U10404 ( .A(n10024), .B(n10025), .C(n10026), .Y(G1080) );
  NAND2X1 U10405 ( .A(G21690), .B(n10015), .Y(n10026) );
  NAND2X1 U10406 ( .A(n10019), .B(G21722), .Y(n10025) );
  NAND2X1 U10407 ( .A(G21649), .B(n10020), .Y(n10024) );
  NAND3X1 U10408 ( .A(n10027), .B(n10028), .C(n10029), .Y(G1079) );
  NAND2X1 U10409 ( .A(G21689), .B(n10015), .Y(n10029) );
  NAND2X1 U10410 ( .A(n10019), .B(G21721), .Y(n10028) );
  NAND2X1 U10411 ( .A(G21650), .B(n10020), .Y(n10027) );
  NAND3X1 U10412 ( .A(n10030), .B(n10031), .C(n10032), .Y(G1078) );
  NAND2X1 U10413 ( .A(G21688), .B(n10015), .Y(n10032) );
  NAND2X1 U10414 ( .A(n10019), .B(G21720), .Y(n10031) );
  NAND2X1 U10415 ( .A(G21651), .B(n10020), .Y(n10030) );
  NAND3X1 U10416 ( .A(n10033), .B(n10034), .C(n10035), .Y(G1077) );
  NAND2X1 U10417 ( .A(G21687), .B(n10015), .Y(n10035) );
  NAND2X1 U10418 ( .A(n10019), .B(G21719), .Y(n10034) );
  NAND2X1 U10419 ( .A(G21652), .B(n10020), .Y(n10033) );
  NAND3X1 U10420 ( .A(n10036), .B(n10037), .C(n10038), .Y(G1076) );
  NAND2X1 U10421 ( .A(G21686), .B(n10015), .Y(n10038) );
  NAND2X1 U10422 ( .A(n10019), .B(G21718), .Y(n10037) );
  NAND2X1 U10423 ( .A(G21653), .B(n10020), .Y(n10036) );
  NAND3X1 U10424 ( .A(n10039), .B(n10040), .C(n10041), .Y(G1075) );
  NAND2X1 U10425 ( .A(G21685), .B(n10015), .Y(n10041) );
  NAND2X1 U10426 ( .A(n10019), .B(G21717), .Y(n10040) );
  NAND2X1 U10427 ( .A(G21654), .B(n10020), .Y(n10039) );
  NAND3X1 U10428 ( .A(n10042), .B(n10043), .C(n10044), .Y(G1074) );
  NAND2X1 U10429 ( .A(G21684), .B(n10015), .Y(n10044) );
  NAND2X1 U10430 ( .A(n10019), .B(G21716), .Y(n10043) );
  NAND2X1 U10431 ( .A(G21655), .B(n10020), .Y(n10042) );
  NAND3X1 U10432 ( .A(n10045), .B(n10046), .C(n10047), .Y(G1073) );
  NAND2X1 U10433 ( .A(G21683), .B(n10015), .Y(n10047) );
  NAND2X1 U10434 ( .A(n10019), .B(G21715), .Y(n10046) );
  NAND2X1 U10435 ( .A(G21656), .B(n10020), .Y(n10045) );
  NAND3X1 U10436 ( .A(n10048), .B(n10049), .C(n10050), .Y(G1072) );
  NAND2X1 U10437 ( .A(G21682), .B(n10015), .Y(n10050) );
  NAND2X1 U10438 ( .A(n10019), .B(G21714), .Y(n10049) );
  NAND2X1 U10439 ( .A(G21657), .B(n10020), .Y(n10048) );
  NAND3X1 U10440 ( .A(n10051), .B(n10052), .C(n10053), .Y(G1071) );
  NAND2X1 U10441 ( .A(G21681), .B(n10015), .Y(n10053) );
  NAND2X1 U10442 ( .A(n10019), .B(G21713), .Y(n10052) );
  NAND2X1 U10443 ( .A(G21658), .B(n10020), .Y(n10051) );
  NAND3X1 U10444 ( .A(n10054), .B(n10055), .C(n10056), .Y(G1070) );
  NAND2X1 U10445 ( .A(G21680), .B(n10015), .Y(n10056) );
  NAND2X1 U10446 ( .A(n10019), .B(G21712), .Y(n10055) );
  NAND2X1 U10447 ( .A(G21659), .B(n10020), .Y(n10054) );
  NAND3X1 U10448 ( .A(n10057), .B(n10058), .C(n10059), .Y(G1069) );
  NAND2X1 U10449 ( .A(G21679), .B(n10015), .Y(n10059) );
  NAND2X1 U10450 ( .A(n10019), .B(G21711), .Y(n10058) );
  NAND2X1 U10451 ( .A(G21660), .B(n10020), .Y(n10057) );
  NAND3X1 U10452 ( .A(n10060), .B(n10061), .C(n10062), .Y(G1068) );
  NAND2X1 U10453 ( .A(G21678), .B(n10015), .Y(n10062) );
  NAND2X1 U10454 ( .A(n10019), .B(G21710), .Y(n10061) );
  AND2X1 U10455 ( .A(n10063), .B(n8711), .Y(n10019) );
  NAND2X1 U10456 ( .A(G21661), .B(n10020), .Y(n10060) );
  NAND3X1 U10457 ( .A(n10064), .B(n10065), .C(n10066), .Y(G1067) );
  NAND2X1 U10458 ( .A(G21677), .B(n10015), .Y(n10066) );
  NAND2X1 U10459 ( .A(n10063), .B(G21709), .Y(n10065) );
  NAND2X1 U10460 ( .A(G21631), .B(n10020), .Y(n10064) );
  NAND3X1 U10461 ( .A(n10067), .B(n10068), .C(n10069), .Y(G1066) );
  NAND2X1 U10462 ( .A(G21676), .B(n10015), .Y(n10069) );
  NAND2X1 U10463 ( .A(n10063), .B(G21708), .Y(n10068) );
  NAND2X1 U10464 ( .A(G21632), .B(n10020), .Y(n10067) );
  NAND3X1 U10465 ( .A(n10070), .B(n10071), .C(n10072), .Y(G1065) );
  NAND2X1 U10466 ( .A(G21675), .B(n10015), .Y(n10072) );
  NAND2X1 U10467 ( .A(n10063), .B(G21707), .Y(n10071) );
  NAND2X1 U10468 ( .A(G21633), .B(n10020), .Y(n10070) );
  NAND3X1 U10469 ( .A(n10073), .B(n10074), .C(n10075), .Y(G1064) );
  NAND2X1 U10470 ( .A(G21674), .B(n10015), .Y(n10075) );
  NAND2X1 U10471 ( .A(n10063), .B(G21706), .Y(n10074) );
  NAND2X1 U10472 ( .A(G21634), .B(n10020), .Y(n10073) );
  NAND3X1 U10473 ( .A(n10076), .B(n10077), .C(n10078), .Y(G1063) );
  NAND2X1 U10474 ( .A(G21673), .B(n10015), .Y(n10078) );
  NAND2X1 U10475 ( .A(n10063), .B(G21705), .Y(n10077) );
  NAND2X1 U10476 ( .A(G21635), .B(n10020), .Y(n10076) );
  NAND3X1 U10477 ( .A(n10079), .B(n10080), .C(n10081), .Y(G1062) );
  NAND2X1 U10478 ( .A(G21672), .B(n10015), .Y(n10081) );
  NAND2X1 U10479 ( .A(n10063), .B(G21704), .Y(n10080) );
  NAND2X1 U10480 ( .A(G21636), .B(n10020), .Y(n10079) );
  NAND3X1 U10481 ( .A(n10082), .B(n10083), .C(n10084), .Y(G1061) );
  NAND2X1 U10482 ( .A(G21671), .B(n10015), .Y(n10084) );
  NAND2X1 U10483 ( .A(n10063), .B(G21703), .Y(n10083) );
  NAND2X1 U10484 ( .A(G21637), .B(n10020), .Y(n10082) );
  NAND3X1 U10485 ( .A(n10085), .B(n10086), .C(n10087), .Y(G1060) );
  NAND2X1 U10486 ( .A(G21670), .B(n10015), .Y(n10087) );
  NAND2X1 U10487 ( .A(n10063), .B(G21702), .Y(n10086) );
  NAND2X1 U10488 ( .A(G21638), .B(n10020), .Y(n10085) );
  NAND3X1 U10489 ( .A(n10088), .B(n10089), .C(n10090), .Y(G1059) );
  NAND2X1 U10490 ( .A(G21669), .B(n10015), .Y(n10090) );
  NAND2X1 U10491 ( .A(n10063), .B(G21701), .Y(n10089) );
  NAND2X1 U10492 ( .A(G21639), .B(n10020), .Y(n10088) );
  NAND3X1 U10493 ( .A(n10091), .B(n10092), .C(n10093), .Y(G1058) );
  NAND2X1 U10494 ( .A(G21668), .B(n10015), .Y(n10093) );
  NAND2X1 U10495 ( .A(n10063), .B(G21700), .Y(n10092) );
  NAND2X1 U10496 ( .A(G21640), .B(n10020), .Y(n10091) );
  NAND3X1 U10497 ( .A(n10094), .B(n10095), .C(n10096), .Y(G1057) );
  NAND2X1 U10498 ( .A(G21667), .B(n10015), .Y(n10096) );
  NAND2X1 U10499 ( .A(n10063), .B(G21699), .Y(n10095) );
  NAND2X1 U10500 ( .A(G21641), .B(n10020), .Y(n10094) );
  NAND3X1 U10501 ( .A(n10097), .B(n10098), .C(n10099), .Y(G1056) );
  NAND2X1 U10502 ( .A(G21666), .B(n10015), .Y(n10099) );
  NAND2X1 U10503 ( .A(n10063), .B(G21698), .Y(n10098) );
  NAND2X1 U10504 ( .A(G21642), .B(n10020), .Y(n10097) );
  NAND3X1 U10505 ( .A(n10100), .B(n10101), .C(n10102), .Y(G1055) );
  NAND2X1 U10506 ( .A(G21665), .B(n10015), .Y(n10102) );
  NAND2X1 U10507 ( .A(n10063), .B(G21697), .Y(n10101) );
  NAND2X1 U10508 ( .A(G21643), .B(n10020), .Y(n10100) );
  NAND3X1 U10509 ( .A(n10103), .B(n10104), .C(n10105), .Y(G1054) );
  NAND2X1 U10510 ( .A(G21664), .B(n10015), .Y(n10105) );
  NAND2X1 U10511 ( .A(n10063), .B(G21696), .Y(n10104) );
  NAND2X1 U10512 ( .A(G21644), .B(n10020), .Y(n10103) );
  NAND3X1 U10513 ( .A(n10106), .B(n10107), .C(n10108), .Y(G1053) );
  NAND2X1 U10514 ( .A(G21663), .B(n10015), .Y(n10108) );
  NAND2X1 U10515 ( .A(n10063), .B(G21695), .Y(n10107) );
  NAND2X1 U10516 ( .A(G21645), .B(n10020), .Y(n10106) );
  NAND3X1 U10517 ( .A(n10109), .B(n10110), .C(n10111), .Y(G1052) );
  NAND2X1 U10518 ( .A(G21662), .B(n10015), .Y(n10111) );
  NAND2X1 U10519 ( .A(n10063), .B(G21694), .Y(n10110) );
  NOR2X1 U10520 ( .A(n8817), .B(n10015), .Y(n10063) );
  NAND2X1 U10521 ( .A(G21646), .B(n10020), .Y(n10109) );
  NAND2X1 U10522 ( .A(n7454), .B(n10114), .Y(n10113) );
  NAND2X1 U10523 ( .A(n9644), .B(n10115), .Y(n10114) );
  NAND3X1 U10524 ( .A(n9175), .B(n7457), .C(n7433), .Y(n10115) );
  NOR2X1 U10525 ( .A(G21392), .B(n10116), .Y(n7454) );
  NAND2X1 U10526 ( .A(n9071), .B(G21427), .Y(n10112) );
  NAND3X1 U10527 ( .A(n10117), .B(n10118), .C(n10119), .Y(G1051) );
  NAND2X1 U10528 ( .A(n10120), .B(G21661), .Y(n10119) );
  NAND2X1 U10529 ( .A(n10121), .B(G21710), .Y(n10117) );
  NAND3X1 U10530 ( .A(n10122), .B(n10123), .C(n10124), .Y(G1050) );
  NAND2X1 U10531 ( .A(n10120), .B(G21660), .Y(n10124) );
  NAND2X1 U10532 ( .A(n10121), .B(G21711), .Y(n10122) );
  NAND3X1 U10533 ( .A(n10125), .B(n10126), .C(n10127), .Y(G1049) );
  NAND2X1 U10534 ( .A(n10120), .B(G21659), .Y(n10127) );
  NAND2X1 U10535 ( .A(n10121), .B(G21712), .Y(n10125) );
  NAND3X1 U10536 ( .A(n10128), .B(n10129), .C(n10130), .Y(G1048) );
  NAND2X1 U10537 ( .A(n10120), .B(G21658), .Y(n10130) );
  NAND2X1 U10538 ( .A(n10121), .B(G21713), .Y(n10128) );
  NAND3X1 U10539 ( .A(n10131), .B(n10132), .C(n10133), .Y(G1047) );
  NAND2X1 U10540 ( .A(n10120), .B(G21657), .Y(n10133) );
  NAND2X1 U10541 ( .A(n10121), .B(G21714), .Y(n10131) );
  NAND3X1 U10542 ( .A(n10134), .B(n10135), .C(n10136), .Y(G1046) );
  NAND2X1 U10543 ( .A(n10120), .B(G21656), .Y(n10136) );
  NAND2X1 U10544 ( .A(n10121), .B(G21715), .Y(n10134) );
  NAND3X1 U10545 ( .A(n10137), .B(n10138), .C(n10139), .Y(G1045) );
  NAND2X1 U10546 ( .A(n10120), .B(G21655), .Y(n10139) );
  NAND2X1 U10547 ( .A(n10121), .B(G21716), .Y(n10137) );
  NAND3X1 U10548 ( .A(n10140), .B(n10141), .C(n10142), .Y(G1044) );
  NAND2X1 U10549 ( .A(n10120), .B(G21654), .Y(n10142) );
  NAND2X1 U10550 ( .A(n10121), .B(G21717), .Y(n10140) );
  NAND3X1 U10551 ( .A(n10143), .B(n10144), .C(n10145), .Y(G1043) );
  NAND2X1 U10552 ( .A(n10120), .B(G21653), .Y(n10145) );
  NAND2X1 U10553 ( .A(n10121), .B(G21718), .Y(n10143) );
  NAND3X1 U10554 ( .A(n10146), .B(n10147), .C(n10148), .Y(G1042) );
  NAND2X1 U10555 ( .A(n10120), .B(G21652), .Y(n10148) );
  NAND2X1 U10556 ( .A(n10121), .B(G21719), .Y(n10146) );
  NAND3X1 U10557 ( .A(n10149), .B(n10150), .C(n10151), .Y(G1041) );
  NAND2X1 U10558 ( .A(n10120), .B(G21651), .Y(n10151) );
  NAND2X1 U10559 ( .A(n10121), .B(G21720), .Y(n10149) );
  NAND3X1 U10560 ( .A(n10152), .B(n10153), .C(n10154), .Y(G1040) );
  NAND2X1 U10561 ( .A(n10120), .B(G21650), .Y(n10154) );
  NAND2X1 U10562 ( .A(n10121), .B(G21721), .Y(n10152) );
  NAND3X1 U10563 ( .A(n10155), .B(n10156), .C(n10157), .Y(G1039) );
  NAND2X1 U10564 ( .A(n10120), .B(G21649), .Y(n10157) );
  NAND2X1 U10565 ( .A(n10121), .B(G21722), .Y(n10155) );
  NAND3X1 U10566 ( .A(n10158), .B(n10159), .C(n10160), .Y(G1038) );
  NAND2X1 U10567 ( .A(n10120), .B(G21648), .Y(n10160) );
  NAND2X1 U10568 ( .A(n10121), .B(G21723), .Y(n10158) );
  NAND3X1 U10569 ( .A(n10161), .B(n10162), .C(n10163), .Y(G1037) );
  NAND2X1 U10570 ( .A(n10120), .B(G21647), .Y(n10163) );
  NAND2X1 U10571 ( .A(n10121), .B(G21724), .Y(n10161) );
  NAND3X1 U10572 ( .A(n10164), .B(n10118), .C(n10165), .Y(G1036) );
  NAND2X1 U10573 ( .A(n10120), .B(G21646), .Y(n10165) );
  NAND2X1 U10574 ( .A(n10166), .B(G32), .Y(n10118) );
  NAND2X1 U10575 ( .A(n10121), .B(G21694), .Y(n10164) );
  NAND3X1 U10576 ( .A(n10167), .B(n10123), .C(n10168), .Y(G1035) );
  NAND2X1 U10577 ( .A(n10120), .B(G21645), .Y(n10168) );
  NAND2X1 U10578 ( .A(n10166), .B(G31), .Y(n10123) );
  NAND2X1 U10579 ( .A(n10121), .B(G21695), .Y(n10167) );
  NAND3X1 U10580 ( .A(n10169), .B(n10126), .C(n10170), .Y(G1034) );
  NAND2X1 U10581 ( .A(n10120), .B(G21644), .Y(n10170) );
  NAND2X1 U10582 ( .A(n10166), .B(G30), .Y(n10126) );
  NAND2X1 U10583 ( .A(n10121), .B(G21696), .Y(n10169) );
  NAND3X1 U10584 ( .A(n10171), .B(n10129), .C(n10172), .Y(G1033) );
  NAND2X1 U10585 ( .A(n10120), .B(G21643), .Y(n10172) );
  NAND2X1 U10586 ( .A(n10166), .B(G29), .Y(n10129) );
  NAND2X1 U10587 ( .A(n10121), .B(G21697), .Y(n10171) );
  NAND3X1 U10588 ( .A(n10173), .B(n10132), .C(n10174), .Y(G1032) );
  NAND2X1 U10589 ( .A(n10120), .B(G21642), .Y(n10174) );
  NAND2X1 U10590 ( .A(n10166), .B(G28), .Y(n10132) );
  NAND2X1 U10591 ( .A(n10121), .B(G21698), .Y(n10173) );
  NAND3X1 U10592 ( .A(n10175), .B(n10135), .C(n10176), .Y(G1031) );
  NAND2X1 U10593 ( .A(n10120), .B(G21641), .Y(n10176) );
  NAND2X1 U10594 ( .A(n10166), .B(G27), .Y(n10135) );
  NAND2X1 U10595 ( .A(n10121), .B(G21699), .Y(n10175) );
  NAND3X1 U10596 ( .A(n10177), .B(n10138), .C(n10178), .Y(G1030) );
  NAND2X1 U10597 ( .A(n10120), .B(G21640), .Y(n10178) );
  NAND2X1 U10598 ( .A(n10166), .B(G26), .Y(n10138) );
  NAND2X1 U10599 ( .A(n10121), .B(G21700), .Y(n10177) );
  NAND3X1 U10600 ( .A(n10179), .B(n10141), .C(n10180), .Y(G1029) );
  NAND2X1 U10601 ( .A(n10120), .B(G21639), .Y(n10180) );
  NAND2X1 U10602 ( .A(n10166), .B(G25), .Y(n10141) );
  NAND2X1 U10603 ( .A(n10121), .B(G21701), .Y(n10179) );
  NAND3X1 U10604 ( .A(n10181), .B(n10144), .C(n10182), .Y(G1028) );
  NAND2X1 U10605 ( .A(n10120), .B(G21638), .Y(n10182) );
  NAND2X1 U10606 ( .A(n10166), .B(G24), .Y(n10144) );
  NAND2X1 U10607 ( .A(n10121), .B(G21702), .Y(n10181) );
  NAND3X1 U10608 ( .A(n10183), .B(n10147), .C(n10184), .Y(G1027) );
  NAND2X1 U10609 ( .A(n10120), .B(G21637), .Y(n10184) );
  NAND2X1 U10610 ( .A(n10166), .B(G23), .Y(n10147) );
  NAND2X1 U10611 ( .A(n10121), .B(G21703), .Y(n10183) );
  NAND3X1 U10612 ( .A(n10185), .B(n10150), .C(n10186), .Y(G1026) );
  NAND2X1 U10613 ( .A(n10120), .B(G21636), .Y(n10186) );
  NAND2X1 U10614 ( .A(n10166), .B(G22), .Y(n10150) );
  NAND2X1 U10615 ( .A(n10121), .B(G21704), .Y(n10185) );
  NAND3X1 U10616 ( .A(n10187), .B(n10153), .C(n10188), .Y(G1025) );
  NAND2X1 U10617 ( .A(n10120), .B(G21635), .Y(n10188) );
  NAND2X1 U10618 ( .A(n10166), .B(G21), .Y(n10153) );
  NAND2X1 U10619 ( .A(n10121), .B(G21705), .Y(n10187) );
  NAND3X1 U10620 ( .A(n10189), .B(n10156), .C(n10190), .Y(G1024) );
  NAND2X1 U10621 ( .A(n10120), .B(G21634), .Y(n10190) );
  NAND2X1 U10622 ( .A(n10166), .B(G20), .Y(n10156) );
  NAND2X1 U10623 ( .A(n10121), .B(G21706), .Y(n10189) );
  NAND3X1 U10624 ( .A(n10191), .B(n10159), .C(n10192), .Y(G1023) );
  NAND2X1 U10625 ( .A(n10120), .B(G21633), .Y(n10192) );
  NAND2X1 U10626 ( .A(n10166), .B(G19), .Y(n10159) );
  NAND2X1 U10627 ( .A(n10121), .B(G21707), .Y(n10191) );
  NAND3X1 U10628 ( .A(n10193), .B(n10162), .C(n10194), .Y(G1022) );
  NAND2X1 U10629 ( .A(n10120), .B(G21632), .Y(n10194) );
  NAND2X1 U10630 ( .A(n10166), .B(G18), .Y(n10162) );
  NAND2X1 U10631 ( .A(n10121), .B(G21708), .Y(n10193) );
  NAND3X1 U10632 ( .A(n10195), .B(n10196), .C(n10197), .Y(G1021) );
  NAND2X1 U10633 ( .A(n10120), .B(G21631), .Y(n10197) );
  NAND2X1 U10634 ( .A(n10166), .B(G17), .Y(n10196) );
  NOR2X1 U10635 ( .A(n7451), .B(n10120), .Y(n10166) );
  NAND2X1 U10636 ( .A(n10121), .B(G21709), .Y(n10195) );
  NAND3X1 U10637 ( .A(n8856), .B(n7457), .C(n7433), .Y(n9644) );
  NOR2X1 U10638 ( .A(n8828), .B(n8817), .Y(n7433) );
  INVX1 U10639 ( .A(n8818), .Y(n8828) );
  NAND4X1 U10640 ( .A(n8818), .B(n9260), .C(n7441), .D(n7445), .Y(n10198) );
  INVX1 U10641 ( .A(G35), .Y(n7445) );
  NOR2X1 U10642 ( .A(n7430), .B(G21427), .Y(n8818) );
  NAND4X1 U10643 ( .A(n10199), .B(n10200), .C(n10201), .D(n10202), .Y(G1020)
         );
  NOR2X1 U10644 ( .A(n10203), .B(n10204), .Y(n10202) );
  NOR2X1 U10645 ( .A(n6891), .B(n9318), .Y(n10204) );
  NOR2X1 U10646 ( .A(n6901), .B(n7018), .Y(n10203) );
  NAND2X1 U10647 ( .A(n6905), .B(n7023), .Y(n10201) );
  NAND2X1 U10648 ( .A(n6903), .B(n7021), .Y(n10200) );
  ADDFXL U10649 ( .A(n9908), .B(n10205), .CI(n10206), .S(n7021) );
  NAND2X1 U10650 ( .A(n10207), .B(n10208), .Y(n10206) );
  NAND2X1 U10651 ( .A(n9926), .B(n10209), .Y(n10208) );
  OR2X1 U10652 ( .A(n10210), .B(n10211), .Y(n10209) );
  NAND2X1 U10653 ( .A(n10211), .B(n10210), .Y(n10207) );
  NOR4X1 U10654 ( .A(n10212), .B(n10213), .C(n10214), .D(n10215), .Y(n10205)
         );
  NOR2X1 U10655 ( .A(n10216), .B(n7014), .Y(n10215) );
  NOR2X1 U10656 ( .A(n10217), .B(n9323), .Y(n10214) );
  INVX1 U10657 ( .A(n7023), .Y(n9323) );
  ADDHXL U10658 ( .A(n10218), .B(n10219), .S(n7023) );
  NAND2X1 U10659 ( .A(n9085), .B(n10220), .Y(n10218) );
  NAND3X1 U10660 ( .A(n10221), .B(n10222), .C(n10223), .Y(n10220) );
  NAND2X1 U10661 ( .A(G21789), .B(n9260), .Y(n10223) );
  NAND2X1 U10662 ( .A(G21598), .B(n10224), .Y(n10222) );
  NAND2X1 U10663 ( .A(G21630), .B(n10225), .Y(n10221) );
  NOR2X1 U10664 ( .A(n9908), .B(n9640), .Y(n10213) );
  NOR2X1 U10665 ( .A(n10226), .B(n7018), .Y(n10212) );
  INVX1 U10666 ( .A(G21789), .Y(n7018) );
  NAND2X1 U10667 ( .A(n7025), .B(n6882), .Y(n10199) );
  INVX1 U10668 ( .A(n9640), .Y(n7025) );
  ADDFXL U10669 ( .A(n10227), .B(n10228), .CI(n10229), .S(n9640) );
  NOR4X1 U10670 ( .A(n10230), .B(n10231), .C(n10232), .D(n10233), .Y(n10228)
         );
  NOR2X1 U10671 ( .A(n10234), .B(n7014), .Y(n10233) );
  NOR2X1 U10672 ( .A(n10235), .B(n9320), .Y(n10232) );
  AND2X1 U10673 ( .A(n10236), .B(G21725), .Y(n10231) );
  NOR2X1 U10674 ( .A(n9085), .B(n9318), .Y(n10230) );
  INVX1 U10675 ( .A(G21630), .Y(n9318) );
  NAND4X1 U10676 ( .A(n10237), .B(n10238), .C(n10239), .D(n10240), .Y(G1019)
         );
  NOR2X1 U10677 ( .A(n10241), .B(n10242), .Y(n10240) );
  NOR2X1 U10678 ( .A(n6891), .B(n9334), .Y(n10242) );
  NOR2X1 U10679 ( .A(n6901), .B(n7033), .Y(n10241) );
  NAND2X1 U10680 ( .A(n7039), .B(n6882), .Y(n10239) );
  NAND2X1 U10681 ( .A(n6903), .B(n7037), .Y(n10238) );
  ADDFXL U10682 ( .A(n9926), .B(n10210), .CI(n10211), .S(n7037) );
  NAND2X1 U10683 ( .A(n10243), .B(n10244), .Y(n10211) );
  NAND2X1 U10684 ( .A(n9926), .B(n10245), .Y(n10244) );
  OR2X1 U10685 ( .A(n10246), .B(n10247), .Y(n10245) );
  NAND2X1 U10686 ( .A(n10247), .B(n10246), .Y(n10243) );
  NAND4X1 U10687 ( .A(n10248), .B(n10249), .C(n10250), .D(n10251), .Y(n10210)
         );
  NOR2X1 U10688 ( .A(n10252), .B(n10253), .Y(n10251) );
  NOR2X1 U10689 ( .A(n10216), .B(n7035), .Y(n10253) );
  NOR2X1 U10690 ( .A(n10226), .B(n7033), .Y(n10252) );
  NAND2X1 U10691 ( .A(n7039), .B(n9926), .Y(n10250) );
  NAND2X1 U10692 ( .A(n7038), .B(n10257), .Y(n10255) );
  NAND2X1 U10693 ( .A(n10258), .B(n9336), .Y(n10254) );
  NAND2X1 U10694 ( .A(n10259), .B(n10257), .Y(n10258) );
  NOR2X1 U10695 ( .A(n9356), .B(n7048), .Y(n10257) );
  NAND2X1 U10696 ( .A(n7038), .B(n10260), .Y(n10248) );
  NAND2X1 U10697 ( .A(n7038), .B(n6905), .Y(n10237) );
  INVX1 U10698 ( .A(n9336), .Y(n7038) );
  NAND2X1 U10699 ( .A(n10219), .B(n10261), .Y(n9336) );
  NAND2X1 U10700 ( .A(n10262), .B(n10263), .Y(n10261) );
  OR2X1 U10701 ( .A(n10263), .B(n10262), .Y(n10219) );
  ADDHXL U10702 ( .A(n10264), .B(n9085), .S(n10262) );
  NAND4X1 U10703 ( .A(n10265), .B(n10266), .C(n10267), .D(n10268), .Y(n10264)
         );
  NOR2X1 U10704 ( .A(n10269), .B(n10270), .Y(n10268) );
  NOR2X1 U10705 ( .A(n10271), .B(n9334), .Y(n10270) );
  INVX1 U10706 ( .A(G21629), .Y(n9334) );
  NOR2X1 U10707 ( .A(n10227), .B(n7033), .Y(n10269) );
  INVX1 U10708 ( .A(G21788), .Y(n7033) );
  NAND2X1 U10709 ( .A(G21597), .B(n10224), .Y(n10267) );
  NAND2X1 U10710 ( .A(n7039), .B(n10272), .Y(n10266) );
  INVX1 U10711 ( .A(n9770), .Y(n7039) );
  NAND2X1 U10712 ( .A(n10229), .B(n10273), .Y(n9770) );
  NAND2X1 U10713 ( .A(n10274), .B(n10275), .Y(n10273) );
  OR2X1 U10714 ( .A(n10275), .B(n10274), .Y(n10229) );
  ADDHXL U10715 ( .A(n9260), .B(n10276), .S(n10274) );
  NOR3X1 U10716 ( .A(n10277), .B(n10278), .C(n10279), .Y(n10276) );
  NOR2X1 U10717 ( .A(n9266), .B(n7034), .Y(n10279) );
  NAND2X1 U10718 ( .A(n7012), .B(n10280), .Y(n7034) );
  NAND2X1 U10719 ( .A(n10281), .B(n10282), .Y(n10280) );
  INVX1 U10720 ( .A(n7017), .Y(n7012) );
  NOR2X1 U10721 ( .A(n10282), .B(n10281), .Y(n7017) );
  NAND2X1 U10722 ( .A(n10283), .B(n10284), .Y(n10281) );
  NAND2X1 U10723 ( .A(n9076), .B(n7035), .Y(n10284) );
  NAND4X1 U10724 ( .A(n10285), .B(n10286), .C(n10287), .D(n8711), .Y(n10283)
         );
  NOR2X1 U10725 ( .A(n10288), .B(n10289), .Y(n10287) );
  NAND4X1 U10726 ( .A(n10290), .B(n10291), .C(n10292), .D(n10293), .Y(n10289)
         );
  NAND2X1 U10727 ( .A(n10294), .B(G21493), .Y(n10293) );
  NAND2X1 U10728 ( .A(n10295), .B(G21501), .Y(n10292) );
  NAND2X1 U10729 ( .A(n10296), .B(G21509), .Y(n10291) );
  NAND2X1 U10730 ( .A(n10297), .B(G21517), .Y(n10290) );
  NAND4X1 U10731 ( .A(n10298), .B(n10299), .C(n10300), .D(n10301), .Y(n10288)
         );
  NAND2X1 U10732 ( .A(n10302), .B(G21525), .Y(n10301) );
  NAND2X1 U10733 ( .A(n10303), .B(G21533), .Y(n10300) );
  NAND2X1 U10734 ( .A(n10304), .B(G21541), .Y(n10299) );
  NAND2X1 U10735 ( .A(n10305), .B(G21549), .Y(n10298) );
  NOR4X1 U10736 ( .A(n10306), .B(n10307), .C(n10308), .D(n10309), .Y(n10286)
         );
  NOR2X1 U10737 ( .A(n10310), .B(n10311), .Y(n10309) );
  NOR2X1 U10738 ( .A(n10312), .B(n10313), .Y(n10308) );
  NOR2X1 U10739 ( .A(n10314), .B(n10315), .Y(n10307) );
  NOR2X1 U10740 ( .A(n10316), .B(n10317), .Y(n10306) );
  NOR4X1 U10741 ( .A(n10318), .B(n10319), .C(n10320), .D(n10321), .Y(n10285)
         );
  NOR2X1 U10742 ( .A(n10322), .B(n10323), .Y(n10321) );
  NOR2X1 U10743 ( .A(n10324), .B(n10325), .Y(n10320) );
  NOR2X1 U10744 ( .A(n10326), .B(n10327), .Y(n10319) );
  NOR2X1 U10745 ( .A(n10328), .B(n10329), .Y(n10318) );
  NOR2X1 U10746 ( .A(n10234), .B(n7035), .Y(n10278) );
  INVX1 U10747 ( .A(G21597), .Y(n7035) );
  NAND3X1 U10748 ( .A(n10330), .B(n10331), .C(n10332), .Y(n10277) );
  NAND2X1 U10749 ( .A(G21756), .B(n10333), .Y(n10332) );
  NAND2X1 U10750 ( .A(G21629), .B(n7564), .Y(n10331) );
  NAND2X1 U10751 ( .A(G21724), .B(n10236), .Y(n10330) );
  NAND2X1 U10752 ( .A(n10334), .B(n10335), .Y(n10275) );
  NAND2X1 U10753 ( .A(n10014), .B(n10336), .Y(n10265) );
  NAND2X1 U10754 ( .A(n10337), .B(n10338), .Y(n10263) );
  INVX1 U10755 ( .A(n10339), .Y(n10337) );
  NAND4X1 U10756 ( .A(n10340), .B(n10341), .C(n10342), .D(n10343), .Y(G1018)
         );
  NOR2X1 U10757 ( .A(n10344), .B(n10345), .Y(n10343) );
  NOR2X1 U10758 ( .A(n6891), .B(n9344), .Y(n10345) );
  NOR2X1 U10759 ( .A(n6901), .B(n10346), .Y(n10344) );
  NAND2X1 U10760 ( .A(n9346), .B(n6882), .Y(n10342) );
  NAND2X1 U10761 ( .A(n6903), .B(n7053), .Y(n10341) );
  ADDFXL U10762 ( .A(n9926), .B(n10247), .CI(n10246), .S(n7053) );
  NAND2X1 U10763 ( .A(n10347), .B(n10348), .Y(n10246) );
  NAND2X1 U10764 ( .A(n9926), .B(n10349), .Y(n10348) );
  OR2X1 U10765 ( .A(n10350), .B(n10351), .Y(n10349) );
  NAND2X1 U10766 ( .A(n10351), .B(n10350), .Y(n10347) );
  NAND4X1 U10767 ( .A(n10352), .B(n10353), .C(n10354), .D(n10355), .Y(n10247)
         );
  NOR2X1 U10768 ( .A(n10356), .B(n10357), .Y(n10355) );
  NOR2X1 U10769 ( .A(n10216), .B(n10358), .Y(n10357) );
  NOR2X1 U10770 ( .A(n10226), .B(n10346), .Y(n10356) );
  NAND2X1 U10771 ( .A(n9346), .B(n9926), .Y(n10354) );
  NAND2X1 U10772 ( .A(n7066), .B(n10361), .Y(n10360) );
  NAND2X1 U10773 ( .A(n10259), .B(n7048), .Y(n10361) );
  NAND2X1 U10774 ( .A(n7048), .B(n9356), .Y(n10359) );
  NAND2X1 U10775 ( .A(n9659), .B(n10260), .Y(n10352) );
  NAND2X1 U10776 ( .A(n9659), .B(n6905), .Y(n10340) );
  INVX1 U10777 ( .A(n7048), .Y(n9659) );
  ADDHXL U10778 ( .A(n10338), .B(n10339), .S(n7048) );
  ADDHXL U10779 ( .A(n9085), .B(n10362), .S(n10338) );
  NOR4X1 U10780 ( .A(n10363), .B(n10364), .C(n10365), .D(n10366), .Y(n10362)
         );
  NOR2X1 U10781 ( .A(n10227), .B(n10346), .Y(n10366) );
  INVX1 U10782 ( .A(G21787), .Y(n10346) );
  NOR2X1 U10783 ( .A(n10271), .B(n9344), .Y(n10365) );
  INVX1 U10784 ( .A(G21628), .Y(n9344) );
  NAND2X1 U10785 ( .A(n10367), .B(n10368), .Y(n10364) );
  NAND2X1 U10786 ( .A(n9346), .B(n10272), .Y(n10368) );
  ADDHXL U10787 ( .A(n10335), .B(n10334), .S(n9346) );
  ADDHXL U10788 ( .A(n10227), .B(n10369), .S(n10335) );
  NOR4X1 U10789 ( .A(n10370), .B(n10371), .C(n10372), .D(n10373), .Y(n10369)
         );
  NOR2X1 U10790 ( .A(n10235), .B(n9345), .Y(n10373) );
  INVX1 U10791 ( .A(G21755), .Y(n9345) );
  NOR2X1 U10792 ( .A(n10234), .B(n10358), .Y(n10372) );
  NAND2X1 U10793 ( .A(n10374), .B(n10375), .Y(n10371) );
  NAND2X1 U10794 ( .A(G21628), .B(n7564), .Y(n10375) );
  NAND2X1 U10795 ( .A(G21723), .B(n10236), .Y(n10374) );
  NOR3X1 U10796 ( .A(n9266), .B(n7049), .C(n7050), .Y(n10370) );
  NOR2X1 U10797 ( .A(n10376), .B(n10377), .Y(n7050) );
  INVX1 U10798 ( .A(n10282), .Y(n7049) );
  NAND2X1 U10799 ( .A(n10377), .B(n10376), .Y(n10282) );
  NAND2X1 U10800 ( .A(n10378), .B(n10379), .Y(n10376) );
  NAND2X1 U10801 ( .A(G21596), .B(n9076), .Y(n10379) );
  NAND2X1 U10802 ( .A(n10380), .B(n8711), .Y(n10378) );
  NAND4X1 U10803 ( .A(n10381), .B(n10382), .C(n10383), .D(n10384), .Y(n10380)
         );
  NOR4X1 U10804 ( .A(n10385), .B(n10386), .C(n10387), .D(n10388), .Y(n10384)
         );
  NOR2X1 U10805 ( .A(n10389), .B(n10311), .Y(n10388) );
  NOR2X1 U10806 ( .A(n10390), .B(n10313), .Y(n10387) );
  NOR2X1 U10807 ( .A(n10391), .B(n10315), .Y(n10386) );
  NOR2X1 U10808 ( .A(n10392), .B(n10317), .Y(n10385) );
  NOR4X1 U10809 ( .A(n10393), .B(n10394), .C(n10395), .D(n10396), .Y(n10383)
         );
  NOR2X1 U10810 ( .A(n10397), .B(n10323), .Y(n10396) );
  NOR2X1 U10811 ( .A(n10398), .B(n10325), .Y(n10395) );
  NOR2X1 U10812 ( .A(n10399), .B(n10327), .Y(n10394) );
  NOR2X1 U10813 ( .A(n10400), .B(n10329), .Y(n10393) );
  NOR4X1 U10814 ( .A(n10401), .B(n10402), .C(n10403), .D(n10404), .Y(n10382)
         );
  NOR2X1 U10815 ( .A(n10405), .B(n10406), .Y(n10404) );
  NOR2X1 U10816 ( .A(n10407), .B(n10408), .Y(n10403) );
  NOR2X1 U10817 ( .A(n10409), .B(n10410), .Y(n10402) );
  NOR2X1 U10818 ( .A(n10411), .B(n10412), .Y(n10401) );
  NOR4X1 U10819 ( .A(n10413), .B(n10414), .C(n10415), .D(n10416), .Y(n10381)
         );
  NOR2X1 U10820 ( .A(n10417), .B(n10418), .Y(n10416) );
  NOR2X1 U10821 ( .A(n10419), .B(n10420), .Y(n10415) );
  NOR2X1 U10822 ( .A(n10421), .B(n10422), .Y(n10414) );
  NOR2X1 U10823 ( .A(n10423), .B(n10424), .Y(n10413) );
  NAND2X1 U10824 ( .A(n10014), .B(n10425), .Y(n10367) );
  NOR2X1 U10825 ( .A(n10426), .B(n10358), .Y(n10363) );
  INVX1 U10826 ( .A(G21596), .Y(n10358) );
  NAND4X1 U10827 ( .A(n10427), .B(n10428), .C(n10429), .D(n10430), .Y(G1017)
         );
  NOR2X1 U10828 ( .A(n10431), .B(n10432), .Y(n10430) );
  NOR2X1 U10829 ( .A(n6891), .B(n9354), .Y(n10432) );
  NOR2X1 U10830 ( .A(n6901), .B(n7062), .Y(n10431) );
  NAND2X1 U10831 ( .A(n7067), .B(n6882), .Y(n10429) );
  NAND2X1 U10832 ( .A(n6903), .B(n7065), .Y(n10428) );
  ADDFXL U10833 ( .A(n9926), .B(n10351), .CI(n10350), .S(n7065) );
  NAND2X1 U10834 ( .A(n10433), .B(n10434), .Y(n10350) );
  NAND2X1 U10835 ( .A(n9926), .B(n10435), .Y(n10434) );
  OR2X1 U10836 ( .A(n10436), .B(n10437), .Y(n10435) );
  NAND2X1 U10837 ( .A(n10437), .B(n10436), .Y(n10433) );
  NAND4X1 U10838 ( .A(n10438), .B(n10439), .C(n10440), .D(n10441), .Y(n10351)
         );
  NOR2X1 U10839 ( .A(n10442), .B(n10443), .Y(n10441) );
  NOR2X1 U10840 ( .A(n10226), .B(n7062), .Y(n10443) );
  NOR2X1 U10841 ( .A(n9908), .B(n9787), .Y(n10442) );
  INVX1 U10842 ( .A(n7067), .Y(n9787) );
  NAND2X1 U10843 ( .A(G21595), .B(n10444), .Y(n10440) );
  NAND2X1 U10844 ( .A(n7066), .B(n10260), .Y(n10439) );
  NAND3X1 U10845 ( .A(n10259), .B(n10256), .C(n9356), .Y(n10438) );
  NAND2X1 U10846 ( .A(n7066), .B(n6905), .Y(n10427) );
  INVX1 U10847 ( .A(n9356), .Y(n7066) );
  NAND2X1 U10848 ( .A(n10445), .B(n10339), .Y(n9356) );
  NAND3X1 U10849 ( .A(n10446), .B(n10447), .C(n10448), .Y(n10339) );
  NAND2X1 U10850 ( .A(n10449), .B(n10450), .Y(n10445) );
  NAND2X1 U10851 ( .A(n10448), .B(n10447), .Y(n10450) );
  INVX1 U10852 ( .A(n10446), .Y(n10449) );
  ADDHXL U10853 ( .A(n9085), .B(n10451), .S(n10446) );
  NOR4X1 U10854 ( .A(n10452), .B(n10453), .C(n10454), .D(n10455), .Y(n10451)
         );
  NOR2X1 U10855 ( .A(n10227), .B(n7062), .Y(n10455) );
  INVX1 U10856 ( .A(G21786), .Y(n7062) );
  NOR2X1 U10857 ( .A(n10271), .B(n9354), .Y(n10454) );
  INVX1 U10858 ( .A(G21627), .Y(n9354) );
  AND2X1 U10859 ( .A(n10456), .B(n10014), .Y(n10453) );
  NAND2X1 U10860 ( .A(n10457), .B(n10458), .Y(n10452) );
  NAND2X1 U10861 ( .A(G21595), .B(n10224), .Y(n10458) );
  NAND2X1 U10862 ( .A(n7067), .B(n10272), .Y(n10457) );
  NOR2X1 U10863 ( .A(n10459), .B(n10334), .Y(n7067) );
  NOR3X1 U10864 ( .A(n10460), .B(n10461), .C(n10462), .Y(n10334) );
  AND2X1 U10865 ( .A(n10460), .B(n10463), .Y(n10459) );
  OR2X1 U10866 ( .A(n10462), .B(n10461), .Y(n10463) );
  ADDHXL U10867 ( .A(n9260), .B(n10464), .S(n10460) );
  NOR3X1 U10868 ( .A(n10465), .B(n10466), .C(n10467), .Y(n10464) );
  NOR2X1 U10869 ( .A(n9266), .B(n7063), .Y(n10467) );
  NAND2X1 U10870 ( .A(n10468), .B(n10469), .Y(n7063) );
  NAND2X1 U10871 ( .A(n10470), .B(n10471), .Y(n10469) );
  INVX1 U10872 ( .A(n10377), .Y(n10468) );
  NOR2X1 U10873 ( .A(n10471), .B(n10470), .Y(n10377) );
  NAND2X1 U10874 ( .A(n10472), .B(n10473), .Y(n10470) );
  NAND2X1 U10875 ( .A(n9076), .B(n7064), .Y(n10473) );
  NAND4X1 U10876 ( .A(n10474), .B(n10475), .C(n10476), .D(n8711), .Y(n10472)
         );
  NOR2X1 U10877 ( .A(n10477), .B(n10478), .Y(n10476) );
  NAND4X1 U10878 ( .A(n10479), .B(n10480), .C(n10481), .D(n10482), .Y(n10478)
         );
  NAND2X1 U10879 ( .A(n10294), .B(G21495), .Y(n10482) );
  INVX1 U10880 ( .A(n10424), .Y(n10294) );
  NAND2X1 U10881 ( .A(n10295), .B(G21503), .Y(n10481) );
  INVX1 U10882 ( .A(n10422), .Y(n10295) );
  NAND2X1 U10883 ( .A(n10296), .B(G21511), .Y(n10480) );
  INVX1 U10884 ( .A(n10420), .Y(n10296) );
  NAND2X1 U10885 ( .A(n10297), .B(G21519), .Y(n10479) );
  INVX1 U10886 ( .A(n10418), .Y(n10297) );
  NAND4X1 U10887 ( .A(n10483), .B(n10484), .C(n10485), .D(n10486), .Y(n10477)
         );
  NAND2X1 U10888 ( .A(n10302), .B(G21527), .Y(n10486) );
  INVX1 U10889 ( .A(n10412), .Y(n10302) );
  NAND2X1 U10890 ( .A(n10303), .B(G21535), .Y(n10485) );
  INVX1 U10891 ( .A(n10410), .Y(n10303) );
  NAND2X1 U10892 ( .A(n10304), .B(G21543), .Y(n10484) );
  INVX1 U10893 ( .A(n10408), .Y(n10304) );
  NAND2X1 U10894 ( .A(n10305), .B(G21551), .Y(n10483) );
  INVX1 U10895 ( .A(n10406), .Y(n10305) );
  NOR4X1 U10896 ( .A(n10487), .B(n10488), .C(n10489), .D(n10490), .Y(n10475)
         );
  NOR2X1 U10897 ( .A(n10491), .B(n10311), .Y(n10490) );
  NOR2X1 U10898 ( .A(n10492), .B(n10313), .Y(n10489) );
  NOR2X1 U10899 ( .A(n10493), .B(n10315), .Y(n10488) );
  NOR2X1 U10900 ( .A(n10494), .B(n10317), .Y(n10487) );
  NOR4X1 U10901 ( .A(n10495), .B(n10496), .C(n10497), .D(n10498), .Y(n10474)
         );
  NOR2X1 U10902 ( .A(n10499), .B(n10323), .Y(n10498) );
  NOR2X1 U10903 ( .A(n10500), .B(n10325), .Y(n10497) );
  NOR2X1 U10904 ( .A(n10501), .B(n10327), .Y(n10496) );
  NOR2X1 U10905 ( .A(n10502), .B(n10329), .Y(n10495) );
  NOR2X1 U10906 ( .A(n10234), .B(n7064), .Y(n10466) );
  INVX1 U10907 ( .A(G21595), .Y(n7064) );
  INVX1 U10908 ( .A(n10503), .Y(n10234) );
  NAND3X1 U10909 ( .A(n10504), .B(n10505), .C(n10506), .Y(n10465) );
  NAND2X1 U10910 ( .A(G21754), .B(n10333), .Y(n10506) );
  NAND2X1 U10911 ( .A(G21627), .B(n7564), .Y(n10505) );
  NAND2X1 U10912 ( .A(G21722), .B(n10236), .Y(n10504) );
  NAND4X1 U10913 ( .A(n10507), .B(n10508), .C(n10509), .D(n10510), .Y(G1016)
         );
  NOR2X1 U10914 ( .A(n10511), .B(n10512), .Y(n10510) );
  NOR2X1 U10915 ( .A(n6891), .B(n9364), .Y(n10512) );
  NOR2X1 U10916 ( .A(n6901), .B(n10513), .Y(n10511) );
  NAND2X1 U10917 ( .A(n9366), .B(n6882), .Y(n10509) );
  NAND2X1 U10918 ( .A(n6903), .B(n7079), .Y(n10508) );
  ADDFXL U10919 ( .A(n9926), .B(n10437), .CI(n10436), .S(n7079) );
  NAND2X1 U10920 ( .A(n10514), .B(n10515), .Y(n10436) );
  NAND2X1 U10921 ( .A(n9926), .B(n10516), .Y(n10515) );
  OR2X1 U10922 ( .A(n10517), .B(n10518), .Y(n10516) );
  NAND2X1 U10923 ( .A(n10518), .B(n10517), .Y(n10514) );
  NAND4X1 U10924 ( .A(n10519), .B(n10520), .C(n10521), .D(n10522), .Y(n10437)
         );
  NOR2X1 U10925 ( .A(n10523), .B(n10524), .Y(n10522) );
  NOR2X1 U10926 ( .A(n10216), .B(n10525), .Y(n10524) );
  NOR2X1 U10927 ( .A(n10226), .B(n10513), .Y(n10523) );
  NAND2X1 U10928 ( .A(n9366), .B(n9926), .Y(n10521) );
  NAND4X1 U10929 ( .A(n10526), .B(n9670), .C(n10256), .D(n10527), .Y(n10520)
         );
  NAND2X1 U10930 ( .A(n9666), .B(n10260), .Y(n10519) );
  NAND2X1 U10931 ( .A(n10217), .B(n10528), .Y(n10260) );
  INVX1 U10932 ( .A(n10259), .Y(n10527) );
  NOR3X1 U10933 ( .A(n7075), .B(n7087), .C(n10529), .Y(n10259) );
  INVX1 U10934 ( .A(n9666), .Y(n7075) );
  NAND2X1 U10935 ( .A(n9666), .B(n6905), .Y(n10507) );
  ADDHXL U10936 ( .A(n10448), .B(n10447), .S(n9666) );
  ADDHXL U10937 ( .A(n9085), .B(n10530), .S(n10447) );
  NOR4X1 U10938 ( .A(n10531), .B(n10532), .C(n10533), .D(n10534), .Y(n10530)
         );
  NOR2X1 U10939 ( .A(n10227), .B(n10513), .Y(n10534) );
  INVX1 U10940 ( .A(G21785), .Y(n10513) );
  NOR2X1 U10941 ( .A(n10271), .B(n9364), .Y(n10533) );
  NAND2X1 U10942 ( .A(n10535), .B(n10536), .Y(n10532) );
  NAND2X1 U10943 ( .A(n9366), .B(n10272), .Y(n10536) );
  ADDHXL U10944 ( .A(n10462), .B(n10461), .S(n9366) );
  ADDHXL U10945 ( .A(n9260), .B(n10537), .S(n10461) );
  NOR4X1 U10946 ( .A(n10538), .B(n10539), .C(n10540), .D(n10541), .Y(n10537)
         );
  AND2X1 U10947 ( .A(n10236), .B(G21721), .Y(n10541) );
  NOR2X1 U10948 ( .A(n9085), .B(n9364), .Y(n10540) );
  INVX1 U10949 ( .A(G21626), .Y(n9364) );
  NOR3X1 U10950 ( .A(n9266), .B(n7076), .C(n7077), .Y(n10539) );
  AND3X1 U10951 ( .A(n10542), .B(n10543), .C(n10544), .Y(n7077) );
  NAND2X1 U10952 ( .A(G21594), .B(n9076), .Y(n10543) );
  NAND2X1 U10953 ( .A(n10545), .B(n8711), .Y(n10542) );
  INVX1 U10954 ( .A(n10471), .Y(n7076) );
  NAND3X1 U10955 ( .A(n10546), .B(n10547), .C(n7088), .Y(n10471) );
  NAND2X1 U10956 ( .A(n9076), .B(n10525), .Y(n10547) );
  OR2X1 U10957 ( .A(n10545), .B(n9076), .Y(n10546) );
  NAND4X1 U10958 ( .A(n10548), .B(n10549), .C(n10550), .D(n10551), .Y(n10545)
         );
  NOR4X1 U10959 ( .A(n10552), .B(n10553), .C(n10554), .D(n10555), .Y(n10551)
         );
  NOR2X1 U10960 ( .A(n10556), .B(n10311), .Y(n10555) );
  NOR2X1 U10961 ( .A(n10557), .B(n10313), .Y(n10554) );
  NOR2X1 U10962 ( .A(n10558), .B(n10315), .Y(n10553) );
  NOR2X1 U10963 ( .A(n10559), .B(n10317), .Y(n10552) );
  NOR4X1 U10964 ( .A(n10560), .B(n10561), .C(n10562), .D(n10563), .Y(n10550)
         );
  NOR2X1 U10965 ( .A(n10564), .B(n10323), .Y(n10563) );
  NOR2X1 U10966 ( .A(n10565), .B(n10325), .Y(n10562) );
  NOR2X1 U10967 ( .A(n10566), .B(n10327), .Y(n10561) );
  NOR2X1 U10968 ( .A(n10567), .B(n10329), .Y(n10560) );
  NOR4X1 U10969 ( .A(n10568), .B(n10569), .C(n10570), .D(n10571), .Y(n10549)
         );
  NOR2X1 U10970 ( .A(n10572), .B(n10406), .Y(n10571) );
  NOR2X1 U10971 ( .A(n10573), .B(n10408), .Y(n10570) );
  NOR2X1 U10972 ( .A(n10574), .B(n10410), .Y(n10569) );
  NOR2X1 U10973 ( .A(n10575), .B(n10412), .Y(n10568) );
  NOR4X1 U10974 ( .A(n10576), .B(n10577), .C(n10578), .D(n10579), .Y(n10548)
         );
  NOR2X1 U10975 ( .A(n10580), .B(n10418), .Y(n10579) );
  NOR2X1 U10976 ( .A(n10581), .B(n10420), .Y(n10578) );
  NOR2X1 U10977 ( .A(n10582), .B(n10422), .Y(n10577) );
  NOR2X1 U10978 ( .A(n10583), .B(n10424), .Y(n10576) );
  NAND2X1 U10979 ( .A(n10584), .B(n10585), .Y(n10538) );
  NAND2X1 U10980 ( .A(G21594), .B(n10503), .Y(n10585) );
  NAND2X1 U10981 ( .A(G21753), .B(n10333), .Y(n10584) );
  NAND2X1 U10982 ( .A(n10014), .B(n10586), .Y(n10535) );
  NOR2X1 U10983 ( .A(n10426), .B(n10525), .Y(n10531) );
  INVX1 U10984 ( .A(G21594), .Y(n10525) );
  NAND4X1 U10985 ( .A(n10587), .B(n10588), .C(n10589), .D(n10590), .Y(G1015)
         );
  NOR2X1 U10986 ( .A(n10591), .B(n10592), .Y(n10590) );
  NOR2X1 U10987 ( .A(n6891), .B(n9374), .Y(n10592) );
  NOR2X1 U10988 ( .A(n6901), .B(n10593), .Y(n10591) );
  NAND2X1 U10989 ( .A(n9376), .B(n6882), .Y(n10589) );
  INVX1 U10990 ( .A(n7090), .Y(n9376) );
  NAND2X1 U10991 ( .A(n6903), .B(n7091), .Y(n10588) );
  ADDFXL U10992 ( .A(n9926), .B(n10518), .CI(n10517), .S(n7091) );
  NAND2X1 U10993 ( .A(n10594), .B(n10595), .Y(n10517) );
  NAND2X1 U10994 ( .A(n9926), .B(n10596), .Y(n10595) );
  OR2X1 U10995 ( .A(n10597), .B(n10598), .Y(n10596) );
  NAND2X1 U10996 ( .A(n10598), .B(n10597), .Y(n10594) );
  NAND4X1 U10997 ( .A(n10599), .B(n10600), .C(n10601), .D(n10602), .Y(n10518)
         );
  NOR2X1 U10998 ( .A(n10603), .B(n10604), .Y(n10602) );
  NOR2X1 U10999 ( .A(n10226), .B(n10593), .Y(n10604) );
  INVX1 U11000 ( .A(G21784), .Y(n10593) );
  NOR2X1 U11001 ( .A(n9908), .B(n7090), .Y(n10603) );
  NAND2X1 U11002 ( .A(G21593), .B(n10444), .Y(n10601) );
  NAND2X1 U11003 ( .A(n9670), .B(n10605), .Y(n10600) );
  NAND3X1 U11004 ( .A(n10526), .B(n10256), .C(n7087), .Y(n10599) );
  INVX1 U11005 ( .A(n9670), .Y(n7087) );
  NAND2X1 U11006 ( .A(n9670), .B(n6905), .Y(n10587) );
  NOR2X1 U11007 ( .A(n10448), .B(n10606), .Y(n9670) );
  AND2X1 U11008 ( .A(n10607), .B(n10608), .Y(n10606) );
  NOR2X1 U11009 ( .A(n10608), .B(n10607), .Y(n10448) );
  ADDHXL U11010 ( .A(n7564), .B(n10609), .S(n10607) );
  NOR3X1 U11011 ( .A(n10610), .B(n10611), .C(n10612), .Y(n10609) );
  NOR2X1 U11012 ( .A(n10613), .B(n7090), .Y(n10612) );
  NAND2X1 U11013 ( .A(n10462), .B(n10614), .Y(n7090) );
  NAND2X1 U11014 ( .A(n10615), .B(n10616), .Y(n10614) );
  OR2X1 U11015 ( .A(n10616), .B(n10615), .Y(n10462) );
  ADDHXL U11016 ( .A(n9260), .B(n10617), .S(n10615) );
  NOR4X1 U11017 ( .A(n10618), .B(n10619), .C(n10620), .D(n10621), .Y(n10617)
         );
  NOR2X1 U11018 ( .A(n9085), .B(n9374), .Y(n10621) );
  INVX1 U11019 ( .A(G21625), .Y(n9374) );
  NOR3X1 U11020 ( .A(n9266), .B(n7088), .C(n7089), .Y(n10620) );
  AND3X1 U11021 ( .A(n10622), .B(n10623), .C(n10624), .Y(n7089) );
  NAND2X1 U11022 ( .A(G21593), .B(n9076), .Y(n10623) );
  NAND2X1 U11023 ( .A(n10625), .B(n8711), .Y(n10622) );
  INVX1 U11024 ( .A(n10544), .Y(n7088) );
  NAND3X1 U11025 ( .A(n10626), .B(n10627), .C(n10628), .Y(n10544) );
  INVX1 U11026 ( .A(n10624), .Y(n10628) );
  NAND2X1 U11027 ( .A(n9076), .B(n10629), .Y(n10627) );
  OR2X1 U11028 ( .A(n10625), .B(n9076), .Y(n10626) );
  NAND4X1 U11029 ( .A(n10630), .B(n10631), .C(n10632), .D(n10633), .Y(n10625)
         );
  NOR4X1 U11030 ( .A(n10634), .B(n10635), .C(n10636), .D(n10637), .Y(n10633)
         );
  NOR2X1 U11031 ( .A(n10638), .B(n10311), .Y(n10637) );
  NOR2X1 U11032 ( .A(n10639), .B(n10313), .Y(n10636) );
  NOR2X1 U11033 ( .A(n10640), .B(n10315), .Y(n10635) );
  NOR2X1 U11034 ( .A(n10641), .B(n10317), .Y(n10634) );
  NOR4X1 U11035 ( .A(n10642), .B(n10643), .C(n10644), .D(n10645), .Y(n10632)
         );
  NOR2X1 U11036 ( .A(n10646), .B(n10323), .Y(n10645) );
  NOR2X1 U11037 ( .A(n10647), .B(n10325), .Y(n10644) );
  NOR2X1 U11038 ( .A(n10648), .B(n10327), .Y(n10643) );
  NOR2X1 U11039 ( .A(n10649), .B(n10329), .Y(n10642) );
  NOR4X1 U11040 ( .A(n10650), .B(n10651), .C(n10652), .D(n10653), .Y(n10631)
         );
  NOR2X1 U11041 ( .A(n10654), .B(n10406), .Y(n10653) );
  NOR2X1 U11042 ( .A(n10655), .B(n10408), .Y(n10652) );
  NOR2X1 U11043 ( .A(n10656), .B(n10410), .Y(n10651) );
  NOR2X1 U11044 ( .A(n10657), .B(n10412), .Y(n10650) );
  NOR4X1 U11045 ( .A(n10658), .B(n10659), .C(n10660), .D(n10661), .Y(n10630)
         );
  NOR2X1 U11046 ( .A(n10662), .B(n10418), .Y(n10661) );
  NOR2X1 U11047 ( .A(n10663), .B(n10420), .Y(n10660) );
  NOR2X1 U11048 ( .A(n10664), .B(n10422), .Y(n10659) );
  NOR2X1 U11049 ( .A(n10665), .B(n10424), .Y(n10658) );
  AND2X1 U11050 ( .A(n10236), .B(G21720), .Y(n10619) );
  NAND2X1 U11051 ( .A(n10666), .B(n10667), .Y(n10618) );
  NAND2X1 U11052 ( .A(G21752), .B(n10333), .Y(n10667) );
  NAND2X1 U11053 ( .A(G21593), .B(n10503), .Y(n10666) );
  OR2X1 U11054 ( .A(n10668), .B(n10669), .Y(n10616) );
  NOR2X1 U11055 ( .A(n10426), .B(n10629), .Y(n10611) );
  INVX1 U11056 ( .A(G21593), .Y(n10629) );
  NAND3X1 U11057 ( .A(n10670), .B(n10671), .C(n10672), .Y(n10610) );
  NAND2X1 U11058 ( .A(n10014), .B(n10673), .Y(n10672) );
  NAND2X1 U11059 ( .A(G21625), .B(n10225), .Y(n10671) );
  NAND2X1 U11060 ( .A(G21784), .B(n9260), .Y(n10670) );
  NAND2X1 U11061 ( .A(n10674), .B(n10675), .Y(n10608) );
  INVX1 U11062 ( .A(n10676), .Y(n10674) );
  NAND4X1 U11063 ( .A(n10677), .B(n10678), .C(n10679), .D(n10680), .Y(G1014)
         );
  NOR2X1 U11064 ( .A(n10681), .B(n10682), .Y(n10680) );
  NOR2X1 U11065 ( .A(n6891), .B(n9384), .Y(n10682) );
  NOR2X1 U11066 ( .A(n6901), .B(n7099), .Y(n10681) );
  NAND2X1 U11067 ( .A(n7104), .B(n6882), .Y(n10679) );
  NAND2X1 U11068 ( .A(n6903), .B(n7102), .Y(n10678) );
  ADDFXL U11069 ( .A(n9926), .B(n10598), .CI(n10597), .S(n7102) );
  NAND2X1 U11070 ( .A(n10683), .B(n10684), .Y(n10597) );
  NAND2X1 U11071 ( .A(n9926), .B(n10685), .Y(n10684) );
  OR2X1 U11072 ( .A(n10686), .B(n10687), .Y(n10685) );
  NAND2X1 U11073 ( .A(n10687), .B(n10686), .Y(n10683) );
  NAND4X1 U11074 ( .A(n10688), .B(n10689), .C(n10690), .D(n10691), .Y(n10598)
         );
  NOR2X1 U11075 ( .A(n10692), .B(n10693), .Y(n10691) );
  NOR2X1 U11076 ( .A(n10216), .B(n7101), .Y(n10693) );
  NOR2X1 U11077 ( .A(n10226), .B(n7099), .Y(n10692) );
  NAND2X1 U11078 ( .A(n7104), .B(n9926), .Y(n10690) );
  NAND4X1 U11079 ( .A(n10694), .B(n9677), .C(n7126), .D(n10529), .Y(n10689) );
  NAND2X1 U11080 ( .A(n7103), .B(n10605), .Y(n10688) );
  NAND2X1 U11081 ( .A(n10217), .B(n10695), .Y(n10605) );
  INVX1 U11082 ( .A(n10526), .Y(n10529) );
  NOR4X1 U11083 ( .A(n10696), .B(n7112), .C(n9386), .D(n9406), .Y(n10526) );
  NAND2X1 U11084 ( .A(n7103), .B(n6905), .Y(n10677) );
  INVX1 U11085 ( .A(n9386), .Y(n7103) );
  ADDHXL U11086 ( .A(n10675), .B(n10676), .S(n9386) );
  ADDHXL U11087 ( .A(n9085), .B(n10697), .S(n10675) );
  NOR4X1 U11088 ( .A(n10698), .B(n10699), .C(n10700), .D(n10701), .Y(n10697)
         );
  NOR2X1 U11089 ( .A(n10227), .B(n7099), .Y(n10701) );
  INVX1 U11090 ( .A(G21783), .Y(n7099) );
  NOR2X1 U11091 ( .A(n10271), .B(n9384), .Y(n10700) );
  NAND2X1 U11092 ( .A(n10702), .B(n10703), .Y(n10699) );
  NAND2X1 U11093 ( .A(n7104), .B(n10272), .Y(n10703) );
  ADDHXL U11094 ( .A(n10668), .B(n10669), .S(n7104) );
  ADDHXL U11095 ( .A(n9260), .B(n10704), .S(n10669) );
  NOR4X1 U11096 ( .A(n10705), .B(n10706), .C(n10707), .D(n10708), .Y(n10704)
         );
  NOR2X1 U11097 ( .A(n9085), .B(n9384), .Y(n10708) );
  INVX1 U11098 ( .A(G21624), .Y(n9384) );
  NOR2X1 U11099 ( .A(n9266), .B(n7100), .Y(n10707) );
  NAND2X1 U11100 ( .A(n10709), .B(n10624), .Y(n7100) );
  NAND4X1 U11101 ( .A(n10710), .B(n10711), .C(n10712), .D(n10713), .Y(n10624)
         );
  NAND2X1 U11102 ( .A(n9076), .B(n7101), .Y(n10713) );
  OR2X1 U11103 ( .A(n10714), .B(n9076), .Y(n10712) );
  NAND3X1 U11104 ( .A(n10715), .B(n10716), .C(n10717), .Y(n10709) );
  NAND2X1 U11105 ( .A(n10710), .B(n10711), .Y(n10717) );
  INVX1 U11106 ( .A(n10718), .Y(n10710) );
  NAND2X1 U11107 ( .A(G21592), .B(n9076), .Y(n10716) );
  NAND2X1 U11108 ( .A(n10714), .B(n8711), .Y(n10715) );
  NAND4X1 U11109 ( .A(n10719), .B(n10720), .C(n10721), .D(n10722), .Y(n10714)
         );
  NOR4X1 U11110 ( .A(n10723), .B(n10724), .C(n10725), .D(n10726), .Y(n10722)
         );
  NOR2X1 U11111 ( .A(n10727), .B(n10311), .Y(n10726) );
  NOR2X1 U11112 ( .A(n10728), .B(n10313), .Y(n10725) );
  NOR2X1 U11113 ( .A(n10729), .B(n10315), .Y(n10724) );
  NOR2X1 U11114 ( .A(n10730), .B(n10317), .Y(n10723) );
  NOR4X1 U11115 ( .A(n10731), .B(n10732), .C(n10733), .D(n10734), .Y(n10721)
         );
  NOR2X1 U11116 ( .A(n10735), .B(n10323), .Y(n10734) );
  NOR2X1 U11117 ( .A(n10736), .B(n10325), .Y(n10733) );
  NOR2X1 U11118 ( .A(n10737), .B(n10327), .Y(n10732) );
  NOR2X1 U11119 ( .A(n10738), .B(n10329), .Y(n10731) );
  NOR4X1 U11120 ( .A(n10739), .B(n10740), .C(n10741), .D(n10742), .Y(n10720)
         );
  NOR2X1 U11121 ( .A(n10743), .B(n10406), .Y(n10742) );
  NOR2X1 U11122 ( .A(n10744), .B(n10408), .Y(n10741) );
  NOR2X1 U11123 ( .A(n10745), .B(n10410), .Y(n10740) );
  NOR2X1 U11124 ( .A(n10746), .B(n10412), .Y(n10739) );
  NOR4X1 U11125 ( .A(n10747), .B(n10748), .C(n10749), .D(n10750), .Y(n10719)
         );
  NOR2X1 U11126 ( .A(n10751), .B(n10418), .Y(n10750) );
  NOR2X1 U11127 ( .A(n10752), .B(n10420), .Y(n10749) );
  NOR2X1 U11128 ( .A(n10753), .B(n10422), .Y(n10748) );
  NOR2X1 U11129 ( .A(n10754), .B(n10424), .Y(n10747) );
  AND2X1 U11130 ( .A(n10236), .B(G21719), .Y(n10706) );
  NAND2X1 U11131 ( .A(n10755), .B(n10756), .Y(n10705) );
  NAND2X1 U11132 ( .A(G21751), .B(n10333), .Y(n10756) );
  NAND2X1 U11133 ( .A(G21592), .B(n10503), .Y(n10755) );
  NAND2X1 U11134 ( .A(n10014), .B(n10757), .Y(n10702) );
  NOR2X1 U11135 ( .A(n10426), .B(n7101), .Y(n10698) );
  INVX1 U11136 ( .A(G21592), .Y(n7101) );
  NAND4X1 U11137 ( .A(n10758), .B(n10759), .C(n10760), .D(n10761), .Y(G1013)
         );
  NOR2X1 U11138 ( .A(n10762), .B(n10763), .Y(n10761) );
  NOR2X1 U11139 ( .A(n6891), .B(n9394), .Y(n10763) );
  NOR2X1 U11140 ( .A(n6901), .B(n10764), .Y(n10762) );
  NAND2X1 U11141 ( .A(n9396), .B(n6882), .Y(n10760) );
  NAND2X1 U11142 ( .A(n6903), .B(n7115), .Y(n10759) );
  ADDFXL U11143 ( .A(n9926), .B(n10687), .CI(n10686), .S(n7115) );
  NAND2X1 U11144 ( .A(n10765), .B(n10766), .Y(n10686) );
  NAND2X1 U11145 ( .A(n9926), .B(n10767), .Y(n10766) );
  OR2X1 U11146 ( .A(n10768), .B(n10769), .Y(n10767) );
  NAND2X1 U11147 ( .A(n10769), .B(n10768), .Y(n10765) );
  NAND4X1 U11148 ( .A(n10770), .B(n10771), .C(n10772), .D(n10773), .Y(n10687)
         );
  NOR2X1 U11149 ( .A(n10774), .B(n10775), .Y(n10773) );
  NOR2X1 U11150 ( .A(n10226), .B(n10764), .Y(n10775) );
  NOR2X1 U11151 ( .A(n9908), .B(n7114), .Y(n10774) );
  NAND2X1 U11152 ( .A(G21591), .B(n10444), .Y(n10772) );
  NAND2X1 U11153 ( .A(n9677), .B(n10776), .Y(n10771) );
  NAND2X1 U11154 ( .A(n10777), .B(n10778), .Y(n10776) );
  INVX1 U11155 ( .A(n10779), .Y(n10777) );
  NAND3X1 U11156 ( .A(n10694), .B(n7126), .C(n7112), .Y(n10770) );
  NAND2X1 U11157 ( .A(n9677), .B(n6905), .Y(n10758) );
  INVX1 U11158 ( .A(n7112), .Y(n9677) );
  NAND2X1 U11159 ( .A(n10676), .B(n10780), .Y(n7112) );
  NAND3X1 U11160 ( .A(n10781), .B(n10782), .C(n10783), .Y(n10780) );
  ADDHXL U11161 ( .A(n10784), .B(n9085), .S(n10783) );
  NAND2X1 U11162 ( .A(n10785), .B(n10786), .Y(n10676) );
  NAND2X1 U11163 ( .A(n10781), .B(n10782), .Y(n10786) );
  NAND2X1 U11164 ( .A(n10787), .B(n10788), .Y(n10781) );
  ADDHXL U11165 ( .A(n7564), .B(n10784), .S(n10785) );
  NAND3X1 U11166 ( .A(n10789), .B(n10790), .C(n10791), .Y(n10784) );
  NOR3X1 U11167 ( .A(n10792), .B(n10793), .C(n10794), .Y(n10791) );
  NOR2X1 U11168 ( .A(n10227), .B(n10764), .Y(n10794) );
  INVX1 U11169 ( .A(G21782), .Y(n10764) );
  NOR2X1 U11170 ( .A(n10271), .B(n9394), .Y(n10793) );
  AND2X1 U11171 ( .A(n10795), .B(n10014), .Y(n10792) );
  NAND2X1 U11172 ( .A(G21591), .B(n10224), .Y(n10790) );
  NAND2X1 U11173 ( .A(n9396), .B(n10272), .Y(n10789) );
  INVX1 U11174 ( .A(n7114), .Y(n9396) );
  NAND2X1 U11175 ( .A(n10668), .B(n10796), .Y(n7114) );
  NAND2X1 U11176 ( .A(n10797), .B(n10798), .Y(n10796) );
  OR2X1 U11177 ( .A(n10798), .B(n10797), .Y(n10668) );
  ADDHXL U11178 ( .A(n10799), .B(n10227), .S(n10797) );
  NAND4X1 U11179 ( .A(n10800), .B(n10801), .C(n10802), .D(n10803), .Y(n10799)
         );
  NAND2X1 U11180 ( .A(G21718), .B(n10236), .Y(n10803) );
  NOR2X1 U11181 ( .A(n10804), .B(n10805), .Y(n10802) );
  NOR2X1 U11182 ( .A(n9085), .B(n9394), .Y(n10805) );
  INVX1 U11183 ( .A(G21623), .Y(n9394) );
  NOR2X1 U11184 ( .A(n7113), .B(n9266), .Y(n10804) );
  ADDHXL U11185 ( .A(n10718), .B(n10711), .S(n7113) );
  NAND2X1 U11186 ( .A(n10806), .B(n10807), .Y(n10711) );
  NAND2X1 U11187 ( .A(G21591), .B(n9076), .Y(n10807) );
  NAND2X1 U11188 ( .A(n10808), .B(n8711), .Y(n10806) );
  NAND4X1 U11189 ( .A(n10809), .B(n10810), .C(n10811), .D(n10812), .Y(n10808)
         );
  NOR4X1 U11190 ( .A(n10813), .B(n10814), .C(n10815), .D(n10816), .Y(n10812)
         );
  NOR2X1 U11191 ( .A(n10817), .B(n10311), .Y(n10816) );
  NOR2X1 U11192 ( .A(n10818), .B(n10313), .Y(n10815) );
  NOR2X1 U11193 ( .A(n10819), .B(n10315), .Y(n10814) );
  NOR2X1 U11194 ( .A(n10820), .B(n10317), .Y(n10813) );
  NOR4X1 U11195 ( .A(n10821), .B(n10822), .C(n10823), .D(n10824), .Y(n10811)
         );
  NOR2X1 U11196 ( .A(n10825), .B(n10323), .Y(n10824) );
  NOR2X1 U11197 ( .A(n10826), .B(n10325), .Y(n10823) );
  NOR2X1 U11198 ( .A(n10827), .B(n10327), .Y(n10822) );
  NOR2X1 U11199 ( .A(n10828), .B(n10329), .Y(n10821) );
  NOR4X1 U11200 ( .A(n10829), .B(n10830), .C(n10831), .D(n10832), .Y(n10810)
         );
  NOR2X1 U11201 ( .A(n10833), .B(n10406), .Y(n10832) );
  NOR2X1 U11202 ( .A(n10834), .B(n10408), .Y(n10831) );
  NOR2X1 U11203 ( .A(n10835), .B(n10410), .Y(n10830) );
  NOR2X1 U11204 ( .A(n10836), .B(n10412), .Y(n10829) );
  NOR4X1 U11205 ( .A(n10837), .B(n10838), .C(n10839), .D(n10840), .Y(n10809)
         );
  NOR2X1 U11206 ( .A(n10841), .B(n10418), .Y(n10840) );
  NOR2X1 U11207 ( .A(n10842), .B(n10420), .Y(n10839) );
  NOR2X1 U11208 ( .A(n10843), .B(n10422), .Y(n10838) );
  NOR2X1 U11209 ( .A(n10844), .B(n10424), .Y(n10837) );
  NAND2X1 U11210 ( .A(n10845), .B(n10846), .Y(n10718) );
  NAND2X1 U11211 ( .A(G21750), .B(n10333), .Y(n10801) );
  NAND2X1 U11212 ( .A(G21591), .B(n10503), .Y(n10800) );
  OR2X1 U11213 ( .A(n10847), .B(n10848), .Y(n10798) );
  NAND4X1 U11214 ( .A(n10849), .B(n10850), .C(n10851), .D(n10852), .Y(G1012)
         );
  NOR2X1 U11215 ( .A(n10853), .B(n10854), .Y(n10852) );
  NOR2X1 U11216 ( .A(n6891), .B(n9404), .Y(n10854) );
  NOR2X1 U11217 ( .A(n6901), .B(n7123), .Y(n10853) );
  NAND2X1 U11218 ( .A(n7127), .B(n6882), .Y(n10851) );
  NAND2X1 U11219 ( .A(n6903), .B(n7125), .Y(n10850) );
  ADDFXL U11220 ( .A(n9926), .B(n10769), .CI(n10768), .S(n7125) );
  NAND2X1 U11221 ( .A(n10855), .B(n10856), .Y(n10768) );
  NAND2X1 U11222 ( .A(n9926), .B(n10857), .Y(n10856) );
  OR2X1 U11223 ( .A(n10858), .B(n10859), .Y(n10857) );
  NAND2X1 U11224 ( .A(n10859), .B(n10858), .Y(n10855) );
  NAND4X1 U11225 ( .A(n10860), .B(n10861), .C(n10862), .D(n10863), .Y(n10769)
         );
  NOR2X1 U11226 ( .A(n10864), .B(n10865), .Y(n10863) );
  NOR2X1 U11227 ( .A(n10226), .B(n7123), .Y(n10865) );
  NOR2X1 U11228 ( .A(n9908), .B(n9823), .Y(n10864) );
  INVX1 U11229 ( .A(n7127), .Y(n9823) );
  NAND2X1 U11230 ( .A(G21590), .B(n10444), .Y(n10862) );
  NAND2X1 U11231 ( .A(n10694), .B(n9406), .Y(n10861) );
  NOR2X1 U11232 ( .A(n10696), .B(n9192), .Y(n10694) );
  NAND2X1 U11233 ( .A(n7126), .B(n10779), .Y(n10860) );
  NAND2X1 U11234 ( .A(n7126), .B(n6905), .Y(n10849) );
  INVX1 U11235 ( .A(n9406), .Y(n7126) );
  ADDHXL U11236 ( .A(n10866), .B(n10788), .S(n9406) );
  NAND2X1 U11237 ( .A(n10867), .B(n10868), .Y(n10788) );
  NAND2X1 U11238 ( .A(n10869), .B(n10870), .Y(n10868) );
  NAND3X1 U11239 ( .A(n10014), .B(n10871), .C(n10872), .Y(n10867) );
  ADDHXL U11240 ( .A(n7564), .B(n10873), .S(n10872) );
  NAND2X1 U11241 ( .A(n10782), .B(n10787), .Y(n10866) );
  NAND2X1 U11242 ( .A(n10874), .B(n10875), .Y(n10787) );
  NAND2X1 U11243 ( .A(n10014), .B(n10876), .Y(n10875) );
  ADDHXL U11244 ( .A(n7564), .B(n10877), .S(n10874) );
  NAND3X1 U11245 ( .A(n10878), .B(n10876), .C(n10014), .Y(n10782) );
  NAND2X1 U11246 ( .A(n10877), .B(n9085), .Y(n10878) );
  AND4X1 U11247 ( .A(n10879), .B(n10880), .C(n10881), .D(n10882), .Y(n10877)
         );
  NOR2X1 U11248 ( .A(n10883), .B(n10884), .Y(n10882) );
  NOR2X1 U11249 ( .A(n10227), .B(n7123), .Y(n10884) );
  INVX1 U11250 ( .A(G21781), .Y(n7123) );
  NOR2X1 U11251 ( .A(n10271), .B(n9404), .Y(n10883) );
  NAND2X1 U11252 ( .A(G21590), .B(n10224), .Y(n10881) );
  NAND2X1 U11253 ( .A(n7127), .B(n10272), .Y(n10880) );
  ADDHXL U11254 ( .A(n10847), .B(n10848), .S(n7127) );
  ADDHXL U11255 ( .A(n10885), .B(n10227), .S(n10848) );
  NAND3X1 U11256 ( .A(n10886), .B(n10887), .C(n10888), .Y(n10885) );
  NOR3X1 U11257 ( .A(n10889), .B(n10890), .C(n10891), .Y(n10888) );
  NOR2X1 U11258 ( .A(n9085), .B(n9404), .Y(n10891) );
  INVX1 U11259 ( .A(G21622), .Y(n9404) );
  NOR2X1 U11260 ( .A(n7124), .B(n9266), .Y(n10890) );
  INVX1 U11261 ( .A(n10892), .Y(n7124) );
  ADDHXL U11262 ( .A(n10845), .B(n10846), .S(n10892) );
  NAND2X1 U11263 ( .A(n10893), .B(n10894), .Y(n10846) );
  NAND2X1 U11264 ( .A(G21590), .B(n9076), .Y(n10894) );
  NAND2X1 U11265 ( .A(n10895), .B(n8711), .Y(n10893) );
  NAND4X1 U11266 ( .A(n10896), .B(n10897), .C(n10898), .D(n10899), .Y(n10895)
         );
  NOR4X1 U11267 ( .A(n10900), .B(n10901), .C(n10902), .D(n10903), .Y(n10899)
         );
  NOR2X1 U11268 ( .A(n10904), .B(n10311), .Y(n10903) );
  NAND2X1 U11269 ( .A(n10905), .B(n10906), .Y(n10311) );
  NOR2X1 U11270 ( .A(n10907), .B(n10313), .Y(n10902) );
  NAND2X1 U11271 ( .A(n10905), .B(n10908), .Y(n10313) );
  NOR2X1 U11272 ( .A(n10909), .B(n10315), .Y(n10901) );
  NAND2X1 U11273 ( .A(n10906), .B(n10910), .Y(n10315) );
  NOR2X1 U11274 ( .A(n10911), .B(n10317), .Y(n10900) );
  NAND2X1 U11275 ( .A(n10910), .B(n10908), .Y(n10317) );
  NOR4X1 U11276 ( .A(n10912), .B(n10913), .C(n10914), .D(n10915), .Y(n10898)
         );
  NOR2X1 U11277 ( .A(n10916), .B(n10323), .Y(n10915) );
  NAND2X1 U11278 ( .A(n10917), .B(n10906), .Y(n10323) );
  NOR2X1 U11279 ( .A(n10918), .B(n10325), .Y(n10914) );
  NAND2X1 U11280 ( .A(n10917), .B(n10908), .Y(n10325) );
  NOR2X1 U11281 ( .A(n10919), .B(n10327), .Y(n10913) );
  NAND2X1 U11282 ( .A(n10920), .B(n10906), .Y(n10327) );
  NOR2X1 U11283 ( .A(n8890), .B(n10921), .Y(n10906) );
  NOR2X1 U11284 ( .A(n10922), .B(n10329), .Y(n10912) );
  NAND2X1 U11285 ( .A(n10920), .B(n10908), .Y(n10329) );
  NOR2X1 U11286 ( .A(G21561), .B(n10921), .Y(n10908) );
  NOR4X1 U11287 ( .A(n10923), .B(n10924), .C(n10925), .D(n10926), .Y(n10897)
         );
  NOR2X1 U11288 ( .A(n10927), .B(n10406), .Y(n10926) );
  NAND2X1 U11289 ( .A(n10928), .B(n10920), .Y(n10406) );
  NOR2X1 U11290 ( .A(n10929), .B(n10408), .Y(n10925) );
  NAND2X1 U11291 ( .A(n10930), .B(n10920), .Y(n10408) );
  NOR2X1 U11292 ( .A(n9136), .B(n9158), .Y(n10920) );
  NOR2X1 U11293 ( .A(n10931), .B(n10410), .Y(n10924) );
  NAND2X1 U11294 ( .A(n10928), .B(n10917), .Y(n10410) );
  NOR2X1 U11295 ( .A(n10932), .B(n10412), .Y(n10923) );
  NAND2X1 U11296 ( .A(n10930), .B(n10917), .Y(n10412) );
  NOR2X1 U11297 ( .A(n9158), .B(n10933), .Y(n10917) );
  INVX1 U11298 ( .A(n10934), .Y(n9158) );
  NOR4X1 U11299 ( .A(n10935), .B(n10936), .C(n10937), .D(n10938), .Y(n10896)
         );
  NOR2X1 U11300 ( .A(n10939), .B(n10418), .Y(n10938) );
  NAND2X1 U11301 ( .A(n10928), .B(n10910), .Y(n10418) );
  NOR2X1 U11302 ( .A(n10940), .B(n10420), .Y(n10937) );
  NAND2X1 U11303 ( .A(n10930), .B(n10910), .Y(n10420) );
  NOR2X1 U11304 ( .A(n9136), .B(n10934), .Y(n10910) );
  INVX1 U11305 ( .A(n10933), .Y(n9136) );
  NOR2X1 U11306 ( .A(n10941), .B(n10422), .Y(n10936) );
  NAND2X1 U11307 ( .A(n10928), .B(n10905), .Y(n10422) );
  NOR2X1 U11308 ( .A(n9204), .B(G21561), .Y(n10928) );
  NOR2X1 U11309 ( .A(n10942), .B(n10424), .Y(n10935) );
  NAND2X1 U11310 ( .A(n10930), .B(n10905), .Y(n10424) );
  NOR2X1 U11311 ( .A(n10934), .B(n10933), .Y(n10905) );
  NOR2X1 U11312 ( .A(n10943), .B(n10944), .Y(n10933) );
  NOR2X1 U11313 ( .A(n10945), .B(n9076), .Y(n10943) );
  ADDHXL U11314 ( .A(n8893), .B(n10946), .S(n10934) );
  NOR2X1 U11315 ( .A(n9204), .B(n8890), .Y(n10930) );
  INVX1 U11316 ( .A(n10921), .Y(n9204) );
  NOR2X1 U11317 ( .A(n10947), .B(n10948), .Y(n10921) );
  NOR3X1 U11318 ( .A(n10949), .B(G21559), .C(n10950), .Y(n10948) );
  INVX1 U11319 ( .A(n10946), .Y(n10950) );
  AND2X1 U11320 ( .A(n8870), .B(n10951), .Y(n10947) );
  NAND2X1 U11321 ( .A(n10949), .B(n10946), .Y(n10951) );
  NAND2X1 U11322 ( .A(n9076), .B(n10952), .Y(n10946) );
  NAND2X1 U11323 ( .A(n10953), .B(n10954), .Y(n10845) );
  NAND2X1 U11324 ( .A(n10955), .B(G21589), .Y(n10954) );
  NAND2X1 U11325 ( .A(n10336), .B(n8711), .Y(n10953) );
  NAND4X1 U11326 ( .A(n10956), .B(n10957), .C(n10958), .D(n10959), .Y(n10336)
         );
  NOR4X1 U11327 ( .A(n10960), .B(n10961), .C(n10962), .D(n10963), .Y(n10959)
         );
  NOR2X1 U11328 ( .A(n10964), .B(n7597), .Y(n10963) );
  NOR2X1 U11329 ( .A(n10965), .B(n7677), .Y(n10962) );
  NOR2X1 U11330 ( .A(n10966), .B(n7757), .Y(n10961) );
  NOR2X1 U11331 ( .A(n10967), .B(n7919), .Y(n10960) );
  NOR4X1 U11332 ( .A(n10968), .B(n10969), .C(n10970), .D(n10971), .Y(n10958)
         );
  NOR2X1 U11333 ( .A(n10972), .B(n7997), .Y(n10971) );
  NOR2X1 U11334 ( .A(n10973), .B(n8075), .Y(n10970) );
  NOR2X1 U11335 ( .A(n10326), .B(n8234), .Y(n10969) );
  NOR2X1 U11336 ( .A(n10324), .B(n8312), .Y(n10968) );
  NOR4X1 U11337 ( .A(n10974), .B(n10975), .C(n10976), .D(n10977), .Y(n10957)
         );
  NOR2X1 U11338 ( .A(n10322), .B(n8390), .Y(n10977) );
  NOR2X1 U11339 ( .A(n10314), .B(n8551), .Y(n10976) );
  NOR2X1 U11340 ( .A(n10312), .B(n8629), .Y(n10975) );
  NOR2X1 U11341 ( .A(n10310), .B(n8706), .Y(n10974) );
  NOR4X1 U11342 ( .A(n10978), .B(n10979), .C(n10980), .D(n10981), .Y(n10956)
         );
  NOR2X1 U11343 ( .A(n10982), .B(n7487), .Y(n10981) );
  NOR2X1 U11344 ( .A(n10983), .B(n7839), .Y(n10980) );
  NOR2X1 U11345 ( .A(n10328), .B(n8154), .Y(n10979) );
  NOR2X1 U11346 ( .A(n10316), .B(n8469), .Y(n10978) );
  AND2X1 U11347 ( .A(n10236), .B(G21717), .Y(n10889) );
  NAND2X1 U11348 ( .A(G21749), .B(n10333), .Y(n10887) );
  NAND2X1 U11349 ( .A(G21590), .B(n10503), .Y(n10886) );
  NAND2X1 U11350 ( .A(n10014), .B(n10984), .Y(n10879) );
  NAND4X1 U11351 ( .A(n10985), .B(n10986), .C(n10987), .D(n10988), .Y(G1011)
         );
  NOR2X1 U11352 ( .A(n10989), .B(n10990), .Y(n10988) );
  NOR2X1 U11353 ( .A(n6891), .B(n9414), .Y(n10990) );
  NOR2X1 U11354 ( .A(n6901), .B(n7135), .Y(n10989) );
  NAND2X1 U11355 ( .A(n7140), .B(n6882), .Y(n10987) );
  NAND2X1 U11356 ( .A(n6903), .B(n7138), .Y(n10986) );
  ADDFXL U11357 ( .A(n9926), .B(n10859), .CI(n10858), .S(n7138) );
  NAND2X1 U11358 ( .A(n10991), .B(n10992), .Y(n10858) );
  NAND2X1 U11359 ( .A(n9926), .B(n10993), .Y(n10992) );
  OR2X1 U11360 ( .A(n10994), .B(n10995), .Y(n10993) );
  NAND2X1 U11361 ( .A(n10995), .B(n10994), .Y(n10991) );
  NAND4X1 U11362 ( .A(n10996), .B(n10997), .C(n10998), .D(n10999), .Y(n10859)
         );
  NOR2X1 U11363 ( .A(n11000), .B(n11001), .Y(n10999) );
  NOR2X1 U11364 ( .A(n10216), .B(n7137), .Y(n11001) );
  INVX1 U11365 ( .A(G21589), .Y(n7137) );
  NOR2X1 U11366 ( .A(n10226), .B(n7135), .Y(n11000) );
  INVX1 U11367 ( .A(G21780), .Y(n7135) );
  NAND2X1 U11368 ( .A(n7140), .B(n9926), .Y(n10998) );
  NAND4X1 U11369 ( .A(n7152), .B(n11002), .C(n7164), .D(n10696), .Y(n10997) );
  NAND2X1 U11370 ( .A(n7139), .B(n10779), .Y(n10996) );
  NAND2X1 U11371 ( .A(n10217), .B(n11003), .Y(n10779) );
  OR4X1 U11372 ( .A(n9416), .B(n11004), .C(n9426), .D(n9436), .Y(n10696) );
  INVX1 U11373 ( .A(n7139), .Y(n9416) );
  NAND2X1 U11374 ( .A(n7139), .B(n6905), .Y(n10985) );
  ADDHXL U11375 ( .A(n10870), .B(n10869), .S(n7139) );
  NAND2X1 U11376 ( .A(n11005), .B(n11006), .Y(n10869) );
  NAND2X1 U11377 ( .A(n10014), .B(n10871), .Y(n11006) );
  ADDHXL U11378 ( .A(n10873), .B(n9085), .S(n11005) );
  NAND4X1 U11379 ( .A(n11007), .B(n11008), .C(n11009), .D(n11010), .Y(n10873)
         );
  NAND2X1 U11380 ( .A(G21589), .B(n10224), .Y(n11010) );
  NAND2X1 U11381 ( .A(G21780), .B(n9260), .Y(n11009) );
  NAND2X1 U11382 ( .A(n7140), .B(n10272), .Y(n11008) );
  INVX1 U11383 ( .A(n9831), .Y(n7140) );
  NAND2X1 U11384 ( .A(n10847), .B(n11011), .Y(n9831) );
  NAND2X1 U11385 ( .A(n11012), .B(n11013), .Y(n11011) );
  OR2X1 U11386 ( .A(n11013), .B(n11012), .Y(n10847) );
  ADDHXL U11387 ( .A(n11014), .B(n10227), .S(n11012) );
  NAND3X1 U11388 ( .A(n11015), .B(n11016), .C(n11017), .Y(n11014) );
  NOR3X1 U11389 ( .A(n11018), .B(n11019), .C(n11020), .Y(n11017) );
  AND2X1 U11390 ( .A(n10236), .B(G21716), .Y(n11020) );
  NOR2X1 U11391 ( .A(n9085), .B(n9414), .Y(n11019) );
  INVX1 U11392 ( .A(G21621), .Y(n9414) );
  NOR2X1 U11393 ( .A(n7136), .B(n9266), .Y(n11018) );
  AND2X1 U11394 ( .A(n11021), .B(n11022), .Y(n7136) );
  NAND2X1 U11395 ( .A(n10425), .B(n8711), .Y(n11022) );
  NAND4X1 U11396 ( .A(n11023), .B(n11024), .C(n11025), .D(n11026), .Y(n10425)
         );
  NOR4X1 U11397 ( .A(n11027), .B(n11028), .C(n11029), .D(n11030), .Y(n11026)
         );
  NOR2X1 U11398 ( .A(n10407), .B(n7597), .Y(n11030) );
  NOR2X1 U11399 ( .A(n10409), .B(n7677), .Y(n11029) );
  NOR2X1 U11400 ( .A(n10411), .B(n7757), .Y(n11028) );
  NOR2X1 U11401 ( .A(n10419), .B(n7919), .Y(n11027) );
  NOR4X1 U11402 ( .A(n11031), .B(n11032), .C(n11033), .D(n11034), .Y(n11025)
         );
  NOR2X1 U11403 ( .A(n10421), .B(n7997), .Y(n11034) );
  NOR2X1 U11404 ( .A(n10423), .B(n8075), .Y(n11033) );
  NOR2X1 U11405 ( .A(n10399), .B(n8234), .Y(n11032) );
  NOR2X1 U11406 ( .A(n10398), .B(n8312), .Y(n11031) );
  NOR4X1 U11407 ( .A(n11035), .B(n11036), .C(n11037), .D(n11038), .Y(n11024)
         );
  NOR2X1 U11408 ( .A(n10397), .B(n8390), .Y(n11038) );
  NOR2X1 U11409 ( .A(n10391), .B(n8551), .Y(n11037) );
  NOR2X1 U11410 ( .A(n10390), .B(n8629), .Y(n11036) );
  NOR2X1 U11411 ( .A(n10389), .B(n8706), .Y(n11035) );
  NOR4X1 U11412 ( .A(n11039), .B(n11040), .C(n11041), .D(n11042), .Y(n11023)
         );
  NOR2X1 U11413 ( .A(n10405), .B(n7487), .Y(n11042) );
  NOR2X1 U11414 ( .A(n10417), .B(n7839), .Y(n11041) );
  NOR2X1 U11415 ( .A(n10400), .B(n8154), .Y(n11040) );
  NOR2X1 U11416 ( .A(n10392), .B(n8469), .Y(n11039) );
  NAND2X1 U11417 ( .A(n11043), .B(n9076), .Y(n11021) );
  ADDHXL U11418 ( .A(G21589), .B(n10955), .S(n11043) );
  NOR2X1 U11419 ( .A(n11044), .B(n7150), .Y(n10955) );
  INVX1 U11420 ( .A(G21588), .Y(n7150) );
  NAND2X1 U11421 ( .A(G21589), .B(n10503), .Y(n11016) );
  NAND2X1 U11422 ( .A(G21748), .B(n10333), .Y(n11015) );
  OR2X1 U11423 ( .A(n11045), .B(n11046), .Y(n11013) );
  NAND2X1 U11424 ( .A(G21621), .B(n10225), .Y(n11007) );
  AND2X1 U11425 ( .A(n11047), .B(n11048), .Y(n10870) );
  NAND4X1 U11426 ( .A(n11049), .B(n11050), .C(n11051), .D(n11052), .Y(G1010)
         );
  NOR2X1 U11427 ( .A(n11053), .B(n11054), .Y(n11052) );
  NOR2X1 U11428 ( .A(n6891), .B(n9424), .Y(n11054) );
  NOR2X1 U11429 ( .A(n6901), .B(n7148), .Y(n11053) );
  NAND2X1 U11430 ( .A(n7153), .B(n6882), .Y(n11051) );
  NAND2X1 U11431 ( .A(n6903), .B(n7151), .Y(n11050) );
  ADDFXL U11432 ( .A(n9926), .B(n10995), .CI(n10994), .S(n7151) );
  NAND2X1 U11433 ( .A(n11055), .B(n11056), .Y(n10994) );
  NAND2X1 U11434 ( .A(n9926), .B(n11057), .Y(n11056) );
  OR2X1 U11435 ( .A(n11058), .B(n11059), .Y(n11057) );
  NAND2X1 U11436 ( .A(n11059), .B(n11058), .Y(n11055) );
  NAND4X1 U11437 ( .A(n11060), .B(n11061), .C(n11062), .D(n11063), .Y(n10995)
         );
  NOR2X1 U11438 ( .A(n11064), .B(n11065), .Y(n11063) );
  NOR2X1 U11439 ( .A(n10226), .B(n7148), .Y(n11065) );
  INVX1 U11440 ( .A(G21779), .Y(n7148) );
  NOR2X1 U11441 ( .A(n9908), .B(n9839), .Y(n11064) );
  INVX1 U11442 ( .A(n7153), .Y(n9839) );
  NAND2X1 U11443 ( .A(G21588), .B(n10444), .Y(n11062) );
  NAND2X1 U11444 ( .A(n7152), .B(n11066), .Y(n11061) );
  NAND2X1 U11445 ( .A(n11067), .B(n11068), .Y(n11066) );
  INVX1 U11446 ( .A(n11069), .Y(n11067) );
  NAND3X1 U11447 ( .A(n11002), .B(n7164), .C(n9426), .Y(n11060) );
  INVX1 U11448 ( .A(n7152), .Y(n9426) );
  NAND2X1 U11449 ( .A(n7152), .B(n6905), .Y(n11049) );
  ADDHXL U11450 ( .A(n11048), .B(n11047), .S(n7152) );
  NAND2X1 U11451 ( .A(n11070), .B(n11071), .Y(n11047) );
  NAND2X1 U11452 ( .A(n10014), .B(n11072), .Y(n11071) );
  ADDHXL U11453 ( .A(n9085), .B(n11073), .S(n11070) );
  NAND4X1 U11454 ( .A(n11074), .B(n11075), .C(n11076), .D(n11077), .Y(n11073)
         );
  NAND2X1 U11455 ( .A(n7153), .B(n10272), .Y(n11077) );
  ADDHXL U11456 ( .A(n11045), .B(n11046), .S(n7153) );
  ADDHXL U11457 ( .A(n11078), .B(n10227), .S(n11046) );
  NAND3X1 U11458 ( .A(n11079), .B(n11080), .C(n11081), .Y(n11078) );
  NOR3X1 U11459 ( .A(n11082), .B(n11083), .C(n11084), .Y(n11081) );
  AND2X1 U11460 ( .A(n10236), .B(G21715), .Y(n11084) );
  NOR2X1 U11461 ( .A(n9085), .B(n9424), .Y(n11083) );
  INVX1 U11462 ( .A(G21620), .Y(n9424) );
  NOR2X1 U11463 ( .A(n7149), .B(n9266), .Y(n11082) );
  AND3X1 U11464 ( .A(n11085), .B(n11086), .C(n11087), .Y(n7149) );
  OR2X1 U11465 ( .A(n11044), .B(G21588), .Y(n11087) );
  NAND3X1 U11466 ( .A(G21588), .B(n11044), .C(n9076), .Y(n11086) );
  NAND2X1 U11467 ( .A(n11088), .B(G21587), .Y(n11044) );
  NAND2X1 U11468 ( .A(n10456), .B(n8711), .Y(n11085) );
  NAND4X1 U11469 ( .A(n11089), .B(n11090), .C(n11091), .D(n11092), .Y(n10456)
         );
  NOR4X1 U11470 ( .A(n11093), .B(n11094), .C(n11095), .D(n11096), .Y(n11092)
         );
  NOR2X1 U11471 ( .A(n11097), .B(n7597), .Y(n11096) );
  NOR2X1 U11472 ( .A(n11098), .B(n7677), .Y(n11095) );
  NOR2X1 U11473 ( .A(n11099), .B(n7757), .Y(n11094) );
  NOR2X1 U11474 ( .A(n11100), .B(n7919), .Y(n11093) );
  NOR4X1 U11475 ( .A(n11101), .B(n11102), .C(n11103), .D(n11104), .Y(n11091)
         );
  NOR2X1 U11476 ( .A(n11105), .B(n7997), .Y(n11104) );
  NOR2X1 U11477 ( .A(n11106), .B(n8075), .Y(n11103) );
  NOR2X1 U11478 ( .A(n10501), .B(n8234), .Y(n11102) );
  NOR2X1 U11479 ( .A(n10500), .B(n8312), .Y(n11101) );
  NOR4X1 U11480 ( .A(n11107), .B(n11108), .C(n11109), .D(n11110), .Y(n11090)
         );
  NOR2X1 U11481 ( .A(n10499), .B(n8390), .Y(n11110) );
  NOR2X1 U11482 ( .A(n10493), .B(n8551), .Y(n11109) );
  NOR2X1 U11483 ( .A(n10492), .B(n8629), .Y(n11108) );
  NOR2X1 U11484 ( .A(n10491), .B(n8706), .Y(n11107) );
  NOR4X1 U11485 ( .A(n11111), .B(n11112), .C(n11113), .D(n11114), .Y(n11089)
         );
  NOR2X1 U11486 ( .A(n11115), .B(n7487), .Y(n11114) );
  NOR2X1 U11487 ( .A(n11116), .B(n7839), .Y(n11113) );
  NOR2X1 U11488 ( .A(n10502), .B(n8154), .Y(n11112) );
  NOR2X1 U11489 ( .A(n10494), .B(n8469), .Y(n11111) );
  NAND2X1 U11490 ( .A(G21588), .B(n10503), .Y(n11080) );
  NAND2X1 U11491 ( .A(G21747), .B(n10333), .Y(n11079) );
  NAND2X1 U11492 ( .A(G21588), .B(n10224), .Y(n11076) );
  NAND2X1 U11493 ( .A(G21620), .B(n10225), .Y(n11075) );
  NAND2X1 U11494 ( .A(G21779), .B(n9260), .Y(n11074) );
  NAND2X1 U11495 ( .A(n11117), .B(n11118), .Y(n11048) );
  NAND2X1 U11496 ( .A(n11119), .B(n11120), .Y(n11118) );
  NAND3X1 U11497 ( .A(n11121), .B(n11122), .C(n10014), .Y(n11117) );
  OR2X1 U11498 ( .A(n11123), .B(n7564), .Y(n11121) );
  NAND4X1 U11499 ( .A(n11124), .B(n11125), .C(n11126), .D(n11127), .Y(G1009)
         );
  NOR2X1 U11500 ( .A(n11128), .B(n11129), .Y(n11127) );
  NOR2X1 U11501 ( .A(n6891), .B(n9434), .Y(n11129) );
  NOR2X1 U11502 ( .A(n6901), .B(n7161), .Y(n11128) );
  NAND2X1 U11503 ( .A(n7165), .B(n6882), .Y(n11126) );
  NAND2X1 U11504 ( .A(n6903), .B(n7163), .Y(n11125) );
  ADDFXL U11505 ( .A(n9926), .B(n11059), .CI(n11058), .S(n7163) );
  NAND2X1 U11506 ( .A(n11130), .B(n11131), .Y(n11058) );
  NAND2X1 U11507 ( .A(n9926), .B(n11132), .Y(n11131) );
  OR2X1 U11508 ( .A(n11133), .B(n11134), .Y(n11132) );
  NAND2X1 U11509 ( .A(n11134), .B(n11133), .Y(n11130) );
  NAND4X1 U11510 ( .A(n11135), .B(n11136), .C(n11137), .D(n11138), .Y(n11059)
         );
  NOR2X1 U11511 ( .A(n11139), .B(n11140), .Y(n11138) );
  NOR2X1 U11512 ( .A(n10226), .B(n7161), .Y(n11140) );
  INVX1 U11513 ( .A(G21778), .Y(n7161) );
  NOR2X1 U11514 ( .A(n9908), .B(n9847), .Y(n11139) );
  NAND2X1 U11515 ( .A(G21587), .B(n10444), .Y(n11137) );
  NAND2X1 U11516 ( .A(n9436), .B(n11002), .Y(n11136) );
  NOR2X1 U11517 ( .A(n11004), .B(n9192), .Y(n11002) );
  INVX1 U11518 ( .A(n7164), .Y(n9436) );
  NAND2X1 U11519 ( .A(n7164), .B(n11069), .Y(n11135) );
  NAND2X1 U11520 ( .A(n7164), .B(n6905), .Y(n11124) );
  ADDHXL U11521 ( .A(n11120), .B(n11119), .S(n7164) );
  NAND2X1 U11522 ( .A(n11141), .B(n11142), .Y(n11119) );
  NAND2X1 U11523 ( .A(n10014), .B(n11122), .Y(n11142) );
  ADDHXL U11524 ( .A(n11123), .B(n9085), .S(n11141) );
  NAND4X1 U11525 ( .A(n11143), .B(n11144), .C(n11145), .D(n11146), .Y(n11123)
         );
  NAND2X1 U11526 ( .A(G21587), .B(n10224), .Y(n11146) );
  NAND2X1 U11527 ( .A(G21778), .B(n9260), .Y(n11145) );
  NAND2X1 U11528 ( .A(n7165), .B(n10272), .Y(n11144) );
  INVX1 U11529 ( .A(n9847), .Y(n7165) );
  NAND2X1 U11530 ( .A(n11045), .B(n11147), .Y(n9847) );
  NAND2X1 U11531 ( .A(n11148), .B(n11149), .Y(n11147) );
  OR2X1 U11532 ( .A(n11149), .B(n11148), .Y(n11045) );
  ADDHXL U11533 ( .A(n11150), .B(n10227), .S(n11148) );
  NAND3X1 U11534 ( .A(n11151), .B(n11152), .C(n11153), .Y(n11150) );
  NOR3X1 U11535 ( .A(n11154), .B(n11155), .C(n11156), .Y(n11153) );
  AND2X1 U11536 ( .A(n10236), .B(G21714), .Y(n11156) );
  NOR2X1 U11537 ( .A(n9085), .B(n9434), .Y(n11155) );
  INVX1 U11538 ( .A(G21619), .Y(n9434) );
  NOR2X1 U11539 ( .A(n7162), .B(n9266), .Y(n11154) );
  AND2X1 U11540 ( .A(n11157), .B(n11158), .Y(n7162) );
  NAND2X1 U11541 ( .A(n10586), .B(n8711), .Y(n11158) );
  NAND4X1 U11542 ( .A(n11159), .B(n11160), .C(n11161), .D(n11162), .Y(n10586)
         );
  NOR4X1 U11543 ( .A(n11163), .B(n11164), .C(n11165), .D(n11166), .Y(n11162)
         );
  NOR2X1 U11544 ( .A(n10573), .B(n7597), .Y(n11166) );
  NOR2X1 U11545 ( .A(n10574), .B(n7677), .Y(n11165) );
  NOR2X1 U11546 ( .A(n10575), .B(n7757), .Y(n11164) );
  NOR2X1 U11547 ( .A(n10581), .B(n7919), .Y(n11163) );
  NOR4X1 U11548 ( .A(n11167), .B(n11168), .C(n11169), .D(n11170), .Y(n11161)
         );
  NOR2X1 U11549 ( .A(n10582), .B(n7997), .Y(n11170) );
  NOR2X1 U11550 ( .A(n10583), .B(n8075), .Y(n11169) );
  NOR2X1 U11551 ( .A(n10566), .B(n8234), .Y(n11168) );
  NOR2X1 U11552 ( .A(n10565), .B(n8312), .Y(n11167) );
  NOR4X1 U11553 ( .A(n11171), .B(n11172), .C(n11173), .D(n11174), .Y(n11160)
         );
  NOR2X1 U11554 ( .A(n10564), .B(n8390), .Y(n11174) );
  NOR2X1 U11555 ( .A(n10558), .B(n8551), .Y(n11173) );
  NOR2X1 U11556 ( .A(n10557), .B(n8629), .Y(n11172) );
  NOR2X1 U11557 ( .A(n10556), .B(n8706), .Y(n11171) );
  NOR4X1 U11558 ( .A(n11175), .B(n11176), .C(n11177), .D(n11178), .Y(n11159)
         );
  NOR2X1 U11559 ( .A(n10572), .B(n7487), .Y(n11178) );
  NOR2X1 U11560 ( .A(n10580), .B(n7839), .Y(n11177) );
  NOR2X1 U11561 ( .A(n10567), .B(n8154), .Y(n11176) );
  NOR2X1 U11562 ( .A(n10559), .B(n8469), .Y(n11175) );
  NAND2X1 U11563 ( .A(n11179), .B(n9076), .Y(n11157) );
  ADDHXL U11564 ( .A(G21587), .B(n11088), .S(n11179) );
  NOR2X1 U11565 ( .A(n11180), .B(n7175), .Y(n11088) );
  NAND2X1 U11566 ( .A(G21587), .B(n10503), .Y(n11152) );
  NAND2X1 U11567 ( .A(G21746), .B(n10333), .Y(n11151) );
  OR2X1 U11568 ( .A(n11181), .B(n11182), .Y(n11149) );
  NAND2X1 U11569 ( .A(G21619), .B(n10225), .Y(n11143) );
  NAND2X1 U11570 ( .A(n11183), .B(n11184), .Y(n11120) );
  NAND2X1 U11571 ( .A(n11185), .B(n11186), .Y(n11184) );
  NAND4X1 U11572 ( .A(n11187), .B(n11188), .C(n11189), .D(n11190), .Y(G1008)
         );
  NOR2X1 U11573 ( .A(n11191), .B(n11192), .Y(n11190) );
  NOR2X1 U11574 ( .A(n6891), .B(n9446), .Y(n11192) );
  NOR2X1 U11575 ( .A(n6901), .B(n7173), .Y(n11191) );
  NAND2X1 U11576 ( .A(n7178), .B(n6882), .Y(n11189) );
  NAND2X1 U11577 ( .A(n6903), .B(n7176), .Y(n11188) );
  ADDFXL U11578 ( .A(n9926), .B(n11134), .CI(n11133), .S(n7176) );
  NAND2X1 U11579 ( .A(n11193), .B(n11194), .Y(n11133) );
  NAND2X1 U11580 ( .A(n9926), .B(n11195), .Y(n11194) );
  OR2X1 U11581 ( .A(n11196), .B(n11197), .Y(n11195) );
  NAND2X1 U11582 ( .A(n11197), .B(n11196), .Y(n11193) );
  NAND4X1 U11583 ( .A(n11198), .B(n11199), .C(n11200), .D(n11201), .Y(n11134)
         );
  NOR2X1 U11584 ( .A(n11202), .B(n11203), .Y(n11201) );
  NOR2X1 U11585 ( .A(n10216), .B(n7175), .Y(n11203) );
  INVX1 U11586 ( .A(G21586), .Y(n7175) );
  NOR2X1 U11587 ( .A(n10226), .B(n7173), .Y(n11202) );
  INVX1 U11588 ( .A(G21777), .Y(n7173) );
  NAND2X1 U11589 ( .A(n7178), .B(n9926), .Y(n11200) );
  NAND4X1 U11590 ( .A(n7202), .B(n11204), .C(n7189), .D(n11004), .Y(n11199) );
  NAND2X1 U11591 ( .A(n7177), .B(n11069), .Y(n11198) );
  NAND2X1 U11592 ( .A(n10217), .B(n11205), .Y(n11069) );
  NAND4X1 U11593 ( .A(n7215), .B(n11206), .C(n7189), .D(n11207), .Y(n11004) );
  NOR2X1 U11594 ( .A(n9445), .B(n9465), .Y(n11207) );
  NAND2X1 U11595 ( .A(n7177), .B(n6905), .Y(n11187) );
  INVX1 U11596 ( .A(n9445), .Y(n7177) );
  ADDHXL U11597 ( .A(n11208), .B(n11186), .S(n9445) );
  NAND2X1 U11598 ( .A(n11209), .B(n11210), .Y(n11186) );
  NAND2X1 U11599 ( .A(n11211), .B(n11212), .Y(n11210) );
  NAND3X1 U11600 ( .A(n10014), .B(n11213), .C(n11214), .Y(n11209) );
  ADDHXL U11601 ( .A(n7564), .B(n11215), .S(n11214) );
  NAND2X1 U11602 ( .A(n11183), .B(n11185), .Y(n11208) );
  NAND2X1 U11603 ( .A(n11216), .B(n11217), .Y(n11185) );
  NAND2X1 U11604 ( .A(n10014), .B(n11218), .Y(n11217) );
  ADDHXL U11605 ( .A(n9085), .B(n11219), .S(n11216) );
  NAND3X1 U11606 ( .A(n10014), .B(n11218), .C(n11220), .Y(n11183) );
  ADDHXL U11607 ( .A(n11219), .B(n7564), .S(n11220) );
  NAND4X1 U11608 ( .A(n11221), .B(n11222), .C(n11223), .D(n11224), .Y(n11219)
         );
  NAND2X1 U11609 ( .A(n7178), .B(n10272), .Y(n11224) );
  ADDHXL U11610 ( .A(n11181), .B(n11182), .S(n7178) );
  ADDHXL U11611 ( .A(n11225), .B(n10227), .S(n11182) );
  NAND3X1 U11612 ( .A(n11226), .B(n11227), .C(n11228), .Y(n11225) );
  NOR3X1 U11613 ( .A(n11229), .B(n11230), .C(n11231), .Y(n11228) );
  AND2X1 U11614 ( .A(n10236), .B(G21713), .Y(n11231) );
  NOR2X1 U11615 ( .A(n9085), .B(n9446), .Y(n11230) );
  INVX1 U11616 ( .A(G21618), .Y(n9446) );
  NOR2X1 U11617 ( .A(n7174), .B(n9266), .Y(n11229) );
  AND3X1 U11618 ( .A(n11232), .B(n11233), .C(n11234), .Y(n7174) );
  OR2X1 U11619 ( .A(n11180), .B(G21586), .Y(n11234) );
  NAND3X1 U11620 ( .A(G21586), .B(n11180), .C(n9076), .Y(n11233) );
  NAND2X1 U11621 ( .A(n11235), .B(G21585), .Y(n11180) );
  NAND2X1 U11622 ( .A(n10673), .B(n8711), .Y(n11232) );
  NAND4X1 U11623 ( .A(n11236), .B(n11237), .C(n11238), .D(n11239), .Y(n10673)
         );
  NOR4X1 U11624 ( .A(n11240), .B(n11241), .C(n11242), .D(n11243), .Y(n11239)
         );
  NOR2X1 U11625 ( .A(n10655), .B(n7597), .Y(n11243) );
  NOR2X1 U11626 ( .A(n10656), .B(n7677), .Y(n11242) );
  NOR2X1 U11627 ( .A(n10657), .B(n7757), .Y(n11241) );
  NOR2X1 U11628 ( .A(n10663), .B(n7919), .Y(n11240) );
  NOR4X1 U11629 ( .A(n11244), .B(n11245), .C(n11246), .D(n11247), .Y(n11238)
         );
  NOR2X1 U11630 ( .A(n10664), .B(n7997), .Y(n11247) );
  NOR2X1 U11631 ( .A(n10665), .B(n8075), .Y(n11246) );
  NOR2X1 U11632 ( .A(n10648), .B(n8234), .Y(n11245) );
  NOR2X1 U11633 ( .A(n10647), .B(n8312), .Y(n11244) );
  NOR4X1 U11634 ( .A(n11248), .B(n11249), .C(n11250), .D(n11251), .Y(n11237)
         );
  NOR2X1 U11635 ( .A(n10646), .B(n8390), .Y(n11251) );
  NOR2X1 U11636 ( .A(n10640), .B(n8551), .Y(n11250) );
  NOR2X1 U11637 ( .A(n10639), .B(n8629), .Y(n11249) );
  NOR2X1 U11638 ( .A(n10638), .B(n8706), .Y(n11248) );
  NOR4X1 U11639 ( .A(n11252), .B(n11253), .C(n11254), .D(n11255), .Y(n11236)
         );
  NOR2X1 U11640 ( .A(n10654), .B(n7487), .Y(n11255) );
  NOR2X1 U11641 ( .A(n10662), .B(n7839), .Y(n11254) );
  NOR2X1 U11642 ( .A(n10649), .B(n8154), .Y(n11253) );
  NOR2X1 U11643 ( .A(n10641), .B(n8469), .Y(n11252) );
  NAND2X1 U11644 ( .A(G21586), .B(n10503), .Y(n11227) );
  NAND2X1 U11645 ( .A(G21745), .B(n10333), .Y(n11226) );
  NAND2X1 U11646 ( .A(G21586), .B(n10224), .Y(n11223) );
  NAND2X1 U11647 ( .A(G21618), .B(n10225), .Y(n11222) );
  NAND2X1 U11648 ( .A(G21777), .B(n9260), .Y(n11221) );
  NAND4X1 U11649 ( .A(n11256), .B(n11257), .C(n11258), .D(n11259), .Y(G1007)
         );
  NOR2X1 U11650 ( .A(n11260), .B(n11261), .Y(n11259) );
  NOR2X1 U11651 ( .A(n6891), .B(n9456), .Y(n11261) );
  NOR2X1 U11652 ( .A(n6901), .B(n7186), .Y(n11260) );
  NAND2X1 U11653 ( .A(n7190), .B(n6882), .Y(n11258) );
  NAND2X1 U11654 ( .A(n6903), .B(n7188), .Y(n11257) );
  ADDFXL U11655 ( .A(n9926), .B(n11197), .CI(n11196), .S(n7188) );
  NAND2X1 U11656 ( .A(n11262), .B(n11263), .Y(n11196) );
  NAND2X1 U11657 ( .A(n9926), .B(n11264), .Y(n11263) );
  OR2X1 U11658 ( .A(n11265), .B(n11266), .Y(n11264) );
  NAND2X1 U11659 ( .A(n11266), .B(n11265), .Y(n11262) );
  NAND4X1 U11660 ( .A(n11267), .B(n11268), .C(n11269), .D(n11270), .Y(n11197)
         );
  NOR2X1 U11661 ( .A(n11271), .B(n11272), .Y(n11270) );
  NOR2X1 U11662 ( .A(n10226), .B(n7186), .Y(n11272) );
  INVX1 U11663 ( .A(G21776), .Y(n7186) );
  NOR2X1 U11664 ( .A(n9908), .B(n9862), .Y(n11271) );
  NAND2X1 U11665 ( .A(G21585), .B(n10444), .Y(n11269) );
  NAND2X1 U11666 ( .A(n7189), .B(n11273), .Y(n11268) );
  NAND2X1 U11667 ( .A(n11274), .B(n11275), .Y(n11273) );
  NAND2X1 U11668 ( .A(n10256), .B(n9465), .Y(n11275) );
  NAND3X1 U11669 ( .A(n11204), .B(n7202), .C(n9455), .Y(n11267) );
  INVX1 U11670 ( .A(n7189), .Y(n9455) );
  NAND2X1 U11671 ( .A(n7189), .B(n6905), .Y(n11256) );
  ADDHXL U11672 ( .A(n11211), .B(n11212), .S(n7189) );
  NAND2X1 U11673 ( .A(n11276), .B(n11277), .Y(n11212) );
  NAND2X1 U11674 ( .A(n11278), .B(n11279), .Y(n11277) );
  NAND2X1 U11675 ( .A(n11280), .B(n11281), .Y(n11211) );
  NAND2X1 U11676 ( .A(n10014), .B(n11213), .Y(n11281) );
  ADDHXL U11677 ( .A(n11215), .B(n9085), .S(n11280) );
  NAND4X1 U11678 ( .A(n11282), .B(n11283), .C(n11284), .D(n11285), .Y(n11215)
         );
  NAND2X1 U11679 ( .A(G21585), .B(n10224), .Y(n11285) );
  NAND2X1 U11680 ( .A(G21776), .B(n9260), .Y(n11284) );
  NAND2X1 U11681 ( .A(n7190), .B(n10272), .Y(n11283) );
  INVX1 U11682 ( .A(n9862), .Y(n7190) );
  NAND2X1 U11683 ( .A(n11181), .B(n11286), .Y(n9862) );
  NAND2X1 U11684 ( .A(n11287), .B(n11288), .Y(n11286) );
  OR2X1 U11685 ( .A(n11288), .B(n11287), .Y(n11181) );
  ADDHXL U11686 ( .A(n11289), .B(n10227), .S(n11287) );
  NAND3X1 U11687 ( .A(n11290), .B(n11291), .C(n11292), .Y(n11289) );
  NOR3X1 U11688 ( .A(n11293), .B(n11294), .C(n11295), .Y(n11292) );
  AND2X1 U11689 ( .A(n10236), .B(G21712), .Y(n11295) );
  NOR2X1 U11690 ( .A(n9085), .B(n9456), .Y(n11294) );
  INVX1 U11691 ( .A(G21617), .Y(n9456) );
  NOR2X1 U11692 ( .A(n7187), .B(n9266), .Y(n11293) );
  AND2X1 U11693 ( .A(n11296), .B(n11297), .Y(n7187) );
  NAND2X1 U11694 ( .A(n10757), .B(n8711), .Y(n11297) );
  NAND4X1 U11695 ( .A(n11298), .B(n11299), .C(n11300), .D(n11301), .Y(n10757)
         );
  NOR4X1 U11696 ( .A(n11302), .B(n11303), .C(n11304), .D(n11305), .Y(n11301)
         );
  NOR2X1 U11697 ( .A(n10744), .B(n7597), .Y(n11305) );
  NOR2X1 U11698 ( .A(n10745), .B(n7677), .Y(n11304) );
  NOR2X1 U11699 ( .A(n10746), .B(n7757), .Y(n11303) );
  NOR2X1 U11700 ( .A(n10752), .B(n7919), .Y(n11302) );
  NOR4X1 U11701 ( .A(n11306), .B(n11307), .C(n11308), .D(n11309), .Y(n11300)
         );
  NOR2X1 U11702 ( .A(n10753), .B(n7997), .Y(n11309) );
  NOR2X1 U11703 ( .A(n10754), .B(n8075), .Y(n11308) );
  NOR2X1 U11704 ( .A(n10737), .B(n8234), .Y(n11307) );
  NOR2X1 U11705 ( .A(n10736), .B(n8312), .Y(n11306) );
  NOR4X1 U11706 ( .A(n11310), .B(n11311), .C(n11312), .D(n11313), .Y(n11299)
         );
  NOR2X1 U11707 ( .A(n10735), .B(n8390), .Y(n11313) );
  NOR2X1 U11708 ( .A(n10729), .B(n8551), .Y(n11312) );
  NOR2X1 U11709 ( .A(n10728), .B(n8629), .Y(n11311) );
  NOR2X1 U11710 ( .A(n10727), .B(n8706), .Y(n11310) );
  NOR4X1 U11711 ( .A(n11314), .B(n11315), .C(n11316), .D(n11317), .Y(n11298)
         );
  NOR2X1 U11712 ( .A(n10743), .B(n7487), .Y(n11317) );
  NOR2X1 U11713 ( .A(n10751), .B(n7839), .Y(n11316) );
  NOR2X1 U11714 ( .A(n10738), .B(n8154), .Y(n11315) );
  NOR2X1 U11715 ( .A(n10730), .B(n8469), .Y(n11314) );
  NAND2X1 U11716 ( .A(n11318), .B(n9076), .Y(n11296) );
  ADDHXL U11717 ( .A(G21585), .B(n11235), .S(n11318) );
  NOR2X1 U11718 ( .A(n11319), .B(n7200), .Y(n11235) );
  INVX1 U11719 ( .A(G21584), .Y(n7200) );
  NAND2X1 U11720 ( .A(G21585), .B(n10503), .Y(n11291) );
  NAND2X1 U11721 ( .A(G21744), .B(n10333), .Y(n11290) );
  OR2X1 U11722 ( .A(n11320), .B(n11321), .Y(n11288) );
  NAND2X1 U11723 ( .A(G21617), .B(n10225), .Y(n11282) );
  NAND4X1 U11724 ( .A(n11322), .B(n11323), .C(n11324), .D(n11325), .Y(G1006)
         );
  NOR2X1 U11725 ( .A(n11326), .B(n11327), .Y(n11325) );
  NOR2X1 U11726 ( .A(n6891), .B(n9466), .Y(n11327) );
  NAND2X1 U11727 ( .A(n7203), .B(n6882), .Y(n11324) );
  NAND2X1 U11728 ( .A(n6903), .B(n7201), .Y(n11323) );
  ADDFXL U11729 ( .A(n9926), .B(n11266), .CI(n11265), .S(n7201) );
  NAND2X1 U11730 ( .A(n11328), .B(n11329), .Y(n11265) );
  NAND2X1 U11731 ( .A(n9926), .B(n11330), .Y(n11329) );
  OR2X1 U11732 ( .A(n11331), .B(n11332), .Y(n11330) );
  NAND2X1 U11733 ( .A(n11332), .B(n11331), .Y(n11328) );
  NAND4X1 U11734 ( .A(n11333), .B(n11334), .C(n11335), .D(n11336), .Y(n11266)
         );
  NOR2X1 U11735 ( .A(n11337), .B(n11338), .Y(n11336) );
  NOR2X1 U11736 ( .A(n10226), .B(n7198), .Y(n11338) );
  INVX1 U11737 ( .A(G21775), .Y(n7198) );
  NOR2X1 U11738 ( .A(n9908), .B(n9870), .Y(n11337) );
  INVX1 U11739 ( .A(n7203), .Y(n9870) );
  NAND2X1 U11740 ( .A(G21584), .B(n10444), .Y(n11335) );
  NAND2X1 U11741 ( .A(n11204), .B(n9465), .Y(n11334) );
  NOR3X1 U11742 ( .A(n9475), .B(n11339), .C(n9192), .Y(n11204) );
  OR2X1 U11743 ( .A(n9465), .B(n11274), .Y(n11333) );
  NOR2X1 U11744 ( .A(n11340), .B(n11341), .Y(n11274) );
  NOR2X1 U11745 ( .A(n7215), .B(n9192), .Y(n11341) );
  NAND2X1 U11746 ( .A(n7202), .B(n6905), .Y(n11322) );
  INVX1 U11747 ( .A(n9465), .Y(n7202) );
  ADDHXL U11748 ( .A(n11342), .B(n11279), .S(n9465) );
  NAND2X1 U11749 ( .A(n11343), .B(n11344), .Y(n11279) );
  NAND2X1 U11750 ( .A(n11345), .B(n11346), .Y(n11344) );
  INVX1 U11751 ( .A(n11347), .Y(n11345) );
  NAND2X1 U11752 ( .A(n11276), .B(n11278), .Y(n11342) );
  NAND2X1 U11753 ( .A(n11348), .B(n11349), .Y(n11278) );
  NAND2X1 U11754 ( .A(n10014), .B(n11350), .Y(n11349) );
  ADDHXL U11755 ( .A(n9085), .B(n11351), .S(n11348) );
  NAND3X1 U11756 ( .A(n10014), .B(n11350), .C(n11352), .Y(n11276) );
  ADDHXL U11757 ( .A(n11351), .B(n7564), .S(n11352) );
  NAND4X1 U11758 ( .A(n11353), .B(n11354), .C(n11355), .D(n11356), .Y(n11351)
         );
  NAND2X1 U11759 ( .A(n7203), .B(n10272), .Y(n11356) );
  ADDHXL U11760 ( .A(n11320), .B(n11321), .S(n7203) );
  ADDHXL U11761 ( .A(n11357), .B(n10227), .S(n11321) );
  NAND3X1 U11762 ( .A(n11358), .B(n11359), .C(n11360), .Y(n11357) );
  NOR3X1 U11763 ( .A(n11361), .B(n11362), .C(n11363), .Y(n11360) );
  AND2X1 U11764 ( .A(n10236), .B(G21711), .Y(n11363) );
  NOR2X1 U11765 ( .A(n9085), .B(n9466), .Y(n11362) );
  INVX1 U11766 ( .A(G21616), .Y(n9466) );
  NOR2X1 U11767 ( .A(n7199), .B(n9266), .Y(n11361) );
  AND3X1 U11768 ( .A(n11364), .B(n11365), .C(n11366), .Y(n7199) );
  OR2X1 U11769 ( .A(n11319), .B(G21584), .Y(n11366) );
  NAND3X1 U11770 ( .A(G21584), .B(n11319), .C(n9076), .Y(n11365) );
  NAND2X1 U11771 ( .A(n11367), .B(G21583), .Y(n11319) );
  NAND2X1 U11772 ( .A(n10795), .B(n8711), .Y(n11364) );
  NAND4X1 U11773 ( .A(n11368), .B(n11369), .C(n11370), .D(n11371), .Y(n10795)
         );
  NOR4X1 U11774 ( .A(n11372), .B(n11373), .C(n11374), .D(n11375), .Y(n11371)
         );
  NOR2X1 U11775 ( .A(n10834), .B(n7597), .Y(n11375) );
  NOR2X1 U11776 ( .A(n10835), .B(n7677), .Y(n11374) );
  NOR2X1 U11777 ( .A(n10836), .B(n7757), .Y(n11373) );
  NOR2X1 U11778 ( .A(n10842), .B(n7919), .Y(n11372) );
  NOR4X1 U11779 ( .A(n11376), .B(n11377), .C(n11378), .D(n11379), .Y(n11370)
         );
  NOR2X1 U11780 ( .A(n10843), .B(n7997), .Y(n11379) );
  NOR2X1 U11781 ( .A(n10844), .B(n8075), .Y(n11378) );
  NOR2X1 U11782 ( .A(n10827), .B(n8234), .Y(n11377) );
  NOR2X1 U11783 ( .A(n10826), .B(n8312), .Y(n11376) );
  NOR4X1 U11784 ( .A(n11380), .B(n11381), .C(n11382), .D(n11383), .Y(n11369)
         );
  NOR2X1 U11785 ( .A(n10825), .B(n8390), .Y(n11383) );
  NOR2X1 U11786 ( .A(n10819), .B(n8551), .Y(n11382) );
  NOR2X1 U11787 ( .A(n10818), .B(n8629), .Y(n11381) );
  NOR2X1 U11788 ( .A(n10817), .B(n8706), .Y(n11380) );
  NOR4X1 U11789 ( .A(n11384), .B(n11385), .C(n11386), .D(n11387), .Y(n11368)
         );
  NOR2X1 U11790 ( .A(n10833), .B(n7487), .Y(n11387) );
  NOR2X1 U11791 ( .A(n10841), .B(n7839), .Y(n11386) );
  NOR2X1 U11792 ( .A(n10828), .B(n8154), .Y(n11385) );
  NOR2X1 U11793 ( .A(n10820), .B(n8469), .Y(n11384) );
  NAND2X1 U11794 ( .A(G21584), .B(n10503), .Y(n11359) );
  NAND2X1 U11795 ( .A(G21743), .B(n10333), .Y(n11358) );
  NAND2X1 U11796 ( .A(G21584), .B(n10224), .Y(n11355) );
  NAND2X1 U11797 ( .A(G21616), .B(n10225), .Y(n11354) );
  NAND2X1 U11798 ( .A(G21775), .B(n9260), .Y(n11353) );
  NAND4X1 U11799 ( .A(n11388), .B(n11389), .C(n11390), .D(n11391), .Y(G1005)
         );
  NOR2X1 U11800 ( .A(n11392), .B(n11393), .Y(n11391) );
  NOR2X1 U11801 ( .A(n6891), .B(n9476), .Y(n11393) );
  NOR2X1 U11802 ( .A(n6901), .B(n7211), .Y(n11392) );
  NAND2X1 U11803 ( .A(n7216), .B(n6882), .Y(n11390) );
  NAND2X1 U11804 ( .A(n6903), .B(n7214), .Y(n11389) );
  ADDFXL U11805 ( .A(n9926), .B(n11332), .CI(n11331), .S(n7214) );
  NAND2X1 U11806 ( .A(n11394), .B(n11395), .Y(n11331) );
  NAND2X1 U11807 ( .A(n9926), .B(n11396), .Y(n11395) );
  OR2X1 U11808 ( .A(n11397), .B(n11398), .Y(n11396) );
  NAND2X1 U11809 ( .A(n11398), .B(n11397), .Y(n11394) );
  NAND4X1 U11810 ( .A(n11399), .B(n11400), .C(n11401), .D(n11402), .Y(n11332)
         );
  NOR2X1 U11811 ( .A(n11403), .B(n11404), .Y(n11402) );
  NOR2X1 U11812 ( .A(n10226), .B(n7211), .Y(n11404) );
  INVX1 U11813 ( .A(G21774), .Y(n7211) );
  NOR2X1 U11814 ( .A(n9908), .B(n9878), .Y(n11403) );
  NAND2X1 U11815 ( .A(G21583), .B(n10444), .Y(n11401) );
  NAND2X1 U11816 ( .A(n7215), .B(n11340), .Y(n11400) );
  NAND2X1 U11817 ( .A(n10217), .B(n11405), .Y(n11340) );
  INVX1 U11818 ( .A(n11206), .Y(n11339) );
  NAND3X1 U11819 ( .A(n10256), .B(n11206), .C(n9475), .Y(n11399) );
  INVX1 U11820 ( .A(n7215), .Y(n9475) );
  NAND2X1 U11821 ( .A(n11406), .B(n11407), .Y(n11206) );
  NAND2X1 U11822 ( .A(n11408), .B(n11409), .Y(n11407) );
  NAND2X1 U11823 ( .A(n9485), .B(n11410), .Y(n11408) );
  OR2X1 U11824 ( .A(n9485), .B(n11410), .Y(n11406) );
  NAND2X1 U11825 ( .A(n6905), .B(n7215), .Y(n11388) );
  ADDHXL U11826 ( .A(n11411), .B(n11347), .S(n7215) );
  NAND2X1 U11827 ( .A(n11343), .B(n11346), .Y(n11411) );
  NAND2X1 U11828 ( .A(n11412), .B(n11413), .Y(n11346) );
  NAND2X1 U11829 ( .A(n10014), .B(n11414), .Y(n11413) );
  ADDHXL U11830 ( .A(n11415), .B(n7564), .S(n11412) );
  NAND3X1 U11831 ( .A(n10014), .B(n11414), .C(n11416), .Y(n11343) );
  ADDHXL U11832 ( .A(n9085), .B(n11415), .S(n11416) );
  AND4X1 U11833 ( .A(n11417), .B(n11418), .C(n11419), .D(n11420), .Y(n11415)
         );
  NAND2X1 U11834 ( .A(G21583), .B(n10224), .Y(n11420) );
  NAND2X1 U11835 ( .A(G21774), .B(n9260), .Y(n11419) );
  NAND2X1 U11836 ( .A(n7216), .B(n10272), .Y(n11418) );
  INVX1 U11837 ( .A(n9878), .Y(n7216) );
  NAND2X1 U11838 ( .A(n11320), .B(n11421), .Y(n9878) );
  NAND3X1 U11839 ( .A(n11422), .B(n11423), .C(n11424), .Y(n11421) );
  ADDHXL U11840 ( .A(n11425), .B(n10227), .S(n11424) );
  NAND2X1 U11841 ( .A(n11426), .B(n11427), .Y(n11320) );
  NAND2X1 U11842 ( .A(n11422), .B(n11423), .Y(n11427) );
  NAND2X1 U11843 ( .A(n11428), .B(n11429), .Y(n11422) );
  ADDHXL U11844 ( .A(n11425), .B(n9260), .S(n11426) );
  NAND3X1 U11845 ( .A(n11430), .B(n11431), .C(n11432), .Y(n11425) );
  NOR3X1 U11846 ( .A(n11433), .B(n11434), .C(n11435), .Y(n11432) );
  AND2X1 U11847 ( .A(n10236), .B(G21710), .Y(n11435) );
  NOR2X1 U11848 ( .A(n9085), .B(n9476), .Y(n11434) );
  INVX1 U11849 ( .A(G21615), .Y(n9476) );
  NOR2X1 U11850 ( .A(n7212), .B(n9266), .Y(n11433) );
  INVX1 U11851 ( .A(n9755), .Y(n9266) );
  AND2X1 U11852 ( .A(n11436), .B(n11437), .Y(n7212) );
  NAND2X1 U11853 ( .A(n11367), .B(n7213), .Y(n11437) );
  INVX1 U11854 ( .A(G21583), .Y(n7213) );
  NAND2X1 U11855 ( .A(n11438), .B(n11439), .Y(n11436) );
  INVX1 U11856 ( .A(n11367), .Y(n11439) );
  NOR3X1 U11857 ( .A(n7224), .B(n7227), .C(n7225), .Y(n11367) );
  OR3X1 U11858 ( .A(n7257), .B(n7254), .C(n7255), .Y(n7225) );
  NAND3X1 U11859 ( .A(G21578), .B(G21577), .C(n7302), .Y(n7255) );
  NOR2X1 U11860 ( .A(n7312), .B(n7313), .Y(n7302) );
  NAND2X1 U11861 ( .A(n7323), .B(G21575), .Y(n7313) );
  NOR3X1 U11862 ( .A(n7336), .B(n7333), .C(n7334), .Y(n7323) );
  NAND3X1 U11863 ( .A(G21572), .B(G21571), .C(n7377), .Y(n7334) );
  NOR2X1 U11864 ( .A(n7375), .B(n7378), .Y(n7377) );
  AND2X1 U11865 ( .A(n7391), .B(n7390), .Y(n7378) );
  NAND2X1 U11866 ( .A(G21569), .B(n9076), .Y(n7390) );
  NAND2X1 U11867 ( .A(n7401), .B(G21568), .Y(n7391) );
  NOR2X1 U11868 ( .A(n8711), .B(n11440), .Y(n7401) );
  INVX1 U11869 ( .A(G21573), .Y(n7333) );
  INVX1 U11870 ( .A(G21574), .Y(n7336) );
  NAND2X1 U11871 ( .A(G21576), .B(n9076), .Y(n7312) );
  NAND2X1 U11872 ( .A(n11441), .B(n11442), .Y(n11438) );
  NAND2X1 U11873 ( .A(G21583), .B(n9076), .Y(n11442) );
  NAND2X1 U11874 ( .A(n10984), .B(n8711), .Y(n11441) );
  NAND4X1 U11875 ( .A(n11443), .B(n11444), .C(n11445), .D(n11446), .Y(n10984)
         );
  NOR4X1 U11876 ( .A(n11447), .B(n11448), .C(n11449), .D(n11450), .Y(n11446)
         );
  NOR2X1 U11877 ( .A(n10929), .B(n7597), .Y(n11450) );
  NAND2X1 U11878 ( .A(n11451), .B(n11452), .Y(n7597) );
  NOR2X1 U11879 ( .A(n10931), .B(n7677), .Y(n11449) );
  NAND2X1 U11880 ( .A(n11453), .B(n11454), .Y(n7677) );
  NOR2X1 U11881 ( .A(n10932), .B(n7757), .Y(n11448) );
  NAND2X1 U11882 ( .A(n11451), .B(n11454), .Y(n7757) );
  NOR2X1 U11883 ( .A(n10940), .B(n7919), .Y(n11447) );
  NAND2X1 U11884 ( .A(n11452), .B(n11455), .Y(n7919) );
  NOR4X1 U11885 ( .A(n11456), .B(n11457), .C(n11458), .D(n11459), .Y(n11445)
         );
  NOR2X1 U11886 ( .A(n10941), .B(n7997), .Y(n11459) );
  NAND2X1 U11887 ( .A(n11460), .B(n11454), .Y(n7997) );
  NOR2X1 U11888 ( .A(n10942), .B(n8075), .Y(n11458) );
  NAND2X1 U11889 ( .A(n11454), .B(n11455), .Y(n8075) );
  NOR2X1 U11890 ( .A(n11461), .B(n9132), .Y(n11454) );
  NOR2X1 U11891 ( .A(n10919), .B(n8234), .Y(n11457) );
  NAND2X1 U11892 ( .A(n11462), .B(n11451), .Y(n8234) );
  NOR2X1 U11893 ( .A(n10918), .B(n8312), .Y(n11456) );
  NAND2X1 U11894 ( .A(n11463), .B(n11453), .Y(n8312) );
  NOR4X1 U11895 ( .A(n11464), .B(n11465), .C(n11466), .D(n11467), .Y(n11444)
         );
  NOR2X1 U11896 ( .A(n10916), .B(n8390), .Y(n11467) );
  NAND2X1 U11897 ( .A(n11463), .B(n11451), .Y(n8390) );
  NOR2X1 U11898 ( .A(n11468), .B(n9110), .Y(n11451) );
  NOR2X1 U11899 ( .A(n10909), .B(n8551), .Y(n11466) );
  NAND2X1 U11900 ( .A(n11462), .B(n11455), .Y(n8551) );
  NOR2X1 U11901 ( .A(n10907), .B(n8629), .Y(n11465) );
  NAND2X1 U11902 ( .A(n11460), .B(n11463), .Y(n8629) );
  NOR2X1 U11903 ( .A(n10904), .B(n8706), .Y(n11464) );
  NAND2X1 U11904 ( .A(n11463), .B(n11455), .Y(n8706) );
  NOR2X1 U11905 ( .A(n9110), .B(n9155), .Y(n11455) );
  NOR2X1 U11906 ( .A(n9132), .B(n9173), .Y(n11463) );
  NOR4X1 U11907 ( .A(n11469), .B(n11470), .C(n11471), .D(n11472), .Y(n11443)
         );
  NOR2X1 U11908 ( .A(n10927), .B(n7487), .Y(n11472) );
  NAND2X1 U11909 ( .A(n11453), .B(n11452), .Y(n7487) );
  NOR2X1 U11910 ( .A(n10939), .B(n7839), .Y(n11471) );
  NAND2X1 U11911 ( .A(n11460), .B(n11452), .Y(n7839) );
  NOR2X1 U11912 ( .A(n11461), .B(n11473), .Y(n11452) );
  INVX1 U11913 ( .A(n9173), .Y(n11461) );
  NOR2X1 U11914 ( .A(n10922), .B(n8154), .Y(n11470) );
  NAND2X1 U11915 ( .A(n11462), .B(n11453), .Y(n8154) );
  NOR2X1 U11916 ( .A(n11468), .B(n11474), .Y(n11453) );
  INVX1 U11917 ( .A(n9155), .Y(n11468) );
  NOR2X1 U11918 ( .A(n10911), .B(n8469), .Y(n11469) );
  NAND2X1 U11919 ( .A(n11460), .B(n11462), .Y(n8469) );
  NOR2X1 U11920 ( .A(n9173), .B(n11473), .Y(n11462) );
  INVX1 U11921 ( .A(n9132), .Y(n11473) );
  NOR2X1 U11922 ( .A(n9155), .B(n11474), .Y(n11460) );
  INVX1 U11923 ( .A(n9110), .Y(n11474) );
  NAND2X1 U11924 ( .A(G21583), .B(n10503), .Y(n11431) );
  NAND2X1 U11925 ( .A(G21742), .B(n10333), .Y(n11430) );
  NAND2X1 U11926 ( .A(G21615), .B(n10225), .Y(n11417) );
  NAND4X1 U11927 ( .A(n11475), .B(n11476), .C(n11477), .D(n11478), .Y(G1004)
         );
  NOR2X1 U11928 ( .A(n11479), .B(n11480), .Y(n11478) );
  NOR2X1 U11929 ( .A(n6891), .B(n9486), .Y(n11480) );
  INVX1 U11930 ( .A(G21614), .Y(n9486) );
  NOR2X1 U11931 ( .A(n6901), .B(n7230), .Y(n11479) );
  NAND2X1 U11932 ( .A(n7233), .B(n6882), .Y(n11477) );
  NAND2X1 U11933 ( .A(n6903), .B(n7231), .Y(n11476) );
  ADDFXL U11934 ( .A(n9926), .B(n11398), .CI(n11397), .S(n7231) );
  NAND2X1 U11935 ( .A(n11481), .B(n11482), .Y(n11397) );
  NAND2X1 U11936 ( .A(n9926), .B(n11483), .Y(n11482) );
  OR2X1 U11937 ( .A(n11484), .B(n11485), .Y(n11483) );
  NAND2X1 U11938 ( .A(n11485), .B(n11484), .Y(n11481) );
  NAND4X1 U11939 ( .A(n11486), .B(n11487), .C(n11488), .D(n11489), .Y(n11398)
         );
  NOR2X1 U11940 ( .A(n11490), .B(n11491), .Y(n11489) );
  NOR2X1 U11941 ( .A(n10216), .B(n7227), .Y(n11491) );
  INVX1 U11942 ( .A(G21582), .Y(n7227) );
  NOR2X1 U11943 ( .A(n10226), .B(n7230), .Y(n11490) );
  INVX1 U11944 ( .A(G21773), .Y(n7230) );
  NAND2X1 U11945 ( .A(n7233), .B(n9926), .Y(n11488) );
  ADDFXL U11946 ( .A(n11409), .B(n9485), .CI(n11410), .S(n11492) );
  NAND2X1 U11947 ( .A(n11493), .B(n11494), .Y(n11410) );
  NAND2X1 U11948 ( .A(n11495), .B(n11496), .Y(n11494) );
  OR2X1 U11949 ( .A(n9495), .B(n11497), .Y(n11496) );
  INVX1 U11950 ( .A(n11498), .Y(n11495) );
  NAND2X1 U11951 ( .A(n11497), .B(n9495), .Y(n11493) );
  NAND2X1 U11952 ( .A(n7232), .B(n11499), .Y(n11486) );
  NAND2X1 U11953 ( .A(n7232), .B(n6905), .Y(n11475) );
  INVX1 U11954 ( .A(n9485), .Y(n7232) );
  NAND2X1 U11955 ( .A(n11347), .B(n11500), .Y(n9485) );
  NAND2X1 U11956 ( .A(n11501), .B(n11502), .Y(n11500) );
  ADDHXL U11957 ( .A(n9085), .B(n11503), .S(n11501) );
  NAND2X1 U11958 ( .A(n11504), .B(n11505), .Y(n11347) );
  ADDHXL U11959 ( .A(n11503), .B(n7564), .S(n11504) );
  NAND4X1 U11960 ( .A(n11506), .B(n11507), .C(n11508), .D(n11509), .Y(n11503)
         );
  NAND2X1 U11961 ( .A(n7233), .B(n10272), .Y(n11509) );
  ADDHXL U11962 ( .A(n11429), .B(n11510), .S(n7233) );
  AND2X1 U11963 ( .A(n11428), .B(n11423), .Y(n11510) );
  NAND3X1 U11964 ( .A(n11511), .B(n11409), .C(n9755), .Y(n11423) );
  NAND2X1 U11965 ( .A(n11512), .B(n11513), .Y(n11428) );
  NAND2X1 U11966 ( .A(n9755), .B(n11409), .Y(n11513) );
  NAND4X1 U11967 ( .A(n11514), .B(n11515), .C(n11516), .D(n11517), .Y(n11409)
         );
  NOR4X1 U11968 ( .A(n11518), .B(n11519), .C(n11520), .D(n11521), .Y(n11517)
         );
  NOR2X1 U11969 ( .A(n10312), .B(n11522), .Y(n11521) );
  NOR2X1 U11970 ( .A(n10314), .B(n11523), .Y(n11520) );
  NOR2X1 U11971 ( .A(n10316), .B(n11524), .Y(n11519) );
  NOR2X1 U11972 ( .A(n10324), .B(n11525), .Y(n11518) );
  NOR4X1 U11973 ( .A(n11526), .B(n11527), .C(n11528), .D(n11529), .Y(n11516)
         );
  NOR2X1 U11974 ( .A(n10326), .B(n11530), .Y(n11529) );
  NOR2X1 U11975 ( .A(n10328), .B(n11531), .Y(n11528) );
  NOR2X1 U11976 ( .A(n10964), .B(n11532), .Y(n11527) );
  NOR2X1 U11977 ( .A(n10965), .B(n11533), .Y(n11526) );
  NOR4X1 U11978 ( .A(n11534), .B(n11535), .C(n11536), .D(n11537), .Y(n11515)
         );
  NOR2X1 U11979 ( .A(n10966), .B(n11538), .Y(n11537) );
  NOR2X1 U11980 ( .A(n10967), .B(n11539), .Y(n11536) );
  NOR2X1 U11981 ( .A(n10972), .B(n11540), .Y(n11535) );
  NOR2X1 U11982 ( .A(n10973), .B(n11541), .Y(n11534) );
  NOR4X1 U11983 ( .A(n11542), .B(n11543), .C(n11544), .D(n11545), .Y(n11514)
         );
  NOR2X1 U11984 ( .A(n10310), .B(n11546), .Y(n11545) );
  NOR2X1 U11985 ( .A(n10322), .B(n11547), .Y(n11544) );
  NOR2X1 U11986 ( .A(n10982), .B(n11548), .Y(n11543) );
  NOR2X1 U11987 ( .A(n10983), .B(n11549), .Y(n11542) );
  ADDHXL U11988 ( .A(n10227), .B(n11511), .S(n11512) );
  NAND4X1 U11989 ( .A(n11550), .B(n11551), .C(n11552), .D(n11553), .Y(n11511)
         );
  NAND2X1 U11990 ( .A(G21614), .B(n7564), .Y(n11553) );
  NAND2X1 U11991 ( .A(G21709), .B(n10236), .Y(n11552) );
  NAND2X1 U11992 ( .A(G21741), .B(n10333), .Y(n11551) );
  NAND2X1 U11993 ( .A(G21582), .B(n10503), .Y(n11550) );
  NAND2X1 U11994 ( .A(n11554), .B(n11555), .Y(n11429) );
  NAND2X1 U11995 ( .A(n11556), .B(n11557), .Y(n11555) );
  NAND2X1 U11996 ( .A(G21582), .B(n10224), .Y(n11508) );
  NAND2X1 U11997 ( .A(G21614), .B(n10225), .Y(n11507) );
  NAND2X1 U11998 ( .A(G21773), .B(n9260), .Y(n11506) );
  NAND4X1 U11999 ( .A(n11558), .B(n11559), .C(n11560), .D(n11561), .Y(G1003)
         );
  NOR2X1 U12000 ( .A(n11562), .B(n11563), .Y(n11561) );
  NOR2X1 U12001 ( .A(n6891), .B(n9496), .Y(n11563) );
  INVX1 U12002 ( .A(G21613), .Y(n9496) );
  NOR2X1 U12003 ( .A(n6901), .B(n7243), .Y(n11562) );
  NAND2X1 U12004 ( .A(n7246), .B(n6882), .Y(n11560) );
  NAND2X1 U12005 ( .A(n6903), .B(n7244), .Y(n11559) );
  ADDFXL U12006 ( .A(n9926), .B(n11484), .CI(n11485), .S(n7244) );
  NAND2X1 U12007 ( .A(n11564), .B(n11565), .Y(n11485) );
  NAND2X1 U12008 ( .A(n9926), .B(n11566), .Y(n11565) );
  OR2X1 U12009 ( .A(n11567), .B(n11568), .Y(n11566) );
  NAND2X1 U12010 ( .A(n11568), .B(n11567), .Y(n11564) );
  NAND4X1 U12011 ( .A(n11569), .B(n11570), .C(n11571), .D(n11572), .Y(n11484)
         );
  NOR2X1 U12012 ( .A(n11573), .B(n11574), .Y(n11572) );
  NOR2X1 U12013 ( .A(n10216), .B(n7224), .Y(n11574) );
  INVX1 U12014 ( .A(G21581), .Y(n7224) );
  NOR2X1 U12015 ( .A(n10226), .B(n7243), .Y(n11573) );
  INVX1 U12016 ( .A(G21772), .Y(n7243) );
  NAND2X1 U12017 ( .A(n7246), .B(n9926), .Y(n11571) );
  ADDFXL U12018 ( .A(n11498), .B(n9495), .CI(n11497), .S(n11575) );
  NAND2X1 U12019 ( .A(n11576), .B(n11577), .Y(n11497) );
  NAND2X1 U12020 ( .A(n11578), .B(n11579), .Y(n11577) );
  OR2X1 U12021 ( .A(n11580), .B(n9505), .Y(n11579) );
  NAND2X1 U12022 ( .A(n9505), .B(n11580), .Y(n11576) );
  NAND2X1 U12023 ( .A(n7245), .B(n11499), .Y(n11569) );
  NAND2X1 U12024 ( .A(n7245), .B(n6905), .Y(n11558) );
  INVX1 U12025 ( .A(n9495), .Y(n7245) );
  NAND2X1 U12026 ( .A(n11502), .B(n11581), .Y(n9495) );
  NAND2X1 U12027 ( .A(n11582), .B(n11583), .Y(n11581) );
  INVX1 U12028 ( .A(n11505), .Y(n11502) );
  NOR2X1 U12029 ( .A(n11583), .B(n11582), .Y(n11505) );
  ADDHXL U12030 ( .A(n11584), .B(n9085), .S(n11582) );
  NAND4X1 U12031 ( .A(n11585), .B(n11586), .C(n11587), .D(n11588), .Y(n11584)
         );
  NAND2X1 U12032 ( .A(G21581), .B(n10224), .Y(n11588) );
  NAND2X1 U12033 ( .A(G21772), .B(n9260), .Y(n11587) );
  NAND2X1 U12034 ( .A(n7246), .B(n10272), .Y(n11586) );
  ADDHXL U12035 ( .A(n11557), .B(n11589), .S(n7246) );
  AND2X1 U12036 ( .A(n11554), .B(n11556), .Y(n11589) );
  NAND2X1 U12037 ( .A(n11590), .B(n11591), .Y(n11556) );
  NAND2X1 U12038 ( .A(n9755), .B(n11498), .Y(n11591) );
  ADDHXL U12039 ( .A(n10227), .B(n11592), .S(n11590) );
  NAND3X1 U12040 ( .A(n11498), .B(n11592), .C(n9755), .Y(n11554) );
  NAND4X1 U12041 ( .A(n11593), .B(n11594), .C(n11595), .D(n11596), .Y(n11592)
         );
  NAND2X1 U12042 ( .A(G21613), .B(n7564), .Y(n11596) );
  NAND2X1 U12043 ( .A(G21708), .B(n10236), .Y(n11595) );
  NAND2X1 U12044 ( .A(G21740), .B(n10333), .Y(n11594) );
  NAND2X1 U12045 ( .A(G21581), .B(n10503), .Y(n11593) );
  NAND4X1 U12046 ( .A(n11597), .B(n11598), .C(n11599), .D(n11600), .Y(n11498)
         );
  NOR4X1 U12047 ( .A(n11601), .B(n11602), .C(n11603), .D(n11604), .Y(n11600)
         );
  NOR2X1 U12048 ( .A(n10390), .B(n11522), .Y(n11604) );
  NOR2X1 U12049 ( .A(n10391), .B(n11523), .Y(n11603) );
  NOR2X1 U12050 ( .A(n10392), .B(n11524), .Y(n11602) );
  NOR2X1 U12051 ( .A(n10398), .B(n11525), .Y(n11601) );
  NOR4X1 U12052 ( .A(n11605), .B(n11606), .C(n11607), .D(n11608), .Y(n11599)
         );
  NOR2X1 U12053 ( .A(n10399), .B(n11530), .Y(n11608) );
  NOR2X1 U12054 ( .A(n10400), .B(n11531), .Y(n11607) );
  NOR2X1 U12055 ( .A(n10407), .B(n11532), .Y(n11606) );
  NOR2X1 U12056 ( .A(n10409), .B(n11533), .Y(n11605) );
  NOR4X1 U12057 ( .A(n11609), .B(n11610), .C(n11611), .D(n11612), .Y(n11598)
         );
  NOR2X1 U12058 ( .A(n10411), .B(n11538), .Y(n11612) );
  NOR2X1 U12059 ( .A(n10419), .B(n11539), .Y(n11611) );
  NOR2X1 U12060 ( .A(n10421), .B(n11540), .Y(n11610) );
  NOR2X1 U12061 ( .A(n10423), .B(n11541), .Y(n11609) );
  NOR4X1 U12062 ( .A(n11613), .B(n11614), .C(n11615), .D(n11616), .Y(n11597)
         );
  NOR2X1 U12063 ( .A(n10389), .B(n11546), .Y(n11616) );
  NOR2X1 U12064 ( .A(n10397), .B(n11547), .Y(n11615) );
  NOR2X1 U12065 ( .A(n10405), .B(n11548), .Y(n11614) );
  NOR2X1 U12066 ( .A(n10417), .B(n11549), .Y(n11613) );
  NAND2X1 U12067 ( .A(n11617), .B(n11618), .Y(n11557) );
  NAND2X1 U12068 ( .A(n11619), .B(n11620), .Y(n11618) );
  NAND2X1 U12069 ( .A(G21613), .B(n10225), .Y(n11585) );
  NAND2X1 U12070 ( .A(n11621), .B(n11622), .Y(n11583) );
  INVX1 U12071 ( .A(n11623), .Y(n11621) );
  NAND4X1 U12072 ( .A(n11624), .B(n11625), .C(n11626), .D(n11627), .Y(G1002)
         );
  NOR2X1 U12073 ( .A(n11628), .B(n11629), .Y(n11627) );
  NOR2X1 U12074 ( .A(n6891), .B(n9506), .Y(n11629) );
  NOR2X1 U12075 ( .A(n6901), .B(n7260), .Y(n11628) );
  NAND2X1 U12076 ( .A(n7263), .B(n6882), .Y(n11626) );
  NAND2X1 U12077 ( .A(n6903), .B(n7261), .Y(n11625) );
  ADDFXL U12078 ( .A(n9926), .B(n11568), .CI(n11567), .S(n7261) );
  NAND2X1 U12079 ( .A(n11630), .B(n11631), .Y(n11567) );
  NAND2X1 U12080 ( .A(n9926), .B(n11632), .Y(n11631) );
  OR2X1 U12081 ( .A(n11633), .B(n11634), .Y(n11632) );
  NAND2X1 U12082 ( .A(n11634), .B(n11633), .Y(n11630) );
  NAND4X1 U12083 ( .A(n11635), .B(n11636), .C(n11637), .D(n11638), .Y(n11568)
         );
  NOR2X1 U12084 ( .A(n11639), .B(n11640), .Y(n11638) );
  NOR2X1 U12085 ( .A(n10216), .B(n7257), .Y(n11640) );
  NOR2X1 U12086 ( .A(n10226), .B(n7260), .Y(n11639) );
  NAND2X1 U12087 ( .A(n7263), .B(n9926), .Y(n11637) );
  NAND2X1 U12088 ( .A(n10256), .B(n11641), .Y(n11636) );
  ADDFXL U12089 ( .A(n7262), .B(n11578), .CI(n11580), .S(n11641) );
  NAND2X1 U12090 ( .A(n11642), .B(n11643), .Y(n11580) );
  NAND2X1 U12091 ( .A(n11644), .B(n11645), .Y(n11643) );
  OR2X1 U12092 ( .A(n9515), .B(n11646), .Y(n11645) );
  INVX1 U12093 ( .A(n11647), .Y(n11644) );
  NAND2X1 U12094 ( .A(n11646), .B(n9515), .Y(n11642) );
  INVX1 U12095 ( .A(n11648), .Y(n11578) );
  NAND2X1 U12096 ( .A(n7262), .B(n11499), .Y(n11635) );
  NAND2X1 U12097 ( .A(n7262), .B(n6905), .Y(n11624) );
  INVX1 U12098 ( .A(n9505), .Y(n7262) );
  ADDHXL U12099 ( .A(n11622), .B(n11623), .S(n9505) );
  ADDHXL U12100 ( .A(n9085), .B(n11649), .S(n11622) );
  NOR4X1 U12101 ( .A(n11650), .B(n11651), .C(n11652), .D(n11653), .Y(n11649)
         );
  NOR2X1 U12102 ( .A(n10227), .B(n7260), .Y(n11653) );
  INVX1 U12103 ( .A(G21771), .Y(n7260) );
  NOR2X1 U12104 ( .A(n10271), .B(n9506), .Y(n11652) );
  INVX1 U12105 ( .A(G21612), .Y(n9506) );
  NOR2X1 U12106 ( .A(n10426), .B(n7257), .Y(n11651) );
  INVX1 U12107 ( .A(G21580), .Y(n7257) );
  AND2X1 U12108 ( .A(n10272), .B(n7263), .Y(n11650) );
  ADDHXL U12109 ( .A(n11620), .B(n11654), .S(n7263) );
  AND2X1 U12110 ( .A(n11619), .B(n11617), .Y(n11654) );
  NAND3X1 U12111 ( .A(n11655), .B(n11648), .C(n9755), .Y(n11617) );
  NAND2X1 U12112 ( .A(n11656), .B(n11657), .Y(n11619) );
  NAND2X1 U12113 ( .A(n9755), .B(n11648), .Y(n11657) );
  NAND4X1 U12114 ( .A(n11658), .B(n11659), .C(n11660), .D(n11661), .Y(n11648)
         );
  NOR4X1 U12115 ( .A(n11662), .B(n11663), .C(n11664), .D(n11665), .Y(n11661)
         );
  NOR2X1 U12116 ( .A(n11100), .B(n11539), .Y(n11665) );
  NOR2X1 U12117 ( .A(n11116), .B(n11549), .Y(n11664) );
  NOR2X1 U12118 ( .A(n11115), .B(n11548), .Y(n11663) );
  NOR2X1 U12119 ( .A(n10499), .B(n11547), .Y(n11662) );
  NOR4X1 U12120 ( .A(n11666), .B(n11667), .C(n11668), .D(n11669), .Y(n11660)
         );
  NOR2X1 U12121 ( .A(n11097), .B(n11532), .Y(n11669) );
  NOR2X1 U12122 ( .A(n10502), .B(n11531), .Y(n11668) );
  NOR2X1 U12123 ( .A(n11106), .B(n11541), .Y(n11667) );
  NOR2X1 U12124 ( .A(n11105), .B(n11540), .Y(n11666) );
  NOR4X1 U12125 ( .A(n11670), .B(n11671), .C(n11672), .D(n11673), .Y(n11659)
         );
  NOR2X1 U12126 ( .A(n10500), .B(n11525), .Y(n11673) );
  NOR2X1 U12127 ( .A(n10494), .B(n11524), .Y(n11672) );
  NOR2X1 U12128 ( .A(n10493), .B(n11523), .Y(n11671) );
  NOR2X1 U12129 ( .A(n11098), .B(n11533), .Y(n11670) );
  NOR4X1 U12130 ( .A(n11674), .B(n11675), .C(n11676), .D(n11677), .Y(n11658)
         );
  NOR2X1 U12131 ( .A(n10491), .B(n11546), .Y(n11677) );
  NOR2X1 U12132 ( .A(n10492), .B(n11522), .Y(n11676) );
  NOR2X1 U12133 ( .A(n10501), .B(n11530), .Y(n11675) );
  NOR2X1 U12134 ( .A(n11099), .B(n11538), .Y(n11674) );
  ADDHXL U12135 ( .A(n10227), .B(n11655), .S(n11656) );
  NAND4X1 U12136 ( .A(n11678), .B(n11679), .C(n11680), .D(n11681), .Y(n11655)
         );
  NAND2X1 U12137 ( .A(G21612), .B(n7564), .Y(n11681) );
  NAND2X1 U12138 ( .A(G21707), .B(n10236), .Y(n11680) );
  NAND2X1 U12139 ( .A(G21739), .B(n10333), .Y(n11679) );
  NAND2X1 U12140 ( .A(G21580), .B(n10503), .Y(n11678) );
  NAND2X1 U12141 ( .A(n11682), .B(n11683), .Y(n11620) );
  NAND2X1 U12142 ( .A(n11684), .B(n11685), .Y(n11683) );
  NAND4X1 U12143 ( .A(n11686), .B(n11687), .C(n11688), .D(n11689), .Y(G1001)
         );
  NOR2X1 U12144 ( .A(n11690), .B(n11691), .Y(n11689) );
  NOR2X1 U12145 ( .A(n6891), .B(n9516), .Y(n11691) );
  NOR2X1 U12146 ( .A(n6901), .B(n7272), .Y(n11690) );
  NAND2X1 U12147 ( .A(n7275), .B(n6882), .Y(n11688) );
  NAND2X1 U12148 ( .A(n6903), .B(n7273), .Y(n11687) );
  ADDFXL U12149 ( .A(n9926), .B(n11634), .CI(n11633), .S(n7273) );
  NAND2X1 U12150 ( .A(n11692), .B(n11693), .Y(n11633) );
  NAND2X1 U12151 ( .A(n9926), .B(n11694), .Y(n11693) );
  NAND2X1 U12152 ( .A(n11695), .B(n11696), .Y(n11694) );
  NAND2X1 U12153 ( .A(n11697), .B(n11698), .Y(n11692) );
  NAND4X1 U12154 ( .A(n11699), .B(n11700), .C(n11701), .D(n11702), .Y(n11634)
         );
  NOR2X1 U12155 ( .A(n11703), .B(n11704), .Y(n11702) );
  NOR2X1 U12156 ( .A(n10216), .B(n7254), .Y(n11704) );
  INVX1 U12157 ( .A(n10444), .Y(n10216) );
  NOR2X1 U12158 ( .A(n10226), .B(n7272), .Y(n11703) );
  INVX1 U12159 ( .A(n11705), .Y(n10226) );
  NAND2X1 U12160 ( .A(n7275), .B(n9926), .Y(n11701) );
  ADDFXL U12161 ( .A(n11647), .B(n9515), .CI(n11646), .S(n11706) );
  NAND2X1 U12162 ( .A(n11707), .B(n11708), .Y(n11646) );
  NAND2X1 U12163 ( .A(n11709), .B(n11710), .Y(n11708) );
  OR2X1 U12164 ( .A(n11711), .B(n9525), .Y(n11710) );
  NAND2X1 U12165 ( .A(n9525), .B(n11711), .Y(n11707) );
  NAND2X1 U12166 ( .A(n7274), .B(n11499), .Y(n11699) );
  INVX1 U12167 ( .A(n10217), .Y(n11499) );
  NAND2X1 U12168 ( .A(n7274), .B(n6905), .Y(n11686) );
  INVX1 U12169 ( .A(n9515), .Y(n7274) );
  NAND2X1 U12170 ( .A(n11712), .B(n11623), .Y(n9515) );
  NAND3X1 U12171 ( .A(n11713), .B(n11714), .C(n11715), .Y(n11623) );
  INVX1 U12172 ( .A(n11716), .Y(n11713) );
  NAND2X1 U12173 ( .A(n11716), .B(n11717), .Y(n11712) );
  NAND2X1 U12174 ( .A(n11715), .B(n11714), .Y(n11717) );
  ADDHXL U12175 ( .A(n7564), .B(n11718), .S(n11716) );
  NOR4X1 U12176 ( .A(n11719), .B(n11720), .C(n11721), .D(n11722), .Y(n11718)
         );
  NOR2X1 U12177 ( .A(n10227), .B(n7272), .Y(n11722) );
  INVX1 U12178 ( .A(G21770), .Y(n7272) );
  NOR2X1 U12179 ( .A(n10271), .B(n9516), .Y(n11721) );
  INVX1 U12180 ( .A(G21611), .Y(n9516) );
  NOR2X1 U12181 ( .A(n10426), .B(n7254), .Y(n11720) );
  INVX1 U12182 ( .A(G21579), .Y(n7254) );
  AND2X1 U12183 ( .A(n10272), .B(n7275), .Y(n11719) );
  ADDHXL U12184 ( .A(n11685), .B(n11723), .S(n7275) );
  AND2X1 U12185 ( .A(n11684), .B(n11682), .Y(n11723) );
  NAND3X1 U12186 ( .A(n11724), .B(n11647), .C(n9755), .Y(n11682) );
  NAND2X1 U12187 ( .A(n11725), .B(n11726), .Y(n11684) );
  NAND2X1 U12188 ( .A(n9755), .B(n11647), .Y(n11726) );
  NAND4X1 U12189 ( .A(n11727), .B(n11728), .C(n11729), .D(n11730), .Y(n11647)
         );
  NOR4X1 U12190 ( .A(n11731), .B(n11732), .C(n11733), .D(n11734), .Y(n11730)
         );
  NOR2X1 U12191 ( .A(n10581), .B(n11539), .Y(n11734) );
  NOR2X1 U12192 ( .A(n10580), .B(n11549), .Y(n11733) );
  NOR2X1 U12193 ( .A(n10572), .B(n11548), .Y(n11732) );
  NOR2X1 U12194 ( .A(n10564), .B(n11547), .Y(n11731) );
  NOR4X1 U12195 ( .A(n11735), .B(n11736), .C(n11737), .D(n11738), .Y(n11729)
         );
  NOR2X1 U12196 ( .A(n10573), .B(n11532), .Y(n11738) );
  NOR2X1 U12197 ( .A(n10567), .B(n11531), .Y(n11737) );
  NOR2X1 U12198 ( .A(n10583), .B(n11541), .Y(n11736) );
  NOR2X1 U12199 ( .A(n10582), .B(n11540), .Y(n11735) );
  NOR4X1 U12200 ( .A(n11739), .B(n11740), .C(n11741), .D(n11742), .Y(n11728)
         );
  NOR2X1 U12201 ( .A(n10565), .B(n11525), .Y(n11742) );
  NOR2X1 U12202 ( .A(n10559), .B(n11524), .Y(n11741) );
  NOR2X1 U12203 ( .A(n10558), .B(n11523), .Y(n11740) );
  NOR2X1 U12204 ( .A(n10574), .B(n11533), .Y(n11739) );
  NOR4X1 U12205 ( .A(n11743), .B(n11744), .C(n11745), .D(n11746), .Y(n11727)
         );
  NOR2X1 U12206 ( .A(n10556), .B(n11546), .Y(n11746) );
  NOR2X1 U12207 ( .A(n10557), .B(n11522), .Y(n11745) );
  NOR2X1 U12208 ( .A(n10566), .B(n11530), .Y(n11744) );
  NOR2X1 U12209 ( .A(n10575), .B(n11538), .Y(n11743) );
  ADDHXL U12210 ( .A(n10227), .B(n11724), .S(n11725) );
  NAND4X1 U12211 ( .A(n11747), .B(n11748), .C(n11749), .D(n11750), .Y(n11724)
         );
  NAND2X1 U12212 ( .A(G21611), .B(n7564), .Y(n11750) );
  NAND2X1 U12213 ( .A(G21706), .B(n10236), .Y(n11749) );
  NAND2X1 U12214 ( .A(G21738), .B(n10333), .Y(n11748) );
  NAND2X1 U12215 ( .A(G21579), .B(n10503), .Y(n11747) );
  NAND2X1 U12216 ( .A(n11751), .B(n11752), .Y(n11685) );
  NAND2X1 U12217 ( .A(n11753), .B(n11754), .Y(n11752) );
  NAND4X1 U12218 ( .A(n11755), .B(n11756), .C(n11757), .D(n11758), .Y(G1000)
         );
  NOR2X1 U12219 ( .A(n11759), .B(n11760), .Y(n11758) );
  NOR2X1 U12220 ( .A(n6891), .B(n9526), .Y(n11760) );
  INVX1 U12221 ( .A(G21610), .Y(n9526) );
  NOR2X1 U12222 ( .A(n6887), .B(n9525), .Y(n11759) );
  NAND2X1 U12223 ( .A(G21769), .B(n6890), .Y(n11757) );
  INVX1 U12224 ( .A(n6901), .Y(n6890) );
  NAND2X1 U12225 ( .A(n8798), .B(n6891), .Y(n6901) );
  NAND2X1 U12226 ( .A(n7289), .B(n6903), .Y(n11756) );
  NAND2X1 U12227 ( .A(G21428), .B(n6891), .Y(n6889) );
  AND2X1 U12228 ( .A(n11761), .B(n11762), .Y(n7289) );
  NAND2X1 U12229 ( .A(n11763), .B(n9908), .Y(n11762) );
  ADDHXL U12230 ( .A(n9909), .B(n11698), .S(n11763) );
  NAND2X1 U12231 ( .A(n11764), .B(n9926), .Y(n11761) );
  ADDHXL U12232 ( .A(n11695), .B(n11696), .S(n11764) );
  NOR2X1 U12233 ( .A(n9911), .B(n11697), .Y(n11696) );
  INVX1 U12234 ( .A(n9909), .Y(n11697) );
  NAND2X1 U12235 ( .A(n11765), .B(n11766), .Y(n9909) );
  NAND2X1 U12236 ( .A(n11767), .B(n9908), .Y(n11766) );
  NAND2X1 U12237 ( .A(n9912), .B(n9911), .Y(n11767) );
  NOR2X1 U12238 ( .A(n9924), .B(n9925), .Y(n9912) );
  NAND2X1 U12239 ( .A(n9924), .B(n9925), .Y(n11765) );
  INVX1 U12240 ( .A(n9921), .Y(n9925) );
  NAND2X1 U12241 ( .A(n11768), .B(n11769), .Y(n9921) );
  NAND2X1 U12242 ( .A(n9926), .B(n11770), .Y(n11769) );
  OR2X1 U12243 ( .A(n9932), .B(n9931), .Y(n11770) );
  NAND2X1 U12244 ( .A(n9931), .B(n9932), .Y(n11768) );
  NAND2X1 U12245 ( .A(n9939), .B(n11771), .Y(n9932) );
  NAND2X1 U12246 ( .A(n9937), .B(n9940), .Y(n11771) );
  OR2X1 U12247 ( .A(n11772), .B(n11773), .Y(n9940) );
  NAND2X1 U12248 ( .A(n9949), .B(n9948), .Y(n9937) );
  NAND2X1 U12249 ( .A(n11774), .B(n11775), .Y(n9948) );
  ADDHXL U12250 ( .A(n11776), .B(n9926), .S(n11774) );
  NAND2X1 U12251 ( .A(n9953), .B(n11777), .Y(n9949) );
  NAND2X1 U12252 ( .A(n9952), .B(n9951), .Y(n11777) );
  NAND2X1 U12253 ( .A(n11778), .B(n11779), .Y(n9951) );
  NAND2X1 U12254 ( .A(n9960), .B(n9958), .Y(n9952) );
  NAND2X1 U12255 ( .A(n9967), .B(n11780), .Y(n9958) );
  NAND2X1 U12256 ( .A(n9968), .B(n9965), .Y(n11780) );
  NAND2X1 U12257 ( .A(n9977), .B(n11781), .Y(n9965) );
  NAND2X1 U12258 ( .A(n9979), .B(n9978), .Y(n11781) );
  NAND2X1 U12259 ( .A(n11782), .B(n11783), .Y(n9978) );
  ADDHXL U12260 ( .A(n9908), .B(n11784), .S(n11783) );
  INVX1 U12261 ( .A(n11785), .Y(n11782) );
  NAND2X1 U12262 ( .A(n9992), .B(n9989), .Y(n9979) );
  NAND2X1 U12263 ( .A(n11786), .B(n11787), .Y(n9989) );
  ADDHXL U12264 ( .A(n11788), .B(n9926), .S(n11786) );
  NAND2X1 U12265 ( .A(n9990), .B(n11789), .Y(n9992) );
  NAND2X1 U12266 ( .A(n9988), .B(n9987), .Y(n11789) );
  NAND2X1 U12267 ( .A(n11790), .B(n11791), .Y(n9987) );
  NAND2X1 U12268 ( .A(n9999), .B(n9997), .Y(n9988) );
  NAND2X1 U12269 ( .A(n10007), .B(n11792), .Y(n9997) );
  OR2X1 U12270 ( .A(n9908), .B(n10006), .Y(n11792) );
  NOR2X1 U12271 ( .A(n11793), .B(n11794), .Y(n10006) );
  NAND2X1 U12272 ( .A(n11794), .B(n11793), .Y(n10007) );
  NAND4X1 U12273 ( .A(n11795), .B(n11796), .C(n11797), .D(n11798), .Y(n11793)
         );
  NOR2X1 U12274 ( .A(n11799), .B(n7456), .Y(n11798) );
  NOR2X1 U12275 ( .A(n7421), .B(n9908), .Y(n11799) );
  NAND2X1 U12276 ( .A(G21567), .B(n10444), .Y(n11797) );
  NAND2X1 U12277 ( .A(n7003), .B(n11800), .Y(n11796) );
  NAND2X1 U12278 ( .A(n11705), .B(G21758), .Y(n11795) );
  ADDHXL U12279 ( .A(n9926), .B(n11801), .S(n11794) );
  NAND4X1 U12280 ( .A(n11802), .B(n9193), .C(n11803), .D(n11804), .Y(n11801)
         );
  NOR4X1 U12281 ( .A(n11805), .B(n11806), .C(n11807), .D(n11808), .Y(n11804)
         );
  AND2X1 U12282 ( .A(n11414), .B(n11809), .Y(n11807) );
  NAND4X1 U12283 ( .A(n11810), .B(n11811), .C(n11812), .D(n11813), .Y(n11414)
         );
  NOR4X1 U12284 ( .A(n11814), .B(n11815), .C(n11816), .D(n11817), .Y(n11813)
         );
  NOR2X1 U12285 ( .A(n10907), .B(n11818), .Y(n11817) );
  NOR2X1 U12286 ( .A(n10909), .B(n11819), .Y(n11816) );
  NOR2X1 U12287 ( .A(n10911), .B(n11820), .Y(n11815) );
  NOR2X1 U12288 ( .A(n10918), .B(n11821), .Y(n11814) );
  NOR4X1 U12289 ( .A(n11822), .B(n11823), .C(n11824), .D(n11825), .Y(n11812)
         );
  NOR2X1 U12290 ( .A(n10919), .B(n11826), .Y(n11825) );
  NOR2X1 U12291 ( .A(n10922), .B(n11827), .Y(n11824) );
  NOR2X1 U12292 ( .A(n10941), .B(n11828), .Y(n11823) );
  NOR2X1 U12293 ( .A(n10940), .B(n11829), .Y(n11822) );
  NOR4X1 U12294 ( .A(n11830), .B(n11831), .C(n11832), .D(n11833), .Y(n11811)
         );
  NOR2X1 U12295 ( .A(n10939), .B(n11834), .Y(n11833) );
  NOR2X1 U12296 ( .A(n10931), .B(n11835), .Y(n11832) );
  NOR2X1 U12297 ( .A(n10929), .B(n11836), .Y(n11831) );
  NOR2X1 U12298 ( .A(n10927), .B(n11837), .Y(n11830) );
  NOR4X1 U12299 ( .A(n11838), .B(n11839), .C(n11840), .D(n11841), .Y(n11810)
         );
  NOR2X1 U12300 ( .A(n10904), .B(n11842), .Y(n11841) );
  NOR2X1 U12301 ( .A(n10916), .B(n11843), .Y(n11840) );
  NOR2X1 U12302 ( .A(n10942), .B(n11844), .Y(n11839) );
  NOR2X1 U12303 ( .A(n10932), .B(n11845), .Y(n11838) );
  NOR2X1 U12304 ( .A(n11846), .B(n11847), .Y(n11806) );
  NOR4X1 U12305 ( .A(n11848), .B(n11849), .C(n11850), .D(n11851), .Y(n11846)
         );
  NAND4X1 U12306 ( .A(n11852), .B(n11853), .C(n11854), .D(n11855), .Y(n11851)
         );
  NAND2X1 U12307 ( .A(n7813), .B(G21532), .Y(n11855) );
  INVX1 U12308 ( .A(n7816), .Y(n7813) );
  NAND2X1 U12309 ( .A(n8131), .B(G21500), .Y(n11854) );
  INVX1 U12310 ( .A(n8134), .Y(n8131) );
  NAND2X1 U12311 ( .A(n8446), .B(G21468), .Y(n11853) );
  INVX1 U12312 ( .A(n8449), .Y(n8446) );
  NAND2X1 U12313 ( .A(n8788), .B(G21436), .Y(n11852) );
  INVX1 U12314 ( .A(n8803), .Y(n8788) );
  NAND4X1 U12315 ( .A(n11856), .B(n11857), .C(n11858), .D(n11859), .Y(n11850)
         );
  NAND2X1 U12316 ( .A(n7565), .B(G21556), .Y(n11859) );
  INVX1 U12317 ( .A(n7570), .Y(n7565) );
  NAND2X1 U12318 ( .A(n7653), .B(G21548), .Y(n11858) );
  INVX1 U12319 ( .A(n7656), .Y(n7653) );
  NAND2X1 U12320 ( .A(n7733), .B(G21540), .Y(n11857) );
  INVX1 U12321 ( .A(n7736), .Y(n7733) );
  NAND2X1 U12322 ( .A(n7895), .B(G21524), .Y(n11856) );
  INVX1 U12323 ( .A(n7898), .Y(n7895) );
  NAND4X1 U12324 ( .A(n11860), .B(n11861), .C(n11862), .D(n11863), .Y(n11849)
         );
  NAND2X1 U12325 ( .A(n7975), .B(G21516), .Y(n11863) );
  INVX1 U12326 ( .A(n7978), .Y(n7975) );
  NAND2X1 U12327 ( .A(n8053), .B(G21508), .Y(n11862) );
  INVX1 U12328 ( .A(n8056), .Y(n8053) );
  NAND2X1 U12329 ( .A(n8210), .B(G21492), .Y(n11861) );
  INVX1 U12330 ( .A(n8213), .Y(n8210) );
  NAND2X1 U12331 ( .A(n8290), .B(G21484), .Y(n11860) );
  INVX1 U12332 ( .A(n8293), .Y(n8290) );
  NAND4X1 U12333 ( .A(n11864), .B(n11865), .C(n11866), .D(n11867), .Y(n11848)
         );
  NAND2X1 U12334 ( .A(n8368), .B(G21476), .Y(n11867) );
  INVX1 U12335 ( .A(n8371), .Y(n8368) );
  NAND2X1 U12336 ( .A(n8525), .B(G21460), .Y(n11866) );
  INVX1 U12337 ( .A(n8528), .Y(n8525) );
  NAND2X1 U12338 ( .A(n8607), .B(G21452), .Y(n11865) );
  INVX1 U12339 ( .A(n8610), .Y(n8607) );
  NAND2X1 U12340 ( .A(n8685), .B(G21444), .Y(n11864) );
  INVX1 U12341 ( .A(n8688), .Y(n8685) );
  NOR2X1 U12342 ( .A(n7439), .B(n8890), .Y(n11805) );
  NAND2X1 U12343 ( .A(n10256), .B(n11868), .Y(n11803) );
  NAND4X1 U12344 ( .A(n11869), .B(n11870), .C(n11871), .D(n11872), .Y(n11868)
         );
  NOR4X1 U12345 ( .A(n11873), .B(n11874), .C(n11875), .D(n11876), .Y(n11872)
         );
  NOR2X1 U12346 ( .A(n10904), .B(n11877), .Y(n11876) );
  NOR2X1 U12347 ( .A(n10907), .B(n11878), .Y(n11875) );
  NOR2X1 U12348 ( .A(n10909), .B(n11879), .Y(n11874) );
  NOR2X1 U12349 ( .A(n10911), .B(n11880), .Y(n11873) );
  NOR4X1 U12350 ( .A(n11881), .B(n11882), .C(n11883), .D(n11884), .Y(n11871)
         );
  NOR2X1 U12351 ( .A(n10916), .B(n11885), .Y(n11884) );
  NOR2X1 U12352 ( .A(n10918), .B(n11886), .Y(n11883) );
  NOR2X1 U12353 ( .A(n10919), .B(n11887), .Y(n11882) );
  NOR2X1 U12354 ( .A(n10922), .B(n11888), .Y(n11881) );
  NOR4X1 U12355 ( .A(n11889), .B(n11890), .C(n11891), .D(n11892), .Y(n11870)
         );
  NOR2X1 U12356 ( .A(n10942), .B(n11893), .Y(n11892) );
  NOR2X1 U12357 ( .A(n10941), .B(n11894), .Y(n11891) );
  NOR2X1 U12358 ( .A(n10940), .B(n11895), .Y(n11890) );
  NOR2X1 U12359 ( .A(n10939), .B(n11896), .Y(n11889) );
  NOR4X1 U12360 ( .A(n11897), .B(n11898), .C(n11899), .D(n11900), .Y(n11869)
         );
  NOR2X1 U12361 ( .A(n10932), .B(n11901), .Y(n11900) );
  NOR2X1 U12362 ( .A(n10931), .B(n11902), .Y(n11899) );
  NOR2X1 U12363 ( .A(n10929), .B(n11903), .Y(n11898) );
  NOR2X1 U12364 ( .A(n10927), .B(n11904), .Y(n11897) );
  NAND4X1 U12365 ( .A(n11905), .B(n11906), .C(n11907), .D(n11908), .Y(n11802)
         );
  NOR4X1 U12366 ( .A(n11909), .B(n11910), .C(n11911), .D(n11912), .Y(n11908)
         );
  NOR2X1 U12367 ( .A(n10941), .B(n11913), .Y(n11912) );
  NOR2X1 U12368 ( .A(n10940), .B(n11914), .Y(n11911) );
  NAND2X1 U12369 ( .A(n11915), .B(n11916), .Y(n11910) );
  NAND2X1 U12370 ( .A(n11917), .B(G21540), .Y(n11916) );
  NAND2X1 U12371 ( .A(n11918), .B(G21548), .Y(n11915) );
  NOR2X1 U12372 ( .A(n10932), .B(n11919), .Y(n11909) );
  NOR4X1 U12373 ( .A(n11920), .B(n11921), .C(n11922), .D(n11923), .Y(n11907)
         );
  NOR2X1 U12374 ( .A(n10942), .B(n11924), .Y(n11923) );
  NOR2X1 U12375 ( .A(n10907), .B(n11925), .Y(n11922) );
  NOR2X1 U12376 ( .A(n10909), .B(n11926), .Y(n11921) );
  NOR2X1 U12377 ( .A(n10911), .B(n11927), .Y(n11920) );
  NOR4X1 U12378 ( .A(n11928), .B(n11929), .C(n11930), .D(n11931), .Y(n11906)
         );
  NOR2X1 U12379 ( .A(n10918), .B(n11932), .Y(n11931) );
  NOR2X1 U12380 ( .A(n10919), .B(n11933), .Y(n11930) );
  NOR2X1 U12381 ( .A(n10922), .B(n11934), .Y(n11929) );
  NOR2X1 U12382 ( .A(n10927), .B(n11935), .Y(n11928) );
  NOR4X1 U12383 ( .A(n11936), .B(n11937), .C(n11938), .D(n9908), .Y(n11905) );
  NOR2X1 U12384 ( .A(n10904), .B(n11939), .Y(n11938) );
  NOR2X1 U12385 ( .A(n10916), .B(n11940), .Y(n11937) );
  NOR2X1 U12386 ( .A(n10939), .B(n11941), .Y(n11936) );
  OR2X1 U12387 ( .A(n11791), .B(n11790), .Y(n9999) );
  ADDHXL U12388 ( .A(n11942), .B(n9926), .S(n11790) );
  NAND4X1 U12389 ( .A(n11943), .B(n11944), .C(n11945), .D(n11946), .Y(n11942)
         );
  NOR4X1 U12390 ( .A(n9195), .B(n11947), .C(n11948), .D(n11949), .Y(n11946) );
  NOR2X1 U12391 ( .A(n11950), .B(n9192), .Y(n11949) );
  NOR4X1 U12392 ( .A(n11951), .B(n11952), .C(n11953), .D(n11954), .Y(n11950)
         );
  NAND4X1 U12393 ( .A(n11955), .B(n11956), .C(n11957), .D(n11958), .Y(n11954)
         );
  NAND2X1 U12394 ( .A(n11959), .B(G21555), .Y(n11958) );
  NAND2X1 U12395 ( .A(n11960), .B(G21547), .Y(n11957) );
  NAND2X1 U12396 ( .A(n11961), .B(G21539), .Y(n11956) );
  NAND2X1 U12397 ( .A(n11962), .B(G21531), .Y(n11955) );
  NAND4X1 U12398 ( .A(n11963), .B(n11964), .C(n11965), .D(n11966), .Y(n11953)
         );
  NAND2X1 U12399 ( .A(n11967), .B(G21523), .Y(n11966) );
  NAND2X1 U12400 ( .A(n11968), .B(G21515), .Y(n11965) );
  NAND2X1 U12401 ( .A(n11969), .B(G21507), .Y(n11964) );
  NAND2X1 U12402 ( .A(n11970), .B(G21499), .Y(n11963) );
  NAND4X1 U12403 ( .A(n11971), .B(n11972), .C(n11973), .D(n11974), .Y(n11952)
         );
  NAND2X1 U12404 ( .A(n11975), .B(G21491), .Y(n11974) );
  NAND2X1 U12405 ( .A(n11976), .B(G21483), .Y(n11973) );
  NAND2X1 U12406 ( .A(n11977), .B(G21475), .Y(n11972) );
  NAND2X1 U12407 ( .A(n11978), .B(G21467), .Y(n11971) );
  NAND4X1 U12408 ( .A(n11979), .B(n11980), .C(n11981), .D(n11982), .Y(n11951)
         );
  NAND2X1 U12409 ( .A(n11983), .B(G21459), .Y(n11982) );
  NAND2X1 U12410 ( .A(n11984), .B(G21451), .Y(n11981) );
  NAND2X1 U12411 ( .A(n11985), .B(G21443), .Y(n11980) );
  NAND2X1 U12412 ( .A(n11986), .B(G21435), .Y(n11979) );
  NOR2X1 U12413 ( .A(n10116), .B(n11987), .Y(n11948) );
  NOR4X1 U12414 ( .A(n11988), .B(n11989), .C(n11990), .D(n11991), .Y(n11947)
         );
  NAND4X1 U12415 ( .A(n9926), .B(n11992), .C(n11993), .D(n11994), .Y(n11991)
         );
  OR2X1 U12416 ( .A(n11941), .B(n10841), .Y(n11994) );
  OR2X1 U12417 ( .A(n11940), .B(n10825), .Y(n11993) );
  OR2X1 U12418 ( .A(n11939), .B(n10817), .Y(n11992) );
  NAND4X1 U12419 ( .A(n11995), .B(n11996), .C(n11997), .D(n11998), .Y(n11990)
         );
  OR2X1 U12420 ( .A(n11935), .B(n10833), .Y(n11998) );
  OR2X1 U12421 ( .A(n11934), .B(n10828), .Y(n11997) );
  OR2X1 U12422 ( .A(n11933), .B(n10827), .Y(n11996) );
  OR2X1 U12423 ( .A(n11932), .B(n10826), .Y(n11995) );
  NAND4X1 U12424 ( .A(n11999), .B(n12000), .C(n12001), .D(n12002), .Y(n11989)
         );
  OR2X1 U12425 ( .A(n11927), .B(n10820), .Y(n12002) );
  OR2X1 U12426 ( .A(n11926), .B(n10819), .Y(n12001) );
  OR2X1 U12427 ( .A(n11925), .B(n10818), .Y(n12000) );
  OR2X1 U12428 ( .A(n11924), .B(n10844), .Y(n11999) );
  NAND4X1 U12429 ( .A(n12003), .B(n12004), .C(n12005), .D(n12006), .Y(n11988)
         );
  OR2X1 U12430 ( .A(n11919), .B(n10836), .Y(n12006) );
  NOR2X1 U12431 ( .A(n12007), .B(n12008), .Y(n12005) );
  NOR2X1 U12432 ( .A(n10834), .B(n12009), .Y(n12008) );
  NOR2X1 U12433 ( .A(n10835), .B(n12010), .Y(n12007) );
  OR2X1 U12434 ( .A(n11914), .B(n10842), .Y(n12004) );
  OR2X1 U12435 ( .A(n11913), .B(n10843), .Y(n12003) );
  NAND2X1 U12436 ( .A(G21560), .B(n7456), .Y(n11945) );
  NAND2X1 U12437 ( .A(n12011), .B(n12012), .Y(n11944) );
  NAND4X1 U12438 ( .A(n12013), .B(n12014), .C(n12015), .D(n12016), .Y(n12012)
         );
  NOR4X1 U12439 ( .A(n12017), .B(n12018), .C(n12019), .D(n12020), .Y(n12016)
         );
  NOR2X1 U12440 ( .A(n10818), .B(n8688), .Y(n12020) );
  NOR2X1 U12441 ( .A(n10819), .B(n8610), .Y(n12019) );
  NOR2X1 U12442 ( .A(n10820), .B(n8528), .Y(n12018) );
  NOR2X1 U12443 ( .A(n10826), .B(n8371), .Y(n12017) );
  NOR4X1 U12444 ( .A(n12021), .B(n12022), .C(n12023), .D(n12024), .Y(n12015)
         );
  NOR2X1 U12445 ( .A(n10827), .B(n8293), .Y(n12024) );
  NOR2X1 U12446 ( .A(n10828), .B(n8213), .Y(n12023) );
  NOR2X1 U12447 ( .A(n10843), .B(n8056), .Y(n12022) );
  NOR2X1 U12448 ( .A(n10842), .B(n7978), .Y(n12021) );
  NOR4X1 U12449 ( .A(n12025), .B(n12026), .C(n12027), .D(n12028), .Y(n12014)
         );
  NOR2X1 U12450 ( .A(n10841), .B(n7898), .Y(n12028) );
  NOR2X1 U12451 ( .A(n10835), .B(n7736), .Y(n12027) );
  NOR2X1 U12452 ( .A(n10834), .B(n7656), .Y(n12026) );
  NOR2X1 U12453 ( .A(n10833), .B(n7570), .Y(n12025) );
  NOR4X1 U12454 ( .A(n12029), .B(n12030), .C(n12031), .D(n12032), .Y(n12013)
         );
  NOR2X1 U12455 ( .A(n10817), .B(n8803), .Y(n12032) );
  NOR2X1 U12456 ( .A(n10825), .B(n8449), .Y(n12031) );
  NOR2X1 U12457 ( .A(n10844), .B(n8134), .Y(n12030) );
  NOR2X1 U12458 ( .A(n10836), .B(n7816), .Y(n12029) );
  NAND2X1 U12459 ( .A(n11809), .B(n11350), .Y(n11943) );
  NAND4X1 U12460 ( .A(n12033), .B(n12034), .C(n12035), .D(n12036), .Y(n11350)
         );
  NOR4X1 U12461 ( .A(n12037), .B(n12038), .C(n12039), .D(n12040), .Y(n12036)
         );
  NOR2X1 U12462 ( .A(n10818), .B(n11818), .Y(n12040) );
  NOR2X1 U12463 ( .A(n10819), .B(n11819), .Y(n12039) );
  NOR2X1 U12464 ( .A(n10820), .B(n11820), .Y(n12038) );
  NOR2X1 U12465 ( .A(n10826), .B(n11821), .Y(n12037) );
  NOR4X1 U12466 ( .A(n12041), .B(n12042), .C(n12043), .D(n12044), .Y(n12035)
         );
  NOR2X1 U12467 ( .A(n10827), .B(n11826), .Y(n12044) );
  NOR2X1 U12468 ( .A(n10828), .B(n11827), .Y(n12043) );
  NOR2X1 U12469 ( .A(n10843), .B(n11828), .Y(n12042) );
  NOR2X1 U12470 ( .A(n10842), .B(n11829), .Y(n12041) );
  NOR4X1 U12471 ( .A(n12045), .B(n12046), .C(n12047), .D(n12048), .Y(n12034)
         );
  NOR2X1 U12472 ( .A(n10841), .B(n11834), .Y(n12048) );
  NOR2X1 U12473 ( .A(n10835), .B(n11835), .Y(n12047) );
  NOR2X1 U12474 ( .A(n10834), .B(n11836), .Y(n12046) );
  NOR2X1 U12475 ( .A(n10833), .B(n11837), .Y(n12045) );
  NOR4X1 U12476 ( .A(n12049), .B(n12050), .C(n12051), .D(n12052), .Y(n12033)
         );
  NOR2X1 U12477 ( .A(n10817), .B(n11842), .Y(n12052) );
  NOR2X1 U12478 ( .A(n10825), .B(n11843), .Y(n12051) );
  NOR2X1 U12479 ( .A(n10844), .B(n11844), .Y(n12050) );
  NOR2X1 U12480 ( .A(n10836), .B(n11845), .Y(n12049) );
  NAND4X1 U12481 ( .A(n12053), .B(n12054), .C(n12055), .D(n12056), .Y(n11791)
         );
  NAND2X1 U12482 ( .A(n6992), .B(n11800), .Y(n12056) );
  NAND2X1 U12483 ( .A(n11705), .B(G21759), .Y(n12055) );
  NAND2X1 U12484 ( .A(G21568), .B(n10444), .Y(n12054) );
  NAND2X1 U12485 ( .A(n9926), .B(n6990), .Y(n12053) );
  NAND2X1 U12486 ( .A(n12057), .B(n12058), .Y(n9990) );
  ADDHXL U12487 ( .A(n9908), .B(n11788), .S(n12058) );
  NAND4X1 U12488 ( .A(n12059), .B(n12060), .C(n12061), .D(n12062), .Y(n11788)
         );
  NOR3X1 U12489 ( .A(n12063), .B(n12064), .C(n12065), .Y(n12062) );
  AND2X1 U12490 ( .A(n11213), .B(n11809), .Y(n12065) );
  NAND4X1 U12491 ( .A(n12066), .B(n12067), .C(n12068), .D(n12069), .Y(n11213)
         );
  NOR4X1 U12492 ( .A(n12070), .B(n12071), .C(n12072), .D(n12073), .Y(n12069)
         );
  NOR2X1 U12493 ( .A(n10728), .B(n11818), .Y(n12073) );
  NOR2X1 U12494 ( .A(n10729), .B(n11819), .Y(n12072) );
  NOR2X1 U12495 ( .A(n10730), .B(n11820), .Y(n12071) );
  NOR2X1 U12496 ( .A(n10736), .B(n11821), .Y(n12070) );
  NOR4X1 U12497 ( .A(n12074), .B(n12075), .C(n12076), .D(n12077), .Y(n12068)
         );
  NOR2X1 U12498 ( .A(n10737), .B(n11826), .Y(n12077) );
  NOR2X1 U12499 ( .A(n10738), .B(n11827), .Y(n12076) );
  NOR2X1 U12500 ( .A(n10753), .B(n11828), .Y(n12075) );
  NOR2X1 U12501 ( .A(n10752), .B(n11829), .Y(n12074) );
  NOR4X1 U12502 ( .A(n12078), .B(n12079), .C(n12080), .D(n12081), .Y(n12067)
         );
  NOR2X1 U12503 ( .A(n10751), .B(n11834), .Y(n12081) );
  NOR2X1 U12504 ( .A(n10745), .B(n11835), .Y(n12080) );
  NOR2X1 U12505 ( .A(n10744), .B(n11836), .Y(n12079) );
  NOR2X1 U12506 ( .A(n10743), .B(n11837), .Y(n12078) );
  NOR4X1 U12507 ( .A(n12082), .B(n12083), .C(n12084), .D(n12085), .Y(n12066)
         );
  NOR2X1 U12508 ( .A(n10727), .B(n11842), .Y(n12085) );
  NOR2X1 U12509 ( .A(n10735), .B(n11843), .Y(n12084) );
  NOR2X1 U12510 ( .A(n10754), .B(n11844), .Y(n12083) );
  NOR2X1 U12511 ( .A(n10746), .B(n11845), .Y(n12082) );
  NOR2X1 U12512 ( .A(n12086), .B(n9192), .Y(n12064) );
  NOR4X1 U12513 ( .A(n12087), .B(n12088), .C(n12089), .D(n12090), .Y(n12086)
         );
  NAND4X1 U12514 ( .A(n12091), .B(n12092), .C(n12093), .D(n12094), .Y(n12090)
         );
  NAND2X1 U12515 ( .A(n11959), .B(G21554), .Y(n12094) );
  NAND2X1 U12516 ( .A(n11960), .B(G21546), .Y(n12093) );
  NAND2X1 U12517 ( .A(n11961), .B(G21538), .Y(n12092) );
  NAND2X1 U12518 ( .A(n11962), .B(G21530), .Y(n12091) );
  NAND4X1 U12519 ( .A(n12095), .B(n12096), .C(n12097), .D(n12098), .Y(n12089)
         );
  NAND2X1 U12520 ( .A(n11967), .B(G21522), .Y(n12098) );
  NAND2X1 U12521 ( .A(n11968), .B(G21514), .Y(n12097) );
  NAND2X1 U12522 ( .A(n11969), .B(G21506), .Y(n12096) );
  NAND2X1 U12523 ( .A(n11970), .B(G21498), .Y(n12095) );
  NAND4X1 U12524 ( .A(n12099), .B(n12100), .C(n12101), .D(n12102), .Y(n12088)
         );
  NAND2X1 U12525 ( .A(n11975), .B(G21490), .Y(n12102) );
  NAND2X1 U12526 ( .A(n11976), .B(G21482), .Y(n12101) );
  NAND2X1 U12527 ( .A(n11977), .B(G21474), .Y(n12100) );
  NAND2X1 U12528 ( .A(n11978), .B(G21466), .Y(n12099) );
  NAND4X1 U12529 ( .A(n12103), .B(n12104), .C(n12105), .D(n12106), .Y(n12087)
         );
  NAND2X1 U12530 ( .A(n11983), .B(G21458), .Y(n12106) );
  NAND2X1 U12531 ( .A(n11984), .B(G21450), .Y(n12105) );
  NAND2X1 U12532 ( .A(n11985), .B(G21442), .Y(n12104) );
  NAND2X1 U12533 ( .A(n11986), .B(G21434), .Y(n12103) );
  NOR2X1 U12534 ( .A(n7439), .B(n8893), .Y(n12063) );
  NAND2X1 U12535 ( .A(n12011), .B(n12107), .Y(n12061) );
  NAND4X1 U12536 ( .A(n12108), .B(n12109), .C(n12110), .D(n12111), .Y(n12107)
         );
  NOR4X1 U12537 ( .A(n12112), .B(n12113), .C(n12114), .D(n12115), .Y(n12111)
         );
  NOR2X1 U12538 ( .A(n10728), .B(n8688), .Y(n12115) );
  NOR2X1 U12539 ( .A(n10729), .B(n8610), .Y(n12114) );
  NOR2X1 U12540 ( .A(n10730), .B(n8528), .Y(n12113) );
  NOR2X1 U12541 ( .A(n10736), .B(n8371), .Y(n12112) );
  NOR4X1 U12542 ( .A(n12116), .B(n12117), .C(n12118), .D(n12119), .Y(n12110)
         );
  NOR2X1 U12543 ( .A(n10737), .B(n8293), .Y(n12119) );
  NOR2X1 U12544 ( .A(n10738), .B(n8213), .Y(n12118) );
  NOR2X1 U12545 ( .A(n10753), .B(n8056), .Y(n12117) );
  NOR2X1 U12546 ( .A(n10752), .B(n7978), .Y(n12116) );
  NOR4X1 U12547 ( .A(n12120), .B(n12121), .C(n12122), .D(n12123), .Y(n12109)
         );
  NOR2X1 U12548 ( .A(n10751), .B(n7898), .Y(n12123) );
  NOR2X1 U12549 ( .A(n10745), .B(n7736), .Y(n12122) );
  NOR2X1 U12550 ( .A(n10744), .B(n7656), .Y(n12121) );
  NOR2X1 U12551 ( .A(n10743), .B(n7570), .Y(n12120) );
  NOR4X1 U12552 ( .A(n12124), .B(n12125), .C(n12126), .D(n12127), .Y(n12108)
         );
  NOR2X1 U12553 ( .A(n10727), .B(n8803), .Y(n12127) );
  NOR2X1 U12554 ( .A(n10735), .B(n8449), .Y(n12126) );
  NOR2X1 U12555 ( .A(n10754), .B(n8134), .Y(n12125) );
  NOR2X1 U12556 ( .A(n10746), .B(n7816), .Y(n12124) );
  NAND4X1 U12557 ( .A(n12128), .B(n12129), .C(n12130), .D(n12131), .Y(n12059)
         );
  NOR4X1 U12558 ( .A(n12132), .B(n12133), .C(n12134), .D(n12135), .Y(n12131)
         );
  NOR2X1 U12559 ( .A(n10753), .B(n11913), .Y(n12135) );
  NOR2X1 U12560 ( .A(n10752), .B(n11914), .Y(n12134) );
  NAND2X1 U12561 ( .A(n12136), .B(n12137), .Y(n12133) );
  NAND2X1 U12562 ( .A(n11917), .B(G21538), .Y(n12137) );
  NAND2X1 U12563 ( .A(n11918), .B(G21546), .Y(n12136) );
  NOR2X1 U12564 ( .A(n10746), .B(n11919), .Y(n12132) );
  NOR4X1 U12565 ( .A(n12138), .B(n12139), .C(n12140), .D(n12141), .Y(n12130)
         );
  NOR2X1 U12566 ( .A(n10754), .B(n11924), .Y(n12141) );
  NOR2X1 U12567 ( .A(n10728), .B(n11925), .Y(n12140) );
  NOR2X1 U12568 ( .A(n10729), .B(n11926), .Y(n12139) );
  NOR2X1 U12569 ( .A(n10730), .B(n11927), .Y(n12138) );
  NOR4X1 U12570 ( .A(n12142), .B(n12143), .C(n12144), .D(n12145), .Y(n12129)
         );
  NOR2X1 U12571 ( .A(n10736), .B(n11932), .Y(n12145) );
  NOR2X1 U12572 ( .A(n10737), .B(n11933), .Y(n12144) );
  NOR2X1 U12573 ( .A(n10738), .B(n11934), .Y(n12143) );
  NOR2X1 U12574 ( .A(n10743), .B(n11935), .Y(n12142) );
  NOR4X1 U12575 ( .A(n12146), .B(n12147), .C(n12148), .D(n9908), .Y(n12128) );
  NOR2X1 U12576 ( .A(n10727), .B(n11939), .Y(n12148) );
  NOR2X1 U12577 ( .A(n10735), .B(n11940), .Y(n12147) );
  NOR2X1 U12578 ( .A(n10751), .B(n11941), .Y(n12146) );
  INVX1 U12579 ( .A(n11787), .Y(n12057) );
  NAND4X1 U12580 ( .A(n12149), .B(n12150), .C(n12151), .D(n12152), .Y(n11787)
         );
  NAND2X1 U12581 ( .A(n11800), .B(n6981), .Y(n12152) );
  NAND2X1 U12582 ( .A(n11705), .B(G21760), .Y(n12151) );
  NAND2X1 U12583 ( .A(G21569), .B(n10444), .Y(n12150) );
  NAND2X1 U12584 ( .A(n9926), .B(n6979), .Y(n12149) );
  NAND2X1 U12585 ( .A(n12153), .B(n11785), .Y(n9977) );
  NAND4X1 U12586 ( .A(n12154), .B(n12155), .C(n12156), .D(n12157), .Y(n11785)
         );
  NAND2X1 U12587 ( .A(n6971), .B(n11800), .Y(n12157) );
  NAND2X1 U12588 ( .A(n11705), .B(G21761), .Y(n12156) );
  NAND2X1 U12589 ( .A(G21570), .B(n10444), .Y(n12155) );
  NAND2X1 U12590 ( .A(n9926), .B(n6969), .Y(n12154) );
  ADDHXL U12591 ( .A(n11784), .B(n9926), .S(n12153) );
  NAND4X1 U12592 ( .A(n12158), .B(n12159), .C(n12160), .D(n12161), .Y(n11784)
         );
  NOR2X1 U12593 ( .A(n12162), .B(n12163), .Y(n12161) );
  NOR2X1 U12594 ( .A(n7439), .B(n8870), .Y(n12163) );
  AND2X1 U12595 ( .A(n11218), .B(n11809), .Y(n12162) );
  NAND4X1 U12596 ( .A(n12164), .B(n12165), .C(n12166), .D(n12167), .Y(n11218)
         );
  NOR4X1 U12597 ( .A(n12168), .B(n12169), .C(n12170), .D(n12171), .Y(n12167)
         );
  NOR2X1 U12598 ( .A(n10639), .B(n11818), .Y(n12171) );
  NOR2X1 U12599 ( .A(n10640), .B(n11819), .Y(n12170) );
  NOR2X1 U12600 ( .A(n10641), .B(n11820), .Y(n12169) );
  NOR2X1 U12601 ( .A(n10647), .B(n11821), .Y(n12168) );
  NOR4X1 U12602 ( .A(n12172), .B(n12173), .C(n12174), .D(n12175), .Y(n12166)
         );
  NOR2X1 U12603 ( .A(n10648), .B(n11826), .Y(n12175) );
  NOR2X1 U12604 ( .A(n10649), .B(n11827), .Y(n12174) );
  NOR2X1 U12605 ( .A(n10664), .B(n11828), .Y(n12173) );
  NOR2X1 U12606 ( .A(n10663), .B(n11829), .Y(n12172) );
  NOR4X1 U12607 ( .A(n12176), .B(n12177), .C(n12178), .D(n12179), .Y(n12165)
         );
  NOR2X1 U12608 ( .A(n10662), .B(n11834), .Y(n12179) );
  NOR2X1 U12609 ( .A(n10656), .B(n11835), .Y(n12178) );
  NOR2X1 U12610 ( .A(n10655), .B(n11836), .Y(n12177) );
  NOR2X1 U12611 ( .A(n10654), .B(n11837), .Y(n12176) );
  NOR4X1 U12612 ( .A(n12180), .B(n12181), .C(n12182), .D(n12183), .Y(n12164)
         );
  NOR2X1 U12613 ( .A(n10638), .B(n11842), .Y(n12183) );
  NOR2X1 U12614 ( .A(n10646), .B(n11843), .Y(n12182) );
  NOR2X1 U12615 ( .A(n10665), .B(n11844), .Y(n12181) );
  NOR2X1 U12616 ( .A(n10657), .B(n11845), .Y(n12180) );
  NAND2X1 U12617 ( .A(n10256), .B(n12184), .Y(n12160) );
  NAND4X1 U12618 ( .A(n12185), .B(n12186), .C(n12187), .D(n12188), .Y(n12184)
         );
  NOR4X1 U12619 ( .A(n12189), .B(n12190), .C(n12191), .D(n12192), .Y(n12188)
         );
  NOR2X1 U12620 ( .A(n10638), .B(n11877), .Y(n12192) );
  NOR2X1 U12621 ( .A(n10639), .B(n11878), .Y(n12191) );
  NOR2X1 U12622 ( .A(n10640), .B(n11879), .Y(n12190) );
  NOR2X1 U12623 ( .A(n10641), .B(n11880), .Y(n12189) );
  NOR4X1 U12624 ( .A(n12193), .B(n12194), .C(n12195), .D(n12196), .Y(n12187)
         );
  NOR2X1 U12625 ( .A(n10646), .B(n11885), .Y(n12196) );
  NOR2X1 U12626 ( .A(n10647), .B(n11886), .Y(n12195) );
  NOR2X1 U12627 ( .A(n10648), .B(n11887), .Y(n12194) );
  NOR2X1 U12628 ( .A(n10649), .B(n11888), .Y(n12193) );
  NOR4X1 U12629 ( .A(n12197), .B(n12198), .C(n12199), .D(n12200), .Y(n12186)
         );
  NOR2X1 U12630 ( .A(n10665), .B(n11893), .Y(n12200) );
  NOR2X1 U12631 ( .A(n10664), .B(n11894), .Y(n12199) );
  NOR2X1 U12632 ( .A(n10663), .B(n11895), .Y(n12198) );
  NOR2X1 U12633 ( .A(n10662), .B(n11896), .Y(n12197) );
  NOR4X1 U12634 ( .A(n12201), .B(n12202), .C(n12203), .D(n12204), .Y(n12185)
         );
  NOR2X1 U12635 ( .A(n10657), .B(n11901), .Y(n12204) );
  NOR2X1 U12636 ( .A(n10656), .B(n11902), .Y(n12203) );
  NOR2X1 U12637 ( .A(n10655), .B(n11903), .Y(n12202) );
  NOR2X1 U12638 ( .A(n10654), .B(n11904), .Y(n12201) );
  NAND4X1 U12639 ( .A(n12205), .B(n12206), .C(n12207), .D(n12208), .Y(n12159)
         );
  NOR4X1 U12640 ( .A(n12209), .B(n12210), .C(n12211), .D(n12212), .Y(n12208)
         );
  NOR2X1 U12641 ( .A(n10664), .B(n11913), .Y(n12212) );
  NOR2X1 U12642 ( .A(n10663), .B(n11914), .Y(n12211) );
  NAND2X1 U12643 ( .A(n12213), .B(n12214), .Y(n12210) );
  NAND2X1 U12644 ( .A(n11917), .B(G21537), .Y(n12214) );
  NAND2X1 U12645 ( .A(n11918), .B(G21545), .Y(n12213) );
  NOR2X1 U12646 ( .A(n10657), .B(n11919), .Y(n12209) );
  NOR4X1 U12647 ( .A(n12215), .B(n12216), .C(n12217), .D(n12218), .Y(n12207)
         );
  NOR2X1 U12648 ( .A(n10665), .B(n11924), .Y(n12218) );
  NOR2X1 U12649 ( .A(n10639), .B(n11925), .Y(n12217) );
  NOR2X1 U12650 ( .A(n10640), .B(n11926), .Y(n12216) );
  NOR2X1 U12651 ( .A(n10641), .B(n11927), .Y(n12215) );
  NOR4X1 U12652 ( .A(n12219), .B(n12220), .C(n12221), .D(n12222), .Y(n12206)
         );
  NOR2X1 U12653 ( .A(n10647), .B(n11932), .Y(n12222) );
  NOR2X1 U12654 ( .A(n10648), .B(n11933), .Y(n12221) );
  NOR2X1 U12655 ( .A(n10649), .B(n11934), .Y(n12220) );
  NOR2X1 U12656 ( .A(n10654), .B(n11935), .Y(n12219) );
  NOR4X1 U12657 ( .A(n12223), .B(n12224), .C(n12225), .D(n9908), .Y(n12205) );
  NOR2X1 U12658 ( .A(n10638), .B(n11939), .Y(n12225) );
  NOR2X1 U12659 ( .A(n10646), .B(n11940), .Y(n12224) );
  NOR2X1 U12660 ( .A(n10662), .B(n11941), .Y(n12223) );
  NAND2X1 U12661 ( .A(n12011), .B(n12226), .Y(n12158) );
  NAND4X1 U12662 ( .A(n12227), .B(n12228), .C(n12229), .D(n12230), .Y(n12226)
         );
  NOR4X1 U12663 ( .A(n12231), .B(n12232), .C(n12233), .D(n12234), .Y(n12230)
         );
  NOR2X1 U12664 ( .A(n10639), .B(n8688), .Y(n12234) );
  NOR2X1 U12665 ( .A(n10640), .B(n8610), .Y(n12233) );
  NOR2X1 U12666 ( .A(n10641), .B(n8528), .Y(n12232) );
  NOR2X1 U12667 ( .A(n10647), .B(n8371), .Y(n12231) );
  NOR4X1 U12668 ( .A(n12235), .B(n12236), .C(n12237), .D(n12238), .Y(n12229)
         );
  NOR2X1 U12669 ( .A(n10648), .B(n8293), .Y(n12238) );
  NOR2X1 U12670 ( .A(n10649), .B(n8213), .Y(n12237) );
  NOR2X1 U12671 ( .A(n10664), .B(n8056), .Y(n12236) );
  NOR2X1 U12672 ( .A(n10663), .B(n7978), .Y(n12235) );
  NOR4X1 U12673 ( .A(n12239), .B(n12240), .C(n12241), .D(n12242), .Y(n12228)
         );
  NOR2X1 U12674 ( .A(n10662), .B(n7898), .Y(n12242) );
  NOR2X1 U12675 ( .A(n10656), .B(n7736), .Y(n12241) );
  NOR2X1 U12676 ( .A(n10655), .B(n7656), .Y(n12240) );
  NOR2X1 U12677 ( .A(n10654), .B(n7570), .Y(n12239) );
  NOR4X1 U12678 ( .A(n12243), .B(n12244), .C(n12245), .D(n12246), .Y(n12227)
         );
  NOR2X1 U12679 ( .A(n10638), .B(n8803), .Y(n12246) );
  NOR2X1 U12680 ( .A(n10646), .B(n8449), .Y(n12245) );
  NOR2X1 U12681 ( .A(n10665), .B(n8134), .Y(n12244) );
  NOR2X1 U12682 ( .A(n10657), .B(n7816), .Y(n12243) );
  OR2X1 U12683 ( .A(n12247), .B(n12248), .Y(n9968) );
  NAND2X1 U12684 ( .A(n12248), .B(n12247), .Y(n9967) );
  NAND4X1 U12685 ( .A(n12249), .B(n12250), .C(n12251), .D(n12252), .Y(n12247)
         );
  NAND2X1 U12686 ( .A(n6961), .B(n11800), .Y(n12252) );
  ADDHXL U12687 ( .A(n12253), .B(n12254), .S(n6961) );
  AND2X1 U12688 ( .A(n12255), .B(n12256), .Y(n12254) );
  NAND2X1 U12689 ( .A(n11705), .B(G21762), .Y(n12251) );
  NAND2X1 U12690 ( .A(G21571), .B(n10444), .Y(n12250) );
  NAND2X1 U12691 ( .A(n9926), .B(n6959), .Y(n12249) );
  ADDHXL U12692 ( .A(n9926), .B(n12257), .S(n12248) );
  NAND4X1 U12693 ( .A(n12258), .B(n12259), .C(n12260), .D(n12261), .Y(n12257)
         );
  NOR2X1 U12694 ( .A(n12262), .B(n12263), .Y(n12261) );
  NOR2X1 U12695 ( .A(n7439), .B(n8848), .Y(n12263) );
  NOR2X1 U12696 ( .A(n12264), .B(n9192), .Y(n12262) );
  NOR4X1 U12697 ( .A(n12265), .B(n12266), .C(n12267), .D(n12268), .Y(n12264)
         );
  NAND4X1 U12698 ( .A(n12269), .B(n12270), .C(n12271), .D(n12272), .Y(n12268)
         );
  NAND2X1 U12699 ( .A(n11959), .B(G21552), .Y(n12272) );
  INVX1 U12700 ( .A(n11904), .Y(n11959) );
  NAND2X1 U12701 ( .A(n11960), .B(G21544), .Y(n12271) );
  INVX1 U12702 ( .A(n11903), .Y(n11960) );
  NAND2X1 U12703 ( .A(n11961), .B(G21536), .Y(n12270) );
  INVX1 U12704 ( .A(n11902), .Y(n11961) );
  NAND2X1 U12705 ( .A(n11962), .B(G21528), .Y(n12269) );
  INVX1 U12706 ( .A(n11901), .Y(n11962) );
  NAND4X1 U12707 ( .A(n12273), .B(n12274), .C(n12275), .D(n12276), .Y(n12267)
         );
  NAND2X1 U12708 ( .A(n11967), .B(G21520), .Y(n12276) );
  INVX1 U12709 ( .A(n11896), .Y(n11967) );
  NAND2X1 U12710 ( .A(n11968), .B(G21512), .Y(n12275) );
  INVX1 U12711 ( .A(n11895), .Y(n11968) );
  NAND2X1 U12712 ( .A(n11969), .B(G21504), .Y(n12274) );
  INVX1 U12713 ( .A(n11894), .Y(n11969) );
  NAND2X1 U12714 ( .A(n11970), .B(G21496), .Y(n12273) );
  INVX1 U12715 ( .A(n11893), .Y(n11970) );
  NAND4X1 U12716 ( .A(n12277), .B(n12278), .C(n12279), .D(n12280), .Y(n12266)
         );
  NAND2X1 U12717 ( .A(n11975), .B(G21488), .Y(n12280) );
  INVX1 U12718 ( .A(n11888), .Y(n11975) );
  NAND2X1 U12719 ( .A(n11976), .B(G21480), .Y(n12279) );
  INVX1 U12720 ( .A(n11887), .Y(n11976) );
  NAND2X1 U12721 ( .A(n11977), .B(G21472), .Y(n12278) );
  INVX1 U12722 ( .A(n11886), .Y(n11977) );
  NAND2X1 U12723 ( .A(n11978), .B(G21464), .Y(n12277) );
  INVX1 U12724 ( .A(n11885), .Y(n11978) );
  NAND4X1 U12725 ( .A(n12281), .B(n12282), .C(n12283), .D(n12284), .Y(n12265)
         );
  NAND2X1 U12726 ( .A(n11983), .B(G21456), .Y(n12284) );
  INVX1 U12727 ( .A(n11880), .Y(n11983) );
  NAND2X1 U12728 ( .A(n11984), .B(G21448), .Y(n12283) );
  INVX1 U12729 ( .A(n11879), .Y(n11984) );
  NAND2X1 U12730 ( .A(n11985), .B(G21440), .Y(n12282) );
  INVX1 U12731 ( .A(n11878), .Y(n11985) );
  NAND2X1 U12732 ( .A(n11986), .B(G21432), .Y(n12281) );
  INVX1 U12733 ( .A(n11877), .Y(n11986) );
  NAND2X1 U12734 ( .A(n11809), .B(n11122), .Y(n12260) );
  NAND4X1 U12735 ( .A(n12285), .B(n12286), .C(n12287), .D(n12288), .Y(n11122)
         );
  NOR4X1 U12736 ( .A(n12289), .B(n12290), .C(n12291), .D(n12292), .Y(n12288)
         );
  NOR2X1 U12737 ( .A(n10557), .B(n11818), .Y(n12292) );
  NOR2X1 U12738 ( .A(n10558), .B(n11819), .Y(n12291) );
  NOR2X1 U12739 ( .A(n10559), .B(n11820), .Y(n12290) );
  NOR2X1 U12740 ( .A(n10565), .B(n11821), .Y(n12289) );
  NOR4X1 U12741 ( .A(n12293), .B(n12294), .C(n12295), .D(n12296), .Y(n12287)
         );
  NOR2X1 U12742 ( .A(n10566), .B(n11826), .Y(n12296) );
  NOR2X1 U12743 ( .A(n10567), .B(n11827), .Y(n12295) );
  NOR2X1 U12744 ( .A(n10582), .B(n11828), .Y(n12294) );
  NOR2X1 U12745 ( .A(n10581), .B(n11829), .Y(n12293) );
  NOR4X1 U12746 ( .A(n12297), .B(n12298), .C(n12299), .D(n12300), .Y(n12286)
         );
  NOR2X1 U12747 ( .A(n10580), .B(n11834), .Y(n12300) );
  NOR2X1 U12748 ( .A(n10574), .B(n11835), .Y(n12299) );
  NOR2X1 U12749 ( .A(n10573), .B(n11836), .Y(n12298) );
  NOR2X1 U12750 ( .A(n10572), .B(n11837), .Y(n12297) );
  NOR4X1 U12751 ( .A(n12301), .B(n12302), .C(n12303), .D(n12304), .Y(n12285)
         );
  NOR2X1 U12752 ( .A(n10556), .B(n11842), .Y(n12304) );
  NOR2X1 U12753 ( .A(n10564), .B(n11843), .Y(n12303) );
  NOR2X1 U12754 ( .A(n10583), .B(n11844), .Y(n12302) );
  NOR2X1 U12755 ( .A(n10575), .B(n11845), .Y(n12301) );
  NAND4X1 U12756 ( .A(n12305), .B(n12306), .C(n12307), .D(n12308), .Y(n12259)
         );
  NOR4X1 U12757 ( .A(n12309), .B(n12310), .C(n12311), .D(n12312), .Y(n12308)
         );
  NOR2X1 U12758 ( .A(n10582), .B(n11913), .Y(n12312) );
  NOR2X1 U12759 ( .A(n10581), .B(n11914), .Y(n12311) );
  NAND2X1 U12760 ( .A(n12313), .B(n12314), .Y(n12310) );
  NAND2X1 U12761 ( .A(n11917), .B(G21536), .Y(n12314) );
  NAND2X1 U12762 ( .A(n11918), .B(G21544), .Y(n12313) );
  NOR2X1 U12763 ( .A(n10575), .B(n11919), .Y(n12309) );
  NOR4X1 U12764 ( .A(n12315), .B(n12316), .C(n12317), .D(n12318), .Y(n12307)
         );
  NOR2X1 U12765 ( .A(n10583), .B(n11924), .Y(n12318) );
  NOR2X1 U12766 ( .A(n10557), .B(n11925), .Y(n12317) );
  NOR2X1 U12767 ( .A(n10558), .B(n11926), .Y(n12316) );
  NOR2X1 U12768 ( .A(n10559), .B(n11927), .Y(n12315) );
  NOR4X1 U12769 ( .A(n12319), .B(n12320), .C(n12321), .D(n12322), .Y(n12306)
         );
  NOR2X1 U12770 ( .A(n10565), .B(n11932), .Y(n12322) );
  NOR2X1 U12771 ( .A(n10566), .B(n11933), .Y(n12321) );
  NOR2X1 U12772 ( .A(n10567), .B(n11934), .Y(n12320) );
  NOR2X1 U12773 ( .A(n10572), .B(n11935), .Y(n12319) );
  NOR4X1 U12774 ( .A(n12323), .B(n12324), .C(n12325), .D(n9908), .Y(n12305) );
  NOR2X1 U12775 ( .A(n10556), .B(n11939), .Y(n12325) );
  NOR2X1 U12776 ( .A(n10564), .B(n11940), .Y(n12324) );
  NOR2X1 U12777 ( .A(n10580), .B(n11941), .Y(n12323) );
  NAND2X1 U12778 ( .A(n12011), .B(n12326), .Y(n12258) );
  NAND4X1 U12779 ( .A(n12327), .B(n12328), .C(n12329), .D(n12330), .Y(n12326)
         );
  NOR4X1 U12780 ( .A(n12331), .B(n12332), .C(n12333), .D(n12334), .Y(n12330)
         );
  NOR2X1 U12781 ( .A(n10557), .B(n8688), .Y(n12334) );
  NOR2X1 U12782 ( .A(n10558), .B(n8610), .Y(n12333) );
  NOR2X1 U12783 ( .A(n10559), .B(n8528), .Y(n12332) );
  NOR2X1 U12784 ( .A(n10565), .B(n8371), .Y(n12331) );
  NOR4X1 U12785 ( .A(n12335), .B(n12336), .C(n12337), .D(n12338), .Y(n12329)
         );
  NOR2X1 U12786 ( .A(n10566), .B(n8293), .Y(n12338) );
  NOR2X1 U12787 ( .A(n10567), .B(n8213), .Y(n12337) );
  NOR2X1 U12788 ( .A(n10582), .B(n8056), .Y(n12336) );
  NOR2X1 U12789 ( .A(n10581), .B(n7978), .Y(n12335) );
  NOR4X1 U12790 ( .A(n12339), .B(n12340), .C(n12341), .D(n12342), .Y(n12328)
         );
  NOR2X1 U12791 ( .A(n10580), .B(n7898), .Y(n12342) );
  NOR2X1 U12792 ( .A(n10574), .B(n7736), .Y(n12341) );
  NOR2X1 U12793 ( .A(n10573), .B(n7656), .Y(n12340) );
  NOR2X1 U12794 ( .A(n10572), .B(n7570), .Y(n12339) );
  NOR4X1 U12795 ( .A(n12343), .B(n12344), .C(n12345), .D(n12346), .Y(n12327)
         );
  NOR2X1 U12796 ( .A(n10556), .B(n8803), .Y(n12346) );
  NOR2X1 U12797 ( .A(n10564), .B(n8449), .Y(n12345) );
  NOR2X1 U12798 ( .A(n10583), .B(n8134), .Y(n12344) );
  NOR2X1 U12799 ( .A(n10575), .B(n7816), .Y(n12343) );
  OR2X1 U12800 ( .A(n11779), .B(n11778), .Y(n9960) );
  ADDHXL U12801 ( .A(n12347), .B(n9926), .S(n11778) );
  NAND4X1 U12802 ( .A(n12348), .B(n12349), .C(n12350), .D(n12351), .Y(n12347)
         );
  NAND4X1 U12803 ( .A(n12352), .B(n12353), .C(n12354), .D(n12355), .Y(n12351)
         );
  NOR4X1 U12804 ( .A(n12356), .B(n12357), .C(n12358), .D(n12359), .Y(n12355)
         );
  NOR2X1 U12805 ( .A(n11105), .B(n11913), .Y(n12359) );
  NOR2X1 U12806 ( .A(n11100), .B(n11914), .Y(n12358) );
  NAND2X1 U12807 ( .A(n12360), .B(n12361), .Y(n12357) );
  NAND2X1 U12808 ( .A(n11917), .B(G21535), .Y(n12361) );
  NAND2X1 U12809 ( .A(n11918), .B(G21543), .Y(n12360) );
  NOR2X1 U12810 ( .A(n11099), .B(n11919), .Y(n12356) );
  NOR4X1 U12811 ( .A(n12362), .B(n12363), .C(n12364), .D(n12365), .Y(n12354)
         );
  NOR2X1 U12812 ( .A(n11106), .B(n11924), .Y(n12365) );
  NOR2X1 U12813 ( .A(n10492), .B(n11925), .Y(n12364) );
  NOR2X1 U12814 ( .A(n10493), .B(n11926), .Y(n12363) );
  NOR2X1 U12815 ( .A(n10494), .B(n11927), .Y(n12362) );
  NOR4X1 U12816 ( .A(n12366), .B(n12367), .C(n12368), .D(n12369), .Y(n12353)
         );
  NOR2X1 U12817 ( .A(n10500), .B(n11932), .Y(n12369) );
  NOR2X1 U12818 ( .A(n10501), .B(n11933), .Y(n12368) );
  NOR2X1 U12819 ( .A(n10502), .B(n11934), .Y(n12367) );
  NOR2X1 U12820 ( .A(n11115), .B(n11935), .Y(n12366) );
  NOR4X1 U12821 ( .A(n12370), .B(n12371), .C(n12372), .D(n9908), .Y(n12352) );
  NOR2X1 U12822 ( .A(n10491), .B(n11939), .Y(n12372) );
  NOR2X1 U12823 ( .A(n10499), .B(n11940), .Y(n12371) );
  NOR2X1 U12824 ( .A(n11116), .B(n11941), .Y(n12370) );
  NAND2X1 U12825 ( .A(n11809), .B(n11072), .Y(n12350) );
  NAND4X1 U12826 ( .A(n12373), .B(n12374), .C(n12375), .D(n12376), .Y(n11072)
         );
  NOR4X1 U12827 ( .A(n12377), .B(n12378), .C(n12379), .D(n12380), .Y(n12376)
         );
  NOR2X1 U12828 ( .A(n10492), .B(n11818), .Y(n12380) );
  NOR2X1 U12829 ( .A(n10493), .B(n11819), .Y(n12379) );
  NOR2X1 U12830 ( .A(n10494), .B(n11820), .Y(n12378) );
  NOR2X1 U12831 ( .A(n10500), .B(n11821), .Y(n12377) );
  NOR4X1 U12832 ( .A(n12381), .B(n12382), .C(n12383), .D(n12384), .Y(n12375)
         );
  NOR2X1 U12833 ( .A(n10501), .B(n11826), .Y(n12384) );
  NOR2X1 U12834 ( .A(n10502), .B(n11827), .Y(n12383) );
  NOR2X1 U12835 ( .A(n11105), .B(n11828), .Y(n12382) );
  NOR2X1 U12836 ( .A(n11100), .B(n11829), .Y(n12381) );
  NOR4X1 U12837 ( .A(n12385), .B(n12386), .C(n12387), .D(n12388), .Y(n12374)
         );
  NOR2X1 U12838 ( .A(n11116), .B(n11834), .Y(n12388) );
  NOR2X1 U12839 ( .A(n11098), .B(n11835), .Y(n12387) );
  NOR2X1 U12840 ( .A(n11097), .B(n11836), .Y(n12386) );
  NOR2X1 U12841 ( .A(n11115), .B(n11837), .Y(n12385) );
  NOR4X1 U12842 ( .A(n12389), .B(n12390), .C(n12391), .D(n12392), .Y(n12373)
         );
  NOR2X1 U12843 ( .A(n10491), .B(n11842), .Y(n12392) );
  NOR2X1 U12844 ( .A(n10499), .B(n11843), .Y(n12391) );
  NOR2X1 U12845 ( .A(n11106), .B(n11844), .Y(n12390) );
  NOR2X1 U12846 ( .A(n11099), .B(n11845), .Y(n12389) );
  NAND2X1 U12847 ( .A(n10256), .B(n12393), .Y(n12349) );
  NAND4X1 U12848 ( .A(n12394), .B(n12395), .C(n12396), .D(n12397), .Y(n12393)
         );
  NOR4X1 U12849 ( .A(n12398), .B(n12399), .C(n12400), .D(n12401), .Y(n12397)
         );
  NOR2X1 U12850 ( .A(n10491), .B(n11877), .Y(n12401) );
  NOR2X1 U12851 ( .A(n10492), .B(n11878), .Y(n12400) );
  NOR2X1 U12852 ( .A(n10493), .B(n11879), .Y(n12399) );
  NOR2X1 U12853 ( .A(n10494), .B(n11880), .Y(n12398) );
  NOR4X1 U12854 ( .A(n12402), .B(n12403), .C(n12404), .D(n12405), .Y(n12396)
         );
  NOR2X1 U12855 ( .A(n10499), .B(n11885), .Y(n12405) );
  NOR2X1 U12856 ( .A(n10500), .B(n11886), .Y(n12404) );
  NOR2X1 U12857 ( .A(n10501), .B(n11887), .Y(n12403) );
  NOR2X1 U12858 ( .A(n10502), .B(n11888), .Y(n12402) );
  NOR4X1 U12859 ( .A(n12406), .B(n12407), .C(n12408), .D(n12409), .Y(n12395)
         );
  NOR2X1 U12860 ( .A(n11106), .B(n11893), .Y(n12409) );
  NOR2X1 U12861 ( .A(n11105), .B(n11894), .Y(n12408) );
  NOR2X1 U12862 ( .A(n11100), .B(n11895), .Y(n12407) );
  NOR2X1 U12863 ( .A(n11116), .B(n11896), .Y(n12406) );
  NOR4X1 U12864 ( .A(n12410), .B(n12411), .C(n12412), .D(n12413), .Y(n12394)
         );
  NOR2X1 U12865 ( .A(n11099), .B(n11901), .Y(n12413) );
  NOR2X1 U12866 ( .A(n11098), .B(n11902), .Y(n12412) );
  NOR2X1 U12867 ( .A(n11097), .B(n11903), .Y(n12411) );
  NOR2X1 U12868 ( .A(n11115), .B(n11904), .Y(n12410) );
  NAND2X1 U12869 ( .A(n12011), .B(n12414), .Y(n12348) );
  NAND4X1 U12870 ( .A(n12415), .B(n12416), .C(n12417), .D(n12418), .Y(n12414)
         );
  NOR4X1 U12871 ( .A(n12419), .B(n12420), .C(n12421), .D(n12422), .Y(n12418)
         );
  NOR2X1 U12872 ( .A(n10492), .B(n8688), .Y(n12422) );
  NOR2X1 U12873 ( .A(n10493), .B(n8610), .Y(n12421) );
  NOR2X1 U12874 ( .A(n10494), .B(n8528), .Y(n12420) );
  NOR2X1 U12875 ( .A(n10500), .B(n8371), .Y(n12419) );
  NOR4X1 U12876 ( .A(n12423), .B(n12424), .C(n12425), .D(n12426), .Y(n12417)
         );
  NOR2X1 U12877 ( .A(n10501), .B(n8293), .Y(n12426) );
  NOR2X1 U12878 ( .A(n10502), .B(n8213), .Y(n12425) );
  NOR2X1 U12879 ( .A(n11105), .B(n8056), .Y(n12424) );
  NOR2X1 U12880 ( .A(n11100), .B(n7978), .Y(n12423) );
  NOR4X1 U12881 ( .A(n12427), .B(n12428), .C(n12429), .D(n12430), .Y(n12416)
         );
  NOR2X1 U12882 ( .A(n11116), .B(n7898), .Y(n12430) );
  NOR2X1 U12883 ( .A(n11098), .B(n7736), .Y(n12429) );
  NOR2X1 U12884 ( .A(n11097), .B(n7656), .Y(n12428) );
  NOR2X1 U12885 ( .A(n11115), .B(n7570), .Y(n12427) );
  NOR4X1 U12886 ( .A(n12431), .B(n12432), .C(n12433), .D(n12434), .Y(n12415)
         );
  NOR2X1 U12887 ( .A(n10491), .B(n8803), .Y(n12434) );
  NOR2X1 U12888 ( .A(n10499), .B(n8449), .Y(n12433) );
  NOR2X1 U12889 ( .A(n11106), .B(n8134), .Y(n12432) );
  NOR2X1 U12890 ( .A(n11099), .B(n7816), .Y(n12431) );
  NAND4X1 U12891 ( .A(n12435), .B(n12436), .C(n12437), .D(n12438), .Y(n11779)
         );
  NAND2X1 U12892 ( .A(n6950), .B(n11800), .Y(n12438) );
  ADDHXL U12893 ( .A(n12439), .B(n12440), .S(n6950) );
  AND2X1 U12894 ( .A(n12441), .B(n12442), .Y(n12440) );
  NAND2X1 U12895 ( .A(n11705), .B(G21763), .Y(n12437) );
  NAND2X1 U12896 ( .A(G21572), .B(n10444), .Y(n12436) );
  NAND2X1 U12897 ( .A(n9926), .B(n6948), .Y(n12435) );
  NAND2X1 U12898 ( .A(n12443), .B(n12444), .Y(n9953) );
  ADDHXL U12899 ( .A(n9908), .B(n11776), .S(n12444) );
  NAND4X1 U12900 ( .A(n12445), .B(n12446), .C(n12447), .D(n12448), .Y(n11776)
         );
  NAND4X1 U12901 ( .A(n12449), .B(n12450), .C(n12451), .D(n12452), .Y(n12448)
         );
  NOR4X1 U12902 ( .A(n12453), .B(n12454), .C(n12455), .D(n12456), .Y(n12452)
         );
  NOR2X1 U12903 ( .A(n10421), .B(n11913), .Y(n12456) );
  NOR2X1 U12904 ( .A(n10419), .B(n11914), .Y(n12455) );
  NAND2X1 U12905 ( .A(n12457), .B(n12458), .Y(n12454) );
  NAND2X1 U12906 ( .A(n11917), .B(G21534), .Y(n12458) );
  NAND2X1 U12907 ( .A(n11918), .B(G21542), .Y(n12457) );
  NOR2X1 U12908 ( .A(n10411), .B(n11919), .Y(n12453) );
  NOR4X1 U12909 ( .A(n12459), .B(n12460), .C(n12461), .D(n12462), .Y(n12451)
         );
  NOR2X1 U12910 ( .A(n10423), .B(n11924), .Y(n12462) );
  NOR2X1 U12911 ( .A(n10390), .B(n11925), .Y(n12461) );
  NOR2X1 U12912 ( .A(n10391), .B(n11926), .Y(n12460) );
  NOR2X1 U12913 ( .A(n10392), .B(n11927), .Y(n12459) );
  NOR4X1 U12914 ( .A(n12463), .B(n12464), .C(n12465), .D(n12466), .Y(n12450)
         );
  NOR2X1 U12915 ( .A(n10398), .B(n11932), .Y(n12466) );
  NOR2X1 U12916 ( .A(n10399), .B(n11933), .Y(n12465) );
  NOR2X1 U12917 ( .A(n10400), .B(n11934), .Y(n12464) );
  NOR2X1 U12918 ( .A(n10405), .B(n11935), .Y(n12463) );
  NOR4X1 U12919 ( .A(n12467), .B(n12468), .C(n12469), .D(n9908), .Y(n12449) );
  NOR2X1 U12920 ( .A(n10389), .B(n11939), .Y(n12469) );
  NOR2X1 U12921 ( .A(n10397), .B(n11940), .Y(n12468) );
  NOR2X1 U12922 ( .A(n10417), .B(n11941), .Y(n12467) );
  NAND2X1 U12923 ( .A(n11809), .B(n10871), .Y(n12447) );
  NAND4X1 U12924 ( .A(n12470), .B(n12471), .C(n12472), .D(n12473), .Y(n10871)
         );
  NOR4X1 U12925 ( .A(n12474), .B(n12475), .C(n12476), .D(n12477), .Y(n12473)
         );
  NOR2X1 U12926 ( .A(n10390), .B(n11818), .Y(n12477) );
  NOR2X1 U12927 ( .A(n10391), .B(n11819), .Y(n12476) );
  NOR2X1 U12928 ( .A(n10392), .B(n11820), .Y(n12475) );
  NOR2X1 U12929 ( .A(n10398), .B(n11821), .Y(n12474) );
  NOR4X1 U12930 ( .A(n12478), .B(n12479), .C(n12480), .D(n12481), .Y(n12472)
         );
  NOR2X1 U12931 ( .A(n10399), .B(n11826), .Y(n12481) );
  NOR2X1 U12932 ( .A(n10400), .B(n11827), .Y(n12480) );
  NOR2X1 U12933 ( .A(n10421), .B(n11828), .Y(n12479) );
  NOR2X1 U12934 ( .A(n10419), .B(n11829), .Y(n12478) );
  NOR4X1 U12935 ( .A(n12482), .B(n12483), .C(n12484), .D(n12485), .Y(n12471)
         );
  NOR2X1 U12936 ( .A(n10417), .B(n11834), .Y(n12485) );
  NOR2X1 U12937 ( .A(n10409), .B(n11835), .Y(n12484) );
  NOR2X1 U12938 ( .A(n10407), .B(n11836), .Y(n12483) );
  NOR2X1 U12939 ( .A(n10405), .B(n11837), .Y(n12482) );
  NOR4X1 U12940 ( .A(n12486), .B(n12487), .C(n12488), .D(n12489), .Y(n12470)
         );
  NOR2X1 U12941 ( .A(n10389), .B(n11842), .Y(n12489) );
  NOR2X1 U12942 ( .A(n10397), .B(n11843), .Y(n12488) );
  NOR2X1 U12943 ( .A(n10423), .B(n11844), .Y(n12487) );
  NOR2X1 U12944 ( .A(n10411), .B(n11845), .Y(n12486) );
  NAND2X1 U12945 ( .A(n10256), .B(n12490), .Y(n12446) );
  NAND4X1 U12946 ( .A(n12491), .B(n12492), .C(n12493), .D(n12494), .Y(n12490)
         );
  NOR4X1 U12947 ( .A(n12495), .B(n12496), .C(n12497), .D(n12498), .Y(n12494)
         );
  NOR2X1 U12948 ( .A(n10389), .B(n11877), .Y(n12498) );
  NOR2X1 U12949 ( .A(n10390), .B(n11878), .Y(n12497) );
  NOR2X1 U12950 ( .A(n10391), .B(n11879), .Y(n12496) );
  NOR2X1 U12951 ( .A(n10392), .B(n11880), .Y(n12495) );
  NOR4X1 U12952 ( .A(n12499), .B(n12500), .C(n12501), .D(n12502), .Y(n12493)
         );
  NOR2X1 U12953 ( .A(n10397), .B(n11885), .Y(n12502) );
  NOR2X1 U12954 ( .A(n10398), .B(n11886), .Y(n12501) );
  NOR2X1 U12955 ( .A(n10399), .B(n11887), .Y(n12500) );
  NOR2X1 U12956 ( .A(n10400), .B(n11888), .Y(n12499) );
  NOR4X1 U12957 ( .A(n12503), .B(n12504), .C(n12505), .D(n12506), .Y(n12492)
         );
  NOR2X1 U12958 ( .A(n10423), .B(n11893), .Y(n12506) );
  NOR2X1 U12959 ( .A(n10421), .B(n11894), .Y(n12505) );
  NOR2X1 U12960 ( .A(n10419), .B(n11895), .Y(n12504) );
  NOR2X1 U12961 ( .A(n10417), .B(n11896), .Y(n12503) );
  NOR4X1 U12962 ( .A(n12507), .B(n12508), .C(n12509), .D(n12510), .Y(n12491)
         );
  NOR2X1 U12963 ( .A(n10411), .B(n11901), .Y(n12510) );
  NOR2X1 U12964 ( .A(n10409), .B(n11902), .Y(n12509) );
  NOR2X1 U12965 ( .A(n10407), .B(n11903), .Y(n12508) );
  NOR2X1 U12966 ( .A(n10405), .B(n11904), .Y(n12507) );
  NAND2X1 U12967 ( .A(n12011), .B(n12511), .Y(n12445) );
  NAND4X1 U12968 ( .A(n12512), .B(n12513), .C(n12514), .D(n12515), .Y(n12511)
         );
  NOR4X1 U12969 ( .A(n12516), .B(n12517), .C(n12518), .D(n12519), .Y(n12515)
         );
  NOR2X1 U12970 ( .A(n10390), .B(n8688), .Y(n12519) );
  NOR2X1 U12971 ( .A(n10391), .B(n8610), .Y(n12518) );
  NOR2X1 U12972 ( .A(n10392), .B(n8528), .Y(n12517) );
  NOR2X1 U12973 ( .A(n10398), .B(n8371), .Y(n12516) );
  NOR4X1 U12974 ( .A(n12520), .B(n12521), .C(n12522), .D(n12523), .Y(n12514)
         );
  NOR2X1 U12975 ( .A(n10399), .B(n8293), .Y(n12523) );
  NOR2X1 U12976 ( .A(n10400), .B(n8213), .Y(n12522) );
  NOR2X1 U12977 ( .A(n10421), .B(n8056), .Y(n12521) );
  NOR2X1 U12978 ( .A(n10419), .B(n7978), .Y(n12520) );
  NOR4X1 U12979 ( .A(n12524), .B(n12525), .C(n12526), .D(n12527), .Y(n12513)
         );
  NOR2X1 U12980 ( .A(n10417), .B(n7898), .Y(n12527) );
  NOR2X1 U12981 ( .A(n10409), .B(n7736), .Y(n12526) );
  NOR2X1 U12982 ( .A(n10407), .B(n7656), .Y(n12525) );
  NOR2X1 U12983 ( .A(n10405), .B(n7570), .Y(n12524) );
  NOR4X1 U12984 ( .A(n12528), .B(n12529), .C(n12530), .D(n12531), .Y(n12512)
         );
  NOR2X1 U12985 ( .A(n10389), .B(n8803), .Y(n12531) );
  NOR2X1 U12986 ( .A(n10397), .B(n8449), .Y(n12530) );
  NOR2X1 U12987 ( .A(n10423), .B(n8134), .Y(n12529) );
  NOR2X1 U12988 ( .A(n10411), .B(n7816), .Y(n12528) );
  INVX1 U12989 ( .A(n11775), .Y(n12443) );
  NAND4X1 U12990 ( .A(n12532), .B(n12533), .C(n12534), .D(n12535), .Y(n11775)
         );
  NAND2X1 U12991 ( .A(n6939), .B(n11800), .Y(n12535) );
  INVX1 U12992 ( .A(n9570), .Y(n6939) );
  NAND2X1 U12993 ( .A(n12536), .B(n12537), .Y(n9570) );
  NAND2X1 U12994 ( .A(n12538), .B(n12539), .Y(n12537) );
  INVX1 U12995 ( .A(n12540), .Y(n12538) );
  NAND3X1 U12996 ( .A(n12541), .B(n12441), .C(n12542), .Y(n12536) );
  NAND2X1 U12997 ( .A(n12539), .B(n12543), .Y(n12541) );
  NAND2X1 U12998 ( .A(n11705), .B(G21764), .Y(n12534) );
  NAND2X1 U12999 ( .A(G21573), .B(n10444), .Y(n12533) );
  NAND2X1 U13000 ( .A(n9926), .B(n6937), .Y(n12532) );
  NAND2X1 U13001 ( .A(n11773), .B(n11772), .Y(n9939) );
  NAND4X1 U13002 ( .A(n12544), .B(n12545), .C(n12546), .D(n12547), .Y(n11772)
         );
  NAND2X1 U13003 ( .A(n6928), .B(n11800), .Y(n12547) );
  NAND2X1 U13004 ( .A(n10217), .B(n9192), .Y(n11800) );
  ADDHXL U13005 ( .A(n12548), .B(n12549), .S(n6928) );
  AND2X1 U13006 ( .A(n12550), .B(n12551), .Y(n12549) );
  NAND2X1 U13007 ( .A(n11705), .B(G21765), .Y(n12546) );
  NAND2X1 U13008 ( .A(G21574), .B(n10444), .Y(n12545) );
  NAND2X1 U13009 ( .A(n9926), .B(n6926), .Y(n12544) );
  ADDHXL U13010 ( .A(n9926), .B(n12552), .S(n11773) );
  NAND4X1 U13011 ( .A(n12553), .B(n12554), .C(n12555), .D(n12556), .Y(n12552)
         );
  NAND4X1 U13012 ( .A(n12557), .B(n12558), .C(n12559), .D(n12560), .Y(n12556)
         );
  NOR4X1 U13013 ( .A(n12561), .B(n12562), .C(n12563), .D(n12564), .Y(n12560)
         );
  NOR2X1 U13014 ( .A(n10972), .B(n11913), .Y(n12564) );
  NAND2X1 U13015 ( .A(n12565), .B(n12566), .Y(n11913) );
  NOR2X1 U13016 ( .A(n10967), .B(n11914), .Y(n12563) );
  NAND2X1 U13017 ( .A(n12565), .B(n12567), .Y(n11914) );
  NAND2X1 U13018 ( .A(n12568), .B(n12569), .Y(n12562) );
  NAND2X1 U13019 ( .A(n11917), .B(G21533), .Y(n12569) );
  INVX1 U13020 ( .A(n12010), .Y(n11917) );
  NAND2X1 U13021 ( .A(n12566), .B(n12570), .Y(n12010) );
  NAND2X1 U13022 ( .A(n11918), .B(G21541), .Y(n12568) );
  INVX1 U13023 ( .A(n12009), .Y(n11918) );
  NAND2X1 U13024 ( .A(n12567), .B(n12570), .Y(n12009) );
  NOR2X1 U13025 ( .A(n10966), .B(n11919), .Y(n12561) );
  NAND2X1 U13026 ( .A(n12571), .B(n12570), .Y(n11919) );
  NOR4X1 U13027 ( .A(n12572), .B(n12573), .C(n12574), .D(n12575), .Y(n12559)
         );
  NOR2X1 U13028 ( .A(n10973), .B(n11924), .Y(n12575) );
  NAND2X1 U13029 ( .A(n12565), .B(n12571), .Y(n11924) );
  NOR2X1 U13030 ( .A(n10312), .B(n11925), .Y(n12574) );
  NAND2X1 U13031 ( .A(n12576), .B(n12566), .Y(n11925) );
  NOR2X1 U13032 ( .A(n10314), .B(n11926), .Y(n12573) );
  NAND2X1 U13033 ( .A(n12576), .B(n12567), .Y(n11926) );
  NOR2X1 U13034 ( .A(n10316), .B(n11927), .Y(n12572) );
  NAND2X1 U13035 ( .A(n12576), .B(n12577), .Y(n11927) );
  NOR4X1 U13036 ( .A(n12578), .B(n12579), .C(n12580), .D(n12581), .Y(n12558)
         );
  NOR2X1 U13037 ( .A(n10324), .B(n11932), .Y(n12581) );
  NAND2X1 U13038 ( .A(n12582), .B(n12566), .Y(n11932) );
  NOR2X1 U13039 ( .A(n7003), .B(n9615), .Y(n12566) );
  NOR2X1 U13040 ( .A(n10326), .B(n11933), .Y(n12580) );
  NAND2X1 U13041 ( .A(n12582), .B(n12567), .Y(n11933) );
  NOR2X1 U13042 ( .A(n6992), .B(n7410), .Y(n12567) );
  NOR2X1 U13043 ( .A(n10328), .B(n11934), .Y(n12579) );
  NAND2X1 U13044 ( .A(n12582), .B(n12577), .Y(n11934) );
  NOR2X1 U13045 ( .A(n10982), .B(n11935), .Y(n12578) );
  NAND2X1 U13046 ( .A(n12577), .B(n12570), .Y(n11935) );
  NOR2X1 U13047 ( .A(n6981), .B(n6971), .Y(n12570) );
  NOR4X1 U13048 ( .A(n12583), .B(n12584), .C(n12585), .D(n9908), .Y(n12557) );
  NOR2X1 U13049 ( .A(n10310), .B(n11939), .Y(n12585) );
  NAND2X1 U13050 ( .A(n12576), .B(n12571), .Y(n11939) );
  NOR2X1 U13051 ( .A(n7379), .B(n7387), .Y(n12576) );
  NOR2X1 U13052 ( .A(n10322), .B(n11940), .Y(n12584) );
  NAND2X1 U13053 ( .A(n12582), .B(n12571), .Y(n11940) );
  NOR2X1 U13054 ( .A(n9615), .B(n7410), .Y(n12571) );
  INVX1 U13055 ( .A(n7003), .Y(n7410) );
  NOR2X1 U13056 ( .A(n7379), .B(n6981), .Y(n12582) );
  NOR2X1 U13057 ( .A(n10983), .B(n11941), .Y(n12583) );
  NAND2X1 U13058 ( .A(n12577), .B(n12565), .Y(n11941) );
  NOR2X1 U13059 ( .A(n6971), .B(n7387), .Y(n12565) );
  INVX1 U13060 ( .A(n6981), .Y(n7387) );
  NAND2X1 U13061 ( .A(n12586), .B(n12587), .Y(n6981) );
  NAND2X1 U13062 ( .A(n12588), .B(n12589), .Y(n12587) );
  NAND2X1 U13063 ( .A(n12590), .B(n12591), .Y(n12588) );
  NAND2X1 U13064 ( .A(n12592), .B(n12590), .Y(n12586) );
  INVX1 U13065 ( .A(n12593), .Y(n12592) );
  INVX1 U13066 ( .A(n7379), .Y(n6971) );
  ADDHXL U13067 ( .A(n12594), .B(n12593), .S(n7379) );
  NAND2X1 U13068 ( .A(n12595), .B(n12596), .Y(n12594) );
  NOR2X1 U13069 ( .A(n7003), .B(n6992), .Y(n12577) );
  INVX1 U13070 ( .A(n9615), .Y(n6992) );
  ADDHXL U13071 ( .A(n12597), .B(n12598), .S(n9615) );
  NAND2X1 U13072 ( .A(n12599), .B(n12600), .Y(n12597) );
  ADDHXL U13073 ( .A(n7564), .B(n12601), .S(n7003) );
  NOR2X1 U13074 ( .A(n12602), .B(n12603), .Y(n12601) );
  INVX1 U13075 ( .A(n12604), .Y(n12602) );
  NAND2X1 U13076 ( .A(n11809), .B(n10876), .Y(n12555) );
  NAND4X1 U13077 ( .A(n12605), .B(n12606), .C(n12607), .D(n12608), .Y(n10876)
         );
  NOR4X1 U13078 ( .A(n12609), .B(n12610), .C(n12611), .D(n12612), .Y(n12608)
         );
  NOR2X1 U13079 ( .A(n10312), .B(n11818), .Y(n12612) );
  NAND2X1 U13080 ( .A(n12613), .B(n12614), .Y(n11818) );
  NOR2X1 U13081 ( .A(n10314), .B(n11819), .Y(n12611) );
  NAND2X1 U13082 ( .A(n12615), .B(n12613), .Y(n11819) );
  NOR2X1 U13083 ( .A(n10316), .B(n11820), .Y(n12610) );
  NAND2X1 U13084 ( .A(n12613), .B(n12616), .Y(n11820) );
  NOR2X1 U13085 ( .A(n10324), .B(n11821), .Y(n12609) );
  NAND2X1 U13086 ( .A(n12617), .B(n12614), .Y(n11821) );
  NOR4X1 U13087 ( .A(n12618), .B(n12619), .C(n12620), .D(n12621), .Y(n12607)
         );
  NOR2X1 U13088 ( .A(n10326), .B(n11826), .Y(n12621) );
  NAND2X1 U13089 ( .A(n12615), .B(n12617), .Y(n11826) );
  NOR2X1 U13090 ( .A(n10328), .B(n11827), .Y(n12620) );
  NAND2X1 U13091 ( .A(n12616), .B(n12617), .Y(n11827) );
  NOR2X1 U13092 ( .A(n10972), .B(n11828), .Y(n12619) );
  NAND2X1 U13093 ( .A(n12622), .B(n12614), .Y(n11828) );
  NOR2X1 U13094 ( .A(n10967), .B(n11829), .Y(n12618) );
  NAND2X1 U13095 ( .A(n12622), .B(n12615), .Y(n11829) );
  NOR4X1 U13096 ( .A(n12623), .B(n12624), .C(n12625), .D(n12626), .Y(n12606)
         );
  NOR2X1 U13097 ( .A(n10983), .B(n11834), .Y(n12626) );
  NAND2X1 U13098 ( .A(n12622), .B(n12616), .Y(n11834) );
  NOR2X1 U13099 ( .A(n10965), .B(n11835), .Y(n12625) );
  NAND2X1 U13100 ( .A(n12627), .B(n12614), .Y(n11835) );
  NOR2X1 U13101 ( .A(n7001), .B(n12628), .Y(n12614) );
  NOR2X1 U13102 ( .A(n10964), .B(n11836), .Y(n12624) );
  NAND2X1 U13103 ( .A(n12627), .B(n12615), .Y(n11836) );
  NOR2X1 U13104 ( .A(n7421), .B(n6990), .Y(n12615) );
  NOR2X1 U13105 ( .A(n10982), .B(n11837), .Y(n12623) );
  NAND2X1 U13106 ( .A(n12627), .B(n12616), .Y(n11837) );
  NOR2X1 U13107 ( .A(n7001), .B(n6990), .Y(n12616) );
  NOR4X1 U13108 ( .A(n12629), .B(n12630), .C(n12631), .D(n12632), .Y(n12605)
         );
  NOR2X1 U13109 ( .A(n10310), .B(n11842), .Y(n12632) );
  NAND2X1 U13110 ( .A(n12633), .B(n12613), .Y(n11842) );
  NOR2X1 U13111 ( .A(n7392), .B(n9176), .Y(n12613) );
  NOR2X1 U13112 ( .A(n10322), .B(n11843), .Y(n12631) );
  NAND2X1 U13113 ( .A(n12633), .B(n12617), .Y(n11843) );
  NOR2X1 U13114 ( .A(n9176), .B(n6979), .Y(n12617) );
  NOR2X1 U13115 ( .A(n10973), .B(n11844), .Y(n12630) );
  NAND2X1 U13116 ( .A(n12633), .B(n12622), .Y(n11844) );
  NOR2X1 U13117 ( .A(n7392), .B(n6969), .Y(n12622) );
  NOR2X1 U13118 ( .A(n10966), .B(n11845), .Y(n12629) );
  NAND2X1 U13119 ( .A(n12633), .B(n12627), .Y(n11845) );
  NOR2X1 U13120 ( .A(n6969), .B(n6979), .Y(n12627) );
  INVX1 U13121 ( .A(n7392), .Y(n6979) );
  NOR2X1 U13122 ( .A(n12628), .B(n7421), .Y(n12633) );
  INVX1 U13123 ( .A(n7001), .Y(n7421) );
  NAND2X1 U13124 ( .A(n10256), .B(n12634), .Y(n12554) );
  NAND4X1 U13125 ( .A(n12635), .B(n12636), .C(n12637), .D(n12638), .Y(n12634)
         );
  NOR4X1 U13126 ( .A(n12639), .B(n12640), .C(n12641), .D(n12642), .Y(n12638)
         );
  NOR2X1 U13127 ( .A(n10310), .B(n11877), .Y(n12642) );
  NAND2X1 U13128 ( .A(n12643), .B(n12644), .Y(n11877) );
  NOR2X1 U13129 ( .A(n10312), .B(n11878), .Y(n12641) );
  NAND2X1 U13130 ( .A(n12643), .B(n12645), .Y(n11878) );
  NOR2X1 U13131 ( .A(n10314), .B(n11879), .Y(n12640) );
  NAND2X1 U13132 ( .A(n12644), .B(n12646), .Y(n11879) );
  NOR2X1 U13133 ( .A(n10316), .B(n11880), .Y(n12639) );
  NAND2X1 U13134 ( .A(n12646), .B(n12645), .Y(n11880) );
  NOR4X1 U13135 ( .A(n12647), .B(n12648), .C(n12649), .D(n12650), .Y(n12637)
         );
  NOR2X1 U13136 ( .A(n10322), .B(n11885), .Y(n12650) );
  NAND2X1 U13137 ( .A(n12651), .B(n12644), .Y(n11885) );
  NOR2X1 U13138 ( .A(n10324), .B(n11886), .Y(n12649) );
  NAND2X1 U13139 ( .A(n12651), .B(n12645), .Y(n11886) );
  NOR2X1 U13140 ( .A(n10326), .B(n11887), .Y(n12648) );
  NAND2X1 U13141 ( .A(n12652), .B(n12644), .Y(n11887) );
  NOR2X1 U13142 ( .A(n12653), .B(G21561), .Y(n12644) );
  NOR2X1 U13143 ( .A(n10328), .B(n11888), .Y(n12647) );
  NAND2X1 U13144 ( .A(n12652), .B(n12645), .Y(n11888) );
  NOR2X1 U13145 ( .A(n12653), .B(n8890), .Y(n12645) );
  NOR4X1 U13146 ( .A(n12654), .B(n12655), .C(n12656), .D(n12657), .Y(n12636)
         );
  NOR2X1 U13147 ( .A(n10973), .B(n11893), .Y(n12657) );
  NAND2X1 U13148 ( .A(n12658), .B(n12643), .Y(n11893) );
  NOR2X1 U13149 ( .A(n10972), .B(n11894), .Y(n12656) );
  NAND2X1 U13150 ( .A(n12659), .B(n12643), .Y(n11894) );
  AND2X1 U13151 ( .A(n9157), .B(n9139), .Y(n12643) );
  NOR2X1 U13152 ( .A(n10967), .B(n11895), .Y(n12655) );
  NAND2X1 U13153 ( .A(n12658), .B(n12646), .Y(n11895) );
  NOR2X1 U13154 ( .A(n10983), .B(n11896), .Y(n12654) );
  NAND2X1 U13155 ( .A(n12659), .B(n12646), .Y(n11896) );
  AND2X1 U13156 ( .A(n12660), .B(n9157), .Y(n12646) );
  NOR4X1 U13157 ( .A(n12661), .B(n12662), .C(n12663), .D(n12664), .Y(n12635)
         );
  NOR2X1 U13158 ( .A(n10966), .B(n11901), .Y(n12664) );
  NAND2X1 U13159 ( .A(n12658), .B(n12651), .Y(n11901) );
  NOR2X1 U13160 ( .A(n10965), .B(n11902), .Y(n12663) );
  NAND2X1 U13161 ( .A(n12659), .B(n12651), .Y(n11902) );
  NOR2X1 U13162 ( .A(n9157), .B(n12660), .Y(n12651) );
  NOR2X1 U13163 ( .A(n10964), .B(n11903), .Y(n12662) );
  NAND2X1 U13164 ( .A(n12658), .B(n12652), .Y(n11903) );
  NOR2X1 U13165 ( .A(n9196), .B(G21561), .Y(n12658) );
  NOR2X1 U13166 ( .A(n10982), .B(n11904), .Y(n12661) );
  NAND2X1 U13167 ( .A(n12659), .B(n12652), .Y(n11904) );
  NOR2X1 U13168 ( .A(n9157), .B(n9139), .Y(n12652) );
  INVX1 U13169 ( .A(n12660), .Y(n9139) );
  NOR2X1 U13170 ( .A(n9135), .B(n10944), .Y(n12660) );
  NAND2X1 U13171 ( .A(n12665), .B(n12666), .Y(n9157) );
  NAND2X1 U13172 ( .A(n12667), .B(n12668), .Y(n12666) );
  NAND2X1 U13173 ( .A(n9076), .B(n8893), .Y(n12668) );
  INVX1 U13174 ( .A(n12669), .Y(n12667) );
  NAND2X1 U13175 ( .A(n10952), .B(n12670), .Y(n12665) );
  NOR2X1 U13176 ( .A(n8890), .B(n9196), .Y(n12659) );
  INVX1 U13177 ( .A(n12653), .Y(n9196) );
  ADDHXL U13178 ( .A(n12669), .B(n8870), .S(n12653) );
  NAND2X1 U13179 ( .A(n12671), .B(n12670), .Y(n12669) );
  NAND2X1 U13180 ( .A(n12672), .B(n10952), .Y(n12670) );
  ADDHXL U13181 ( .A(n9076), .B(n8893), .S(n12672) );
  NAND2X1 U13182 ( .A(G21559), .B(n8711), .Y(n12671) );
  NAND2X1 U13183 ( .A(n12011), .B(n12673), .Y(n12553) );
  NAND4X1 U13184 ( .A(n12674), .B(n12675), .C(n12676), .D(n12677), .Y(n9931)
         );
  NOR2X1 U13185 ( .A(n12678), .B(n12679), .Y(n12677) );
  AND2X1 U13186 ( .A(n6915), .B(n9926), .Y(n12679) );
  NOR2X1 U13187 ( .A(n10217), .B(n9552), .Y(n12678) );
  NAND2X1 U13188 ( .A(G21575), .B(n10444), .Y(n12676) );
  OR2X1 U13189 ( .A(n12682), .B(n6917), .Y(n12680) );
  NAND2X1 U13190 ( .A(n11705), .B(G21766), .Y(n12674) );
  INVX1 U13191 ( .A(n9922), .Y(n9924) );
  NAND4X1 U13192 ( .A(n12683), .B(n12684), .C(n12685), .D(n12686), .Y(n9922)
         );
  NOR2X1 U13193 ( .A(n12687), .B(n12688), .Y(n12686) );
  NOR2X1 U13194 ( .A(n7314), .B(n9908), .Y(n12688) );
  NOR2X1 U13195 ( .A(n10217), .B(n7310), .Y(n12687) );
  NAND2X1 U13196 ( .A(G21576), .B(n10444), .Y(n12685) );
  NAND2X1 U13197 ( .A(n10256), .B(n12689), .Y(n12684) );
  ADDFXL U13198 ( .A(n12690), .B(n12681), .CI(n7310), .S(n12689) );
  NAND2X1 U13199 ( .A(n11705), .B(G21767), .Y(n12683) );
  NAND4X1 U13200 ( .A(n12691), .B(n12692), .C(n12693), .D(n12694), .Y(n9911)
         );
  NOR2X1 U13201 ( .A(n12695), .B(n12696), .Y(n12694) );
  NOR2X1 U13202 ( .A(n7299), .B(n9908), .Y(n12696) );
  INVX1 U13203 ( .A(n6883), .Y(n7299) );
  NOR2X1 U13204 ( .A(n10217), .B(n6886), .Y(n12695) );
  NAND2X1 U13205 ( .A(G21577), .B(n10444), .Y(n12693) );
  ADDFXL U13206 ( .A(n12698), .B(n6886), .CI(n12699), .S(n12697) );
  NAND2X1 U13207 ( .A(n11705), .B(G21768), .Y(n12691) );
  INVX1 U13208 ( .A(n11698), .Y(n11695) );
  NAND4X1 U13209 ( .A(n12700), .B(n12701), .C(n12702), .D(n12703), .Y(n11698)
         );
  NOR2X1 U13210 ( .A(n12704), .B(n12705), .Y(n12703) );
  AND2X1 U13211 ( .A(n9926), .B(n7291), .Y(n12705) );
  NOR2X1 U13212 ( .A(n10217), .B(n9525), .Y(n12704) );
  INVX1 U13213 ( .A(n7290), .Y(n9525) );
  NOR2X1 U13214 ( .A(n12011), .B(n11809), .Y(n10217) );
  NOR3X1 U13215 ( .A(n9092), .B(n7451), .C(n12707), .Y(n11809) );
  NAND2X1 U13216 ( .A(G21578), .B(n10444), .Y(n12702) );
  NAND3X1 U13217 ( .A(n12060), .B(n12708), .C(n9193), .Y(n10444) );
  NAND2X1 U13218 ( .A(n10256), .B(n12709), .Y(n12701) );
  ADDFXL U13219 ( .A(n7290), .B(n11709), .CI(n11711), .S(n12709) );
  NAND2X1 U13220 ( .A(n12710), .B(n12711), .Y(n11711) );
  NAND2X1 U13221 ( .A(n12712), .B(n12713), .Y(n12711) );
  OR2X1 U13222 ( .A(n12699), .B(n6886), .Y(n12713) );
  INVX1 U13223 ( .A(n12698), .Y(n12712) );
  NAND2X1 U13224 ( .A(n12699), .B(n6886), .Y(n12710) );
  INVX1 U13225 ( .A(n9720), .Y(n6886) );
  NOR2X1 U13226 ( .A(n12714), .B(n11715), .Y(n9720) );
  AND2X1 U13227 ( .A(n12715), .B(n12716), .Y(n12714) );
  OR2X1 U13228 ( .A(n12717), .B(n12718), .Y(n12716) );
  NAND2X1 U13229 ( .A(n12719), .B(n12720), .Y(n12699) );
  NAND2X1 U13230 ( .A(n12721), .B(n12722), .Y(n12720) );
  OR2X1 U13231 ( .A(n12681), .B(n7310), .Y(n12722) );
  INVX1 U13232 ( .A(n12690), .Y(n12721) );
  NAND2X1 U13233 ( .A(n7310), .B(n12681), .Y(n12719) );
  NAND2X1 U13234 ( .A(n6917), .B(n12682), .Y(n12681) );
  INVX1 U13235 ( .A(n9552), .Y(n6917) );
  NAND2X1 U13236 ( .A(n12717), .B(n12723), .Y(n9552) );
  NAND3X1 U13237 ( .A(n12724), .B(n12550), .C(n12725), .Y(n12723) );
  ADDHXL U13238 ( .A(n9085), .B(n12726), .S(n12725) );
  INVX1 U13239 ( .A(n6906), .Y(n7310) );
  ADDHXL U13240 ( .A(n12717), .B(n12718), .S(n6906) );
  INVX1 U13241 ( .A(n12727), .Y(n11709) );
  ADDHXL U13242 ( .A(n11714), .B(n11715), .S(n7290) );
  NOR3X1 U13243 ( .A(n12718), .B(n12717), .C(n12715), .Y(n11715) );
  ADDHXL U13244 ( .A(n12728), .B(n9085), .S(n12715) );
  NAND4X1 U13245 ( .A(n12729), .B(n12730), .C(n12731), .D(n12732), .Y(n12728)
         );
  NAND2X1 U13246 ( .A(n10272), .B(n6883), .Y(n12732) );
  NAND2X1 U13247 ( .A(n12733), .B(n12734), .Y(n6883) );
  NAND2X1 U13248 ( .A(n12735), .B(n12736), .Y(n12734) );
  NAND2X1 U13249 ( .A(n12737), .B(n12738), .Y(n12735) );
  NAND2X1 U13250 ( .A(n12739), .B(n12737), .Y(n12733) );
  INVX1 U13251 ( .A(n11754), .Y(n12739) );
  NAND2X1 U13252 ( .A(G21577), .B(n10224), .Y(n12731) );
  NAND2X1 U13253 ( .A(G21609), .B(n10225), .Y(n12730) );
  NAND2X1 U13254 ( .A(G21768), .B(n9260), .Y(n12729) );
  NAND2X1 U13255 ( .A(n12740), .B(n12741), .Y(n12717) );
  NAND2X1 U13256 ( .A(n12724), .B(n12550), .Y(n12741) );
  NAND3X1 U13257 ( .A(n9755), .B(G21549), .C(n12742), .Y(n12550) );
  ADDHXL U13258 ( .A(n7564), .B(n12743), .S(n12742) );
  NAND2X1 U13259 ( .A(n12548), .B(n12551), .Y(n12724) );
  NAND2X1 U13260 ( .A(n12744), .B(n12745), .Y(n12551) );
  NAND2X1 U13261 ( .A(n9755), .B(G21549), .Y(n12745) );
  ADDHXL U13262 ( .A(n9085), .B(n12743), .S(n12744) );
  NAND4X1 U13263 ( .A(n12746), .B(n12747), .C(n12748), .D(n12749), .Y(n12743)
         );
  NAND2X1 U13264 ( .A(n6926), .B(n10272), .Y(n12749) );
  AND2X1 U13265 ( .A(n12750), .B(n12751), .Y(n6926) );
  NAND2X1 U13266 ( .A(n12752), .B(n12753), .Y(n12751) );
  NAND2X1 U13267 ( .A(G21574), .B(n10224), .Y(n12748) );
  NAND2X1 U13268 ( .A(G21606), .B(n10225), .Y(n12747) );
  NAND2X1 U13269 ( .A(G21765), .B(n9260), .Y(n12746) );
  NAND2X1 U13270 ( .A(n12540), .B(n12539), .Y(n12548) );
  NAND3X1 U13271 ( .A(n9755), .B(G21550), .C(n12754), .Y(n12539) );
  ADDHXL U13272 ( .A(n12755), .B(n7564), .S(n12754) );
  NAND2X1 U13273 ( .A(n12543), .B(n12756), .Y(n12540) );
  NAND2X1 U13274 ( .A(n12542), .B(n12441), .Y(n12756) );
  NAND3X1 U13275 ( .A(n9755), .B(G21551), .C(n12757), .Y(n12441) );
  ADDHXL U13276 ( .A(n12758), .B(n7564), .S(n12757) );
  NAND2X1 U13277 ( .A(n12442), .B(n12439), .Y(n12542) );
  NAND2X1 U13278 ( .A(n12255), .B(n12759), .Y(n12439) );
  NAND2X1 U13279 ( .A(n12256), .B(n12253), .Y(n12759) );
  NAND2X1 U13280 ( .A(n12596), .B(n12760), .Y(n12253) );
  NAND2X1 U13281 ( .A(n12593), .B(n12595), .Y(n12760) );
  NAND2X1 U13282 ( .A(n12761), .B(n12762), .Y(n12595) );
  NAND2X1 U13283 ( .A(n9755), .B(G21553), .Y(n12762) );
  ADDHXL U13284 ( .A(n12763), .B(n9085), .S(n12761) );
  NAND2X1 U13285 ( .A(n12591), .B(n12764), .Y(n12593) );
  NAND2X1 U13286 ( .A(n12589), .B(n12590), .Y(n12764) );
  NAND4X1 U13287 ( .A(n12765), .B(n12766), .C(n12767), .D(n8804), .Y(n12590)
         );
  ADDHXL U13288 ( .A(n9085), .B(n12768), .S(n12765) );
  NAND2X1 U13289 ( .A(n12600), .B(n12769), .Y(n12589) );
  NAND2X1 U13290 ( .A(n12598), .B(n12599), .Y(n12769) );
  NAND2X1 U13291 ( .A(n12770), .B(n12771), .Y(n12599) );
  ADDHXL U13292 ( .A(n9085), .B(n12772), .S(n12771) );
  INVX1 U13293 ( .A(n12773), .Y(n12770) );
  NAND2X1 U13294 ( .A(n12604), .B(n12774), .Y(n12598) );
  OR2X1 U13295 ( .A(n9085), .B(n12603), .Y(n12774) );
  NOR2X1 U13296 ( .A(n12775), .B(n12776), .Y(n12603) );
  NAND2X1 U13297 ( .A(n12776), .B(n12775), .Y(n12604) );
  NAND4X1 U13298 ( .A(n12777), .B(n12778), .C(n12767), .D(n8783), .Y(n12775)
         );
  NAND2X1 U13299 ( .A(G21428), .B(n12779), .Y(n12778) );
  NAND4X1 U13300 ( .A(n12780), .B(n12781), .C(n12782), .D(n12783), .Y(n12779)
         );
  NOR4X1 U13301 ( .A(n9185), .B(n12784), .C(n12785), .D(n12786), .Y(n12783) );
  NOR2X1 U13302 ( .A(n9751), .B(n12787), .Y(n12786) );
  NOR2X1 U13303 ( .A(n12707), .B(n9278), .Y(n12785) );
  NOR2X1 U13304 ( .A(n12788), .B(n12789), .Y(n12782) );
  NAND2X1 U13305 ( .A(n9751), .B(n7442), .Y(n12781) );
  NAND2X1 U13306 ( .A(n12790), .B(n8772), .Y(n12780) );
  NAND2X1 U13307 ( .A(n9755), .B(G21556), .Y(n12777) );
  ADDHXL U13308 ( .A(n12791), .B(n7564), .S(n12776) );
  NAND4X1 U13309 ( .A(n12792), .B(n12793), .C(n12794), .D(n12795), .Y(n12791)
         );
  NOR2X1 U13310 ( .A(n12796), .B(n12797), .Y(n12795) );
  NOR2X1 U13311 ( .A(n10426), .B(n11440), .Y(n12797) );
  NOR2X1 U13312 ( .A(n12798), .B(n8890), .Y(n12796) );
  NAND2X1 U13313 ( .A(n7001), .B(n10272), .Y(n12794) );
  ADDHXL U13314 ( .A(n9260), .B(n12799), .S(n7001) );
  NOR2X1 U13315 ( .A(n12800), .B(n12801), .Y(n12799) );
  INVX1 U13316 ( .A(n12802), .Y(n12800) );
  NAND2X1 U13317 ( .A(G21599), .B(n10225), .Y(n12793) );
  NAND2X1 U13318 ( .A(G21758), .B(n9260), .Y(n12792) );
  NAND2X1 U13319 ( .A(n12803), .B(n12773), .Y(n12600) );
  NAND4X1 U13320 ( .A(n12804), .B(n12805), .C(n12806), .D(n12807), .Y(n12773)
         );
  NOR3X1 U13321 ( .A(n12808), .B(n9260), .C(n9071), .Y(n12807) );
  NOR4X1 U13322 ( .A(n12809), .B(n9223), .C(n11987), .D(n12810), .Y(n12808) );
  OR2X1 U13323 ( .A(n12811), .B(n7451), .Y(n12805) );
  NAND2X1 U13324 ( .A(n9755), .B(G21555), .Y(n12804) );
  ADDHXL U13325 ( .A(n7564), .B(n12772), .S(n12803) );
  NAND4X1 U13326 ( .A(n12812), .B(n12813), .C(n12814), .D(n12815), .Y(n12772)
         );
  NOR2X1 U13327 ( .A(n12816), .B(n12817), .Y(n12815) );
  NOR2X1 U13328 ( .A(n10227), .B(n6989), .Y(n12817) );
  INVX1 U13329 ( .A(G21759), .Y(n6989) );
  NOR2X1 U13330 ( .A(n10271), .B(n6988), .Y(n12816) );
  NAND2X1 U13331 ( .A(G21568), .B(n10224), .Y(n12814) );
  NAND2X1 U13332 ( .A(n6990), .B(n10272), .Y(n12813) );
  INVX1 U13333 ( .A(n12628), .Y(n6990) );
  ADDHXL U13334 ( .A(n12818), .B(n12819), .S(n12628) );
  NAND2X1 U13335 ( .A(n12820), .B(n12821), .Y(n12818) );
  NAND2X1 U13336 ( .A(G21560), .B(n12822), .Y(n12812) );
  NAND2X1 U13337 ( .A(n12823), .B(n12824), .Y(n12591) );
  NAND3X1 U13338 ( .A(n12767), .B(n8804), .C(n12766), .Y(n12824) );
  NAND2X1 U13339 ( .A(n9755), .B(G21554), .Y(n12766) );
  ADDHXL U13340 ( .A(n7564), .B(n12768), .S(n12823) );
  NAND4X1 U13341 ( .A(n12825), .B(n12826), .C(n12827), .D(n12828), .Y(n12768)
         );
  NAND2X1 U13342 ( .A(G21569), .B(n10224), .Y(n12828) );
  NOR2X1 U13343 ( .A(n12829), .B(n12830), .Y(n12827) );
  NOR2X1 U13344 ( .A(n12798), .B(n8893), .Y(n12830) );
  NOR2X1 U13345 ( .A(n10613), .B(n7392), .Y(n12829) );
  NAND2X1 U13346 ( .A(n12831), .B(n12832), .Y(n7392) );
  NAND2X1 U13347 ( .A(n12833), .B(n12834), .Y(n12831) );
  NAND2X1 U13348 ( .A(G21601), .B(n10225), .Y(n12826) );
  NAND2X1 U13349 ( .A(G21760), .B(n9260), .Y(n12825) );
  NAND3X1 U13350 ( .A(n9755), .B(G21553), .C(n12835), .Y(n12596) );
  ADDHXL U13351 ( .A(n7564), .B(n12763), .S(n12835) );
  NAND4X1 U13352 ( .A(n12836), .B(n12837), .C(n12838), .D(n12839), .Y(n12763)
         );
  NOR2X1 U13353 ( .A(n12840), .B(n12841), .Y(n12839) );
  NOR2X1 U13354 ( .A(n12798), .B(n8870), .Y(n12841) );
  INVX1 U13355 ( .A(n12822), .Y(n12798) );
  NAND4X1 U13356 ( .A(n12842), .B(n8783), .C(n12843), .D(n10012), .Y(n12822)
         );
  INVX1 U13357 ( .A(n10236), .Y(n10012) );
  NAND2X1 U13358 ( .A(G21428), .B(n12844), .Y(n12842) );
  NAND2X1 U13359 ( .A(n7423), .B(n12845), .Y(n12844) );
  NAND2X1 U13360 ( .A(n12790), .B(n8861), .Y(n12845) );
  INVX1 U13361 ( .A(n12706), .Y(n12790) );
  NAND2X1 U13362 ( .A(n9092), .B(n7444), .Y(n12706) );
  AND3X1 U13363 ( .A(n9197), .B(n9216), .C(n12846), .Y(n7423) );
  NAND2X1 U13364 ( .A(n12847), .B(n9076), .Y(n9197) );
  NOR2X1 U13365 ( .A(n10426), .B(n7375), .Y(n12840) );
  INVX1 U13366 ( .A(G21570), .Y(n7375) );
  INVX1 U13367 ( .A(n10224), .Y(n10426) );
  NAND2X1 U13368 ( .A(n6969), .B(n10272), .Y(n12838) );
  INVX1 U13369 ( .A(n9176), .Y(n6969) );
  ADDHXL U13370 ( .A(n12848), .B(n12832), .S(n9176) );
  NAND2X1 U13371 ( .A(G21761), .B(n9260), .Y(n12837) );
  NAND2X1 U13372 ( .A(G21602), .B(n10225), .Y(n12836) );
  NAND2X1 U13373 ( .A(n12849), .B(n12850), .Y(n12256) );
  NAND2X1 U13374 ( .A(n9755), .B(G21552), .Y(n12850) );
  ADDHXL U13375 ( .A(n9085), .B(n12851), .S(n12849) );
  NAND3X1 U13376 ( .A(n9755), .B(G21552), .C(n12852), .Y(n12255) );
  ADDHXL U13377 ( .A(n12851), .B(n7564), .S(n12852) );
  NAND4X1 U13378 ( .A(n12853), .B(n12854), .C(n12855), .D(n12856), .Y(n12851)
         );
  NOR2X1 U13379 ( .A(n12857), .B(n12858), .Y(n12856) );
  NOR2X1 U13380 ( .A(n10227), .B(n6958), .Y(n12858) );
  INVX1 U13381 ( .A(G21762), .Y(n6958) );
  NOR2X1 U13382 ( .A(n10271), .B(n6957), .Y(n12857) );
  INVX1 U13383 ( .A(G21603), .Y(n6957) );
  NAND2X1 U13384 ( .A(G21571), .B(n10224), .Y(n12855) );
  NAND2X1 U13385 ( .A(G21557), .B(n12859), .Y(n12854) );
  NAND2X1 U13386 ( .A(n12843), .B(n12860), .Y(n12859) );
  NAND2X1 U13387 ( .A(n9175), .B(G21428), .Y(n12860) );
  INVX1 U13388 ( .A(n9216), .Y(n9175) );
  NAND2X1 U13389 ( .A(n9647), .B(n9185), .Y(n9216) );
  INVX1 U13390 ( .A(n8858), .Y(n9647) );
  NAND2X1 U13391 ( .A(n6959), .B(n10272), .Y(n12853) );
  NOR2X1 U13392 ( .A(n12861), .B(n12862), .Y(n6959) );
  AND2X1 U13393 ( .A(n12863), .B(n12864), .Y(n12861) );
  NAND2X1 U13394 ( .A(n12865), .B(n12848), .Y(n12864) );
  NAND2X1 U13395 ( .A(n12866), .B(n12867), .Y(n12442) );
  NAND2X1 U13396 ( .A(n9755), .B(G21551), .Y(n12867) );
  ADDHXL U13397 ( .A(n9085), .B(n12758), .S(n12866) );
  NAND4X1 U13398 ( .A(n12868), .B(n12869), .C(n12870), .D(n12871), .Y(n12758)
         );
  NAND2X1 U13399 ( .A(n6948), .B(n10272), .Y(n12871) );
  ADDHXL U13400 ( .A(n12872), .B(n12862), .S(n6948) );
  NAND2X1 U13401 ( .A(G21572), .B(n10224), .Y(n12870) );
  NAND2X1 U13402 ( .A(G21604), .B(n10225), .Y(n12869) );
  NAND2X1 U13403 ( .A(G21763), .B(n9260), .Y(n12868) );
  NAND2X1 U13404 ( .A(n12873), .B(n12874), .Y(n12543) );
  NAND2X1 U13405 ( .A(n9755), .B(G21550), .Y(n12874) );
  ADDHXL U13406 ( .A(n9085), .B(n12755), .S(n12873) );
  NAND4X1 U13407 ( .A(n12875), .B(n12876), .C(n12877), .D(n12878), .Y(n12755)
         );
  NAND2X1 U13408 ( .A(n6937), .B(n10272), .Y(n12878) );
  ADDHXL U13409 ( .A(n12879), .B(n12880), .S(n6937) );
  NAND2X1 U13410 ( .A(G21573), .B(n10224), .Y(n12877) );
  NAND2X1 U13411 ( .A(G21605), .B(n10225), .Y(n12876) );
  NAND2X1 U13412 ( .A(G21764), .B(n9260), .Y(n12875) );
  ADDHXL U13413 ( .A(n7564), .B(n12726), .S(n12740) );
  NAND4X1 U13414 ( .A(n12881), .B(n12882), .C(n12883), .D(n12884), .Y(n12726)
         );
  NAND2X1 U13415 ( .A(n6915), .B(n10272), .Y(n12884) );
  ADDHXL U13416 ( .A(n12885), .B(n12750), .S(n6915) );
  INVX1 U13417 ( .A(n12886), .Y(n12750) );
  NAND2X1 U13418 ( .A(n12887), .B(n12888), .Y(n12885) );
  NAND2X1 U13419 ( .A(G21575), .B(n10224), .Y(n12883) );
  NAND2X1 U13420 ( .A(G21607), .B(n10225), .Y(n12882) );
  NAND2X1 U13421 ( .A(G21766), .B(n9260), .Y(n12881) );
  ADDHXL U13422 ( .A(n7564), .B(n12889), .S(n12718) );
  NOR4X1 U13423 ( .A(n12890), .B(n12891), .C(n12892), .D(n12893), .Y(n12889)
         );
  NOR2X1 U13424 ( .A(n10227), .B(n6900), .Y(n12893) );
  INVX1 U13425 ( .A(G21767), .Y(n6900) );
  NOR2X1 U13426 ( .A(n10271), .B(n6899), .Y(n12892) );
  INVX1 U13427 ( .A(G21608), .Y(n6899) );
  AND2X1 U13428 ( .A(n10224), .B(G21576), .Y(n12891) );
  NOR2X1 U13429 ( .A(n10613), .B(n7314), .Y(n12890) );
  INVX1 U13430 ( .A(n6902), .Y(n7314) );
  ADDHXL U13431 ( .A(n12894), .B(n12895), .S(n6902) );
  AND2X1 U13432 ( .A(n12896), .B(n12897), .Y(n12895) );
  ADDHXL U13433 ( .A(n12898), .B(n7564), .S(n11714) );
  NAND4X1 U13434 ( .A(n12899), .B(n12900), .C(n12901), .D(n12902), .Y(n12898)
         );
  NAND2X1 U13435 ( .A(G21578), .B(n10224), .Y(n12902) );
  NAND4X1 U13436 ( .A(n12903), .B(n12811), .C(n12904), .D(n12767), .Y(n10224)
         );
  NAND4X1 U13437 ( .A(G21428), .B(n8772), .C(n7446), .D(n12905), .Y(n12767) );
  NOR2X1 U13438 ( .A(n12809), .B(n11847), .Y(n12905) );
  INVX1 U13439 ( .A(n12011), .Y(n11847) );
  NOR2X1 U13440 ( .A(n12906), .B(n9076), .Y(n12011) );
  NAND2X1 U13441 ( .A(G21428), .B(n7417), .Y(n12904) );
  NAND2X1 U13442 ( .A(n9172), .B(n12907), .Y(n7417) );
  AND2X1 U13443 ( .A(n12908), .B(n12909), .Y(n9172) );
  NAND2X1 U13444 ( .A(n12910), .B(n12784), .Y(n12909) );
  NAND2X1 U13445 ( .A(n12847), .B(n8711), .Y(n12908) );
  INVX1 U13446 ( .A(n12911), .Y(n12847) );
  NAND2X1 U13447 ( .A(n7291), .B(n10272), .Y(n12901) );
  INVX1 U13448 ( .A(n10613), .Y(n10272) );
  NOR2X1 U13449 ( .A(n7564), .B(n9755), .Y(n10613) );
  NAND2X1 U13450 ( .A(G21610), .B(n10225), .Y(n12900) );
  NAND2X1 U13451 ( .A(G21769), .B(n9260), .Y(n12899) );
  NAND2X1 U13452 ( .A(G21769), .B(n11705), .Y(n12700) );
  NOR3X1 U13453 ( .A(n7444), .B(n10116), .C(n11987), .Y(n11705) );
  NAND2X1 U13454 ( .A(n7291), .B(n6882), .Y(n11755) );
  NAND3X1 U13455 ( .A(n9070), .B(n8817), .C(n8897), .Y(n12912) );
  OR2X1 U13456 ( .A(n9257), .B(n9258), .Y(n9269) );
  NAND3X1 U13457 ( .A(n8861), .B(G21426), .C(n9646), .Y(n9258) );
  INVX1 U13458 ( .A(n7441), .Y(n9257) );
  NOR2X1 U13459 ( .A(n12913), .B(n12914), .Y(n7441) );
  AND4X1 U13460 ( .A(n12915), .B(n12916), .C(n12917), .D(n12918), .Y(n12914)
         );
  NAND3X1 U13461 ( .A(n12919), .B(n12920), .C(n12921), .Y(n12918) );
  OR2X1 U13462 ( .A(n12922), .B(n7444), .Y(n12921) );
  NAND3X1 U13463 ( .A(n12923), .B(n12708), .C(n12924), .Y(n12920) );
  INVX1 U13464 ( .A(n12925), .Y(n12924) );
  NAND2X1 U13465 ( .A(n9059), .B(n12926), .Y(n12923) );
  OR2X1 U13466 ( .A(n12926), .B(n9059), .Y(n12919) );
  NAND2X1 U13467 ( .A(n12922), .B(n7444), .Y(n12917) );
  NAND2X1 U13468 ( .A(n12927), .B(n12928), .Y(n12916) );
  ADDHXL U13469 ( .A(n11754), .B(n12929), .S(n7291) );
  AND2X1 U13470 ( .A(n11751), .B(n11753), .Y(n12929) );
  NAND2X1 U13471 ( .A(n12930), .B(n12931), .Y(n11753) );
  NAND2X1 U13472 ( .A(n9755), .B(n12727), .Y(n12931) );
  ADDHXL U13473 ( .A(n10227), .B(n12932), .S(n12930) );
  NAND3X1 U13474 ( .A(n12932), .B(n12727), .C(n9755), .Y(n11751) );
  NAND4X1 U13475 ( .A(n12933), .B(n12934), .C(n12935), .D(n12936), .Y(n12727)
         );
  NOR4X1 U13476 ( .A(n12937), .B(n12938), .C(n12939), .D(n12940), .Y(n12936)
         );
  NOR2X1 U13477 ( .A(n10663), .B(n11539), .Y(n12940) );
  NOR2X1 U13478 ( .A(n10662), .B(n11549), .Y(n12939) );
  NOR2X1 U13479 ( .A(n10654), .B(n11548), .Y(n12938) );
  NOR2X1 U13480 ( .A(n10646), .B(n11547), .Y(n12937) );
  NOR4X1 U13481 ( .A(n12941), .B(n12942), .C(n12943), .D(n12944), .Y(n12935)
         );
  NOR2X1 U13482 ( .A(n10655), .B(n11532), .Y(n12944) );
  NOR2X1 U13483 ( .A(n10649), .B(n11531), .Y(n12943) );
  NOR2X1 U13484 ( .A(n10665), .B(n11541), .Y(n12942) );
  NOR2X1 U13485 ( .A(n10664), .B(n11540), .Y(n12941) );
  NOR4X1 U13486 ( .A(n12945), .B(n12946), .C(n12947), .D(n12948), .Y(n12934)
         );
  NOR2X1 U13487 ( .A(n10647), .B(n11525), .Y(n12948) );
  NOR2X1 U13488 ( .A(n10641), .B(n11524), .Y(n12947) );
  NOR2X1 U13489 ( .A(n10640), .B(n11523), .Y(n12946) );
  NOR2X1 U13490 ( .A(n10656), .B(n11533), .Y(n12945) );
  NOR4X1 U13491 ( .A(n12949), .B(n12950), .C(n12951), .D(n12952), .Y(n12933)
         );
  NOR2X1 U13492 ( .A(n10638), .B(n11546), .Y(n12952) );
  NOR2X1 U13493 ( .A(n10639), .B(n11522), .Y(n12951) );
  NOR2X1 U13494 ( .A(n10648), .B(n11530), .Y(n12950) );
  NOR2X1 U13495 ( .A(n10657), .B(n11538), .Y(n12949) );
  NAND4X1 U13496 ( .A(n12953), .B(n12954), .C(n12955), .D(n12956), .Y(n12932)
         );
  NAND2X1 U13497 ( .A(G21610), .B(n7564), .Y(n12956) );
  NAND2X1 U13498 ( .A(G21705), .B(n10236), .Y(n12955) );
  NAND2X1 U13499 ( .A(G21737), .B(n10333), .Y(n12954) );
  NAND2X1 U13500 ( .A(G21578), .B(n10503), .Y(n12953) );
  NAND2X1 U13501 ( .A(n12738), .B(n12957), .Y(n11754) );
  NAND2X1 U13502 ( .A(n12736), .B(n12737), .Y(n12957) );
  NAND2X1 U13503 ( .A(n12958), .B(n12959), .Y(n12737) );
  NAND2X1 U13504 ( .A(n9755), .B(n12698), .Y(n12959) );
  ADDHXL U13505 ( .A(n10227), .B(n12960), .S(n12958) );
  NAND2X1 U13506 ( .A(n12896), .B(n12961), .Y(n12736) );
  NAND2X1 U13507 ( .A(n12897), .B(n12894), .Y(n12961) );
  NAND2X1 U13508 ( .A(n12888), .B(n12962), .Y(n12894) );
  NAND2X1 U13509 ( .A(n12886), .B(n12887), .Y(n12962) );
  NAND2X1 U13510 ( .A(n12963), .B(n12964), .Y(n12887) );
  NAND2X1 U13511 ( .A(n9755), .B(n12682), .Y(n12964) );
  ADDHXL U13512 ( .A(n10227), .B(n12965), .S(n12963) );
  NOR2X1 U13513 ( .A(n12753), .B(n12752), .Y(n12886) );
  ADDHXL U13514 ( .A(n12966), .B(n10227), .S(n12752) );
  NAND4X1 U13515 ( .A(n12967), .B(n12968), .C(n12969), .D(n12970), .Y(n12966)
         );
  NAND2X1 U13516 ( .A(G21606), .B(n7564), .Y(n12970) );
  NAND2X1 U13517 ( .A(G21701), .B(n10236), .Y(n12969) );
  NAND2X1 U13518 ( .A(G21733), .B(n10333), .Y(n12968) );
  NAND2X1 U13519 ( .A(G21574), .B(n10503), .Y(n12967) );
  NAND2X1 U13520 ( .A(n12880), .B(n12879), .Y(n12753) );
  ADDHXL U13521 ( .A(n12971), .B(n9260), .S(n12879) );
  NAND4X1 U13522 ( .A(n12972), .B(n12973), .C(n12974), .D(n12975), .Y(n12971)
         );
  NAND2X1 U13523 ( .A(G21605), .B(n7564), .Y(n12975) );
  NAND2X1 U13524 ( .A(G21700), .B(n10236), .Y(n12974) );
  NAND2X1 U13525 ( .A(G21732), .B(n10333), .Y(n12973) );
  NAND2X1 U13526 ( .A(G21573), .B(n10503), .Y(n12972) );
  AND2X1 U13527 ( .A(n12862), .B(n12872), .Y(n12880) );
  ADDHXL U13528 ( .A(n12976), .B(n9260), .S(n12872) );
  NAND4X1 U13529 ( .A(n12977), .B(n12978), .C(n12979), .D(n12980), .Y(n12976)
         );
  NAND2X1 U13530 ( .A(G21604), .B(n7564), .Y(n12980) );
  NAND2X1 U13531 ( .A(G21699), .B(n10236), .Y(n12979) );
  NAND2X1 U13532 ( .A(G21731), .B(n10333), .Y(n12978) );
  NAND2X1 U13533 ( .A(G21572), .B(n10503), .Y(n12977) );
  NOR3X1 U13534 ( .A(n12863), .B(n12981), .C(n12832), .Y(n12862) );
  INVX1 U13535 ( .A(n12865), .Y(n12832) );
  NOR2X1 U13536 ( .A(n12834), .B(n12833), .Y(n12865) );
  AND2X1 U13537 ( .A(n12821), .B(n12982), .Y(n12833) );
  NAND2X1 U13538 ( .A(n12820), .B(n12819), .Y(n12982) );
  NAND2X1 U13539 ( .A(n12802), .B(n12983), .Y(n12819) );
  OR2X1 U13540 ( .A(n10227), .B(n12801), .Y(n12983) );
  NOR2X1 U13541 ( .A(n12984), .B(n12985), .Y(n12801) );
  NAND2X1 U13542 ( .A(n12985), .B(n12984), .Y(n12802) );
  NAND4X1 U13543 ( .A(n10271), .B(n12986), .C(n9267), .D(n8783), .Y(n12984) );
  NAND2X1 U13544 ( .A(G21428), .B(n12987), .Y(n12986) );
  NAND4X1 U13545 ( .A(n9219), .B(n12988), .C(n12989), .D(n12990), .Y(n12987)
         );
  NOR3X1 U13546 ( .A(n12991), .B(n12992), .C(n12993), .Y(n12990) );
  NOR2X1 U13547 ( .A(n9751), .B(n12994), .Y(n12993) );
  NOR3X1 U13548 ( .A(n7446), .B(n9194), .C(n12995), .Y(n12992) );
  NOR2X1 U13549 ( .A(n7455), .B(n9751), .Y(n12995) );
  NOR2X1 U13550 ( .A(n12707), .B(n7456), .Y(n12991) );
  INVX1 U13551 ( .A(n12788), .Y(n12989) );
  NAND3X1 U13552 ( .A(n12996), .B(n12997), .C(n12998), .Y(n12788) );
  NAND2X1 U13553 ( .A(n7455), .B(n7456), .Y(n12998) );
  NAND2X1 U13554 ( .A(n9281), .B(n9076), .Y(n12996) );
  NAND2X1 U13555 ( .A(n12784), .B(n7451), .Y(n12988) );
  AND2X1 U13556 ( .A(n12999), .B(n13000), .Y(n9219) );
  NAND2X1 U13557 ( .A(n9224), .B(n7444), .Y(n13000) );
  INVX1 U13558 ( .A(n10225), .Y(n10271) );
  NAND2X1 U13559 ( .A(n8829), .B(n8804), .Y(n10225) );
  ADDHXL U13560 ( .A(n13001), .B(n9260), .S(n12985) );
  NAND4X1 U13561 ( .A(n13002), .B(n13003), .C(n13004), .D(n13005), .Y(n13001)
         );
  NOR4X1 U13562 ( .A(n13006), .B(n13007), .C(n13008), .D(n13009), .Y(n13005)
         );
  AND2X1 U13563 ( .A(n10236), .B(G21694), .Y(n13009) );
  NOR2X1 U13564 ( .A(n9085), .B(n6999), .Y(n13008) );
  INVX1 U13565 ( .A(G21599), .Y(n6999) );
  NOR2X1 U13566 ( .A(n13010), .B(n8890), .Y(n13007) );
  NOR2X1 U13567 ( .A(n8540), .B(n8783), .Y(n13006) );
  NOR2X1 U13568 ( .A(n13011), .B(n13012), .Y(n13004) );
  NOR2X1 U13569 ( .A(n9110), .B(n8804), .Y(n13012) );
  NAND2X1 U13570 ( .A(n13013), .B(n13014), .Y(n9110) );
  NAND2X1 U13571 ( .A(n9053), .B(n13015), .Y(n13014) );
  NOR2X1 U13572 ( .A(n10235), .B(n9624), .Y(n13011) );
  INVX1 U13573 ( .A(G21726), .Y(n9624) );
  NAND2X1 U13574 ( .A(G21567), .B(n10503), .Y(n13003) );
  NAND2X1 U13575 ( .A(n9084), .B(n9071), .Y(n13002) );
  NAND2X1 U13576 ( .A(n13016), .B(n13017), .Y(n12820) );
  ADDHXL U13577 ( .A(n10227), .B(n13018), .S(n13017) );
  INVX1 U13578 ( .A(n13019), .Y(n13016) );
  NAND2X1 U13579 ( .A(n13020), .B(n13019), .Y(n12821) );
  NAND4X1 U13580 ( .A(n9085), .B(n13021), .C(n9267), .D(n13022), .Y(n13019) );
  NOR2X1 U13581 ( .A(n13023), .B(n13024), .Y(n13022) );
  INVX1 U13582 ( .A(n12806), .Y(n13024) );
  NOR2X1 U13583 ( .A(n10013), .B(n13025), .Y(n12806) );
  NOR3X1 U13584 ( .A(n8817), .B(n7442), .C(n9200), .Y(n13025) );
  NOR2X1 U13585 ( .A(n9187), .B(n12810), .Y(n13023) );
  INVX1 U13586 ( .A(n13026), .Y(n12810) );
  INVX1 U13587 ( .A(n8856), .Y(n9187) );
  ADDHXL U13588 ( .A(n13018), .B(n9260), .S(n13020) );
  NAND4X1 U13589 ( .A(n13027), .B(n13028), .C(n13029), .D(n13030), .Y(n13018)
         );
  NOR4X1 U13590 ( .A(n13031), .B(n13032), .C(n13033), .D(n13034), .Y(n13030)
         );
  NOR2X1 U13591 ( .A(n9085), .B(n6988), .Y(n13034) );
  INVX1 U13592 ( .A(G21600), .Y(n6988) );
  NOR2X1 U13593 ( .A(n8880), .B(n8783), .Y(n13033) );
  NOR2X1 U13594 ( .A(n13010), .B(n10945), .Y(n13032) );
  INVX1 U13595 ( .A(n13035), .Y(n13010) );
  NOR2X1 U13596 ( .A(n8804), .B(n9132), .Y(n13031) );
  ADDFXL U13597 ( .A(n13036), .B(n13037), .CI(n13013), .S(n9132) );
  NOR2X1 U13598 ( .A(n13038), .B(n13039), .Y(n13029) );
  NOR2X1 U13599 ( .A(n10235), .B(n9614), .Y(n13039) );
  INVX1 U13600 ( .A(G21727), .Y(n9614) );
  AND2X1 U13601 ( .A(n10236), .B(G21695), .Y(n13038) );
  NAND2X1 U13602 ( .A(G21568), .B(n10503), .Y(n13028) );
  NAND2X1 U13603 ( .A(n9071), .B(n9124), .Y(n13027) );
  ADDHXL U13604 ( .A(n13040), .B(n10227), .S(n12834) );
  NAND4X1 U13605 ( .A(n13041), .B(n13042), .C(n13043), .D(n13044), .Y(n13040)
         );
  NOR4X1 U13606 ( .A(n13045), .B(n13046), .C(n13047), .D(n13048), .Y(n13044)
         );
  NOR2X1 U13607 ( .A(n9085), .B(n6978), .Y(n13048) );
  INVX1 U13608 ( .A(G21601), .Y(n6978) );
  NOR2X1 U13609 ( .A(n8800), .B(n8783), .Y(n13047) );
  NOR2X1 U13610 ( .A(n9155), .B(n8804), .Y(n13046) );
  ADDFXL U13611 ( .A(n13049), .B(n9642), .CI(n13050), .S(n9155) );
  NOR2X1 U13612 ( .A(n10235), .B(n9606), .Y(n13045) );
  INVX1 U13613 ( .A(G21728), .Y(n9606) );
  NOR2X1 U13614 ( .A(n13051), .B(n13052), .Y(n13043) );
  AND2X1 U13615 ( .A(n10236), .B(G21696), .Y(n13052) );
  NOR2X1 U13616 ( .A(n8829), .B(n9154), .Y(n13051) );
  NAND2X1 U13617 ( .A(G21569), .B(n10503), .Y(n13042) );
  NAND2X1 U13618 ( .A(G21559), .B(n13035), .Y(n13041) );
  INVX1 U13619 ( .A(n12848), .Y(n12981) );
  ADDHXL U13620 ( .A(n13053), .B(n9260), .S(n12848) );
  NAND4X1 U13621 ( .A(n13054), .B(n13055), .C(n13056), .D(n13057), .Y(n13053)
         );
  NOR4X1 U13622 ( .A(n13058), .B(n13059), .C(n13060), .D(n13061), .Y(n13057)
         );
  NOR2X1 U13623 ( .A(n9085), .B(n6968), .Y(n13061) );
  INVX1 U13624 ( .A(G21602), .Y(n6968) );
  NOR2X1 U13625 ( .A(n8799), .B(n8783), .Y(n13060) );
  INVX1 U13626 ( .A(n8798), .Y(n8783) );
  NOR2X1 U13627 ( .A(G21427), .B(G21426), .Y(n8798) );
  NOR2X1 U13628 ( .A(n9173), .B(n8804), .Y(n13059) );
  NAND2X1 U13629 ( .A(G21797), .B(G21427), .Y(n8804) );
  ADDHXL U13630 ( .A(n13062), .B(n13063), .S(n9173) );
  NOR2X1 U13631 ( .A(n13064), .B(n13065), .Y(n13063) );
  NOR2X1 U13632 ( .A(n13049), .B(n13050), .Y(n13065) );
  NOR2X1 U13633 ( .A(n13066), .B(n9642), .Y(n13064) );
  AND2X1 U13634 ( .A(n13049), .B(n13050), .Y(n13066) );
  AND2X1 U13635 ( .A(n13067), .B(n13068), .Y(n13050) );
  NAND2X1 U13636 ( .A(n13069), .B(n13070), .Y(n13068) );
  NAND2X1 U13637 ( .A(n13036), .B(n13013), .Y(n13070) );
  INVX1 U13638 ( .A(n13037), .Y(n13069) );
  OR2X1 U13639 ( .A(n13013), .B(n13036), .Y(n13067) );
  NOR2X1 U13640 ( .A(n13071), .B(n7464), .Y(n13036) );
  NOR2X1 U13641 ( .A(n9137), .B(G21426), .Y(n7464) );
  AND2X1 U13642 ( .A(G21560), .B(n13072), .Y(n13071) );
  NAND2X1 U13643 ( .A(n13073), .B(n13074), .Y(n13013) );
  NAND2X1 U13644 ( .A(n13075), .B(n13015), .Y(n13074) );
  NAND2X1 U13645 ( .A(G21561), .B(n13072), .Y(n13015) );
  NAND2X1 U13646 ( .A(n9084), .B(n7430), .Y(n13075) );
  INVX1 U13647 ( .A(n9053), .Y(n13073) );
  NOR2X1 U13648 ( .A(n8711), .B(n7430), .Y(n9053) );
  NOR2X1 U13649 ( .A(n13076), .B(n7469), .Y(n13049) );
  NOR2X1 U13650 ( .A(n9154), .B(G21426), .Y(n7469) );
  AND2X1 U13651 ( .A(G21559), .B(n13072), .Y(n13076) );
  NAND2X1 U13652 ( .A(n13077), .B(n13078), .Y(n13062) );
  NAND2X1 U13653 ( .A(G21558), .B(n13072), .Y(n13078) );
  NAND3X1 U13654 ( .A(n13037), .B(n9642), .C(n13079), .Y(n13072) );
  NAND2X1 U13655 ( .A(n9184), .B(G21426), .Y(n13079) );
  NAND2X1 U13656 ( .A(n7451), .B(G21426), .Y(n9642) );
  NAND2X1 U13657 ( .A(G21426), .B(n13080), .Y(n13037) );
  NAND2X1 U13658 ( .A(n13081), .B(n13082), .Y(n13080) );
  NAND2X1 U13659 ( .A(n9185), .B(n13083), .Y(n13081) );
  INVX1 U13660 ( .A(n10116), .Y(n13083) );
  NAND2X1 U13661 ( .A(n7473), .B(n7430), .Y(n13077) );
  NOR2X1 U13662 ( .A(n10235), .B(n9598), .Y(n13058) );
  INVX1 U13663 ( .A(G21729), .Y(n9598) );
  INVX1 U13664 ( .A(n10333), .Y(n10235) );
  NOR2X1 U13665 ( .A(n13084), .B(n13085), .Y(n13056) );
  AND2X1 U13666 ( .A(n10236), .B(G21697), .Y(n13085) );
  NOR2X1 U13667 ( .A(n8829), .B(n9171), .Y(n13084) );
  INVX1 U13668 ( .A(n9071), .Y(n8829) );
  NAND2X1 U13669 ( .A(G21570), .B(n10503), .Y(n13055) );
  NAND2X1 U13670 ( .A(G21558), .B(n13035), .Y(n13054) );
  NAND3X1 U13671 ( .A(n9267), .B(n12811), .C(n12903), .Y(n13035) );
  AND2X1 U13672 ( .A(n13086), .B(n13087), .Y(n12903) );
  NAND2X1 U13673 ( .A(n13026), .B(n8856), .Y(n13087) );
  NOR4X1 U13674 ( .A(n9632), .B(n11987), .C(n12809), .D(n7458), .Y(n8856) );
  NAND2X1 U13675 ( .A(n7455), .B(n8711), .Y(n11987) );
  NAND2X1 U13676 ( .A(G21428), .B(n13088), .Y(n13086) );
  NAND4X1 U13677 ( .A(n13089), .B(n13090), .C(n13091), .D(n13092), .Y(n13088)
         );
  NOR4X1 U13678 ( .A(n7418), .B(n13093), .C(n13094), .D(n13095), .Y(n13092) );
  NOR2X1 U13679 ( .A(n9077), .B(n9193), .Y(n13095) );
  NOR2X1 U13680 ( .A(n9185), .B(n13096), .Y(n9077) );
  NOR2X1 U13681 ( .A(n7444), .B(n9076), .Y(n13096) );
  NOR2X1 U13682 ( .A(n13097), .B(n9278), .Y(n13094) );
  INVX1 U13683 ( .A(n9224), .Y(n9278) );
  NOR2X1 U13684 ( .A(n8711), .B(n7456), .Y(n9224) );
  NOR2X1 U13685 ( .A(n13098), .B(n9281), .Y(n13097) );
  NOR2X1 U13686 ( .A(n7442), .B(n12906), .Y(n13098) );
  NOR3X1 U13687 ( .A(n12787), .B(n9076), .C(n12784), .Y(n13093) );
  INVX1 U13688 ( .A(n9194), .Y(n12787) );
  NOR2X1 U13689 ( .A(n9200), .B(n7458), .Y(n7418) );
  NOR2X1 U13690 ( .A(n13099), .B(n9186), .Y(n13091) );
  NAND4X1 U13691 ( .A(n13100), .B(n13101), .C(n13102), .D(n13103), .Y(n9186)
         );
  NAND2X1 U13692 ( .A(n12784), .B(n13104), .Y(n13103) );
  NAND3X1 U13693 ( .A(n7446), .B(n12906), .C(n9751), .Y(n13104) );
  NAND3X1 U13694 ( .A(n7442), .B(n7456), .C(n8782), .Y(n13102) );
  NAND2X1 U13695 ( .A(n9194), .B(n9193), .Y(n13101) );
  INVX1 U13696 ( .A(n12789), .Y(n13100) );
  NAND3X1 U13697 ( .A(n13105), .B(n12999), .C(n13106), .Y(n12789) );
  NAND2X1 U13698 ( .A(n13107), .B(n8762), .Y(n13106) );
  NAND2X1 U13699 ( .A(n9218), .B(n9223), .Y(n13107) );
  NAND2X1 U13700 ( .A(n11808), .B(n7451), .Y(n12999) );
  NAND2X1 U13701 ( .A(n13108), .B(n8743), .Y(n13105) );
  NAND2X1 U13702 ( .A(n7439), .B(n13109), .Y(n13108) );
  NAND2X1 U13703 ( .A(n7455), .B(n7458), .Y(n13109) );
  NOR2X1 U13704 ( .A(n7455), .B(n12997), .Y(n13099) );
  INVX1 U13705 ( .A(n9184), .Y(n12997) );
  NOR2X1 U13706 ( .A(n8743), .B(n9076), .Y(n9184) );
  NAND2X1 U13707 ( .A(n9631), .B(n13082), .Y(n13090) );
  OR2X1 U13708 ( .A(n9192), .B(n9179), .Y(n13089) );
  NAND3X1 U13709 ( .A(G21428), .B(n7457), .C(n8861), .Y(n12811) );
  INVX1 U13710 ( .A(n10014), .Y(n9267) );
  NOR2X1 U13711 ( .A(n9134), .B(n8817), .Y(n10014) );
  NAND4X1 U13712 ( .A(n10256), .B(n12994), .C(n9059), .D(n7458), .Y(n9134) );
  NOR3X1 U13713 ( .A(n7456), .B(n12784), .C(n8772), .Y(n12994) );
  NOR2X1 U13714 ( .A(n8711), .B(n9751), .Y(n10256) );
  ADDHXL U13715 ( .A(n13110), .B(n10227), .S(n12863) );
  NAND4X1 U13716 ( .A(n13111), .B(n13112), .C(n13113), .D(n13114), .Y(n13110)
         );
  NAND2X1 U13717 ( .A(G21603), .B(n7564), .Y(n13114) );
  NAND2X1 U13718 ( .A(G21698), .B(n10236), .Y(n13113) );
  NAND2X1 U13719 ( .A(G21730), .B(n10333), .Y(n13112) );
  NAND2X1 U13720 ( .A(G21571), .B(n10503), .Y(n13111) );
  NAND3X1 U13721 ( .A(n12965), .B(n12682), .C(n9755), .Y(n12888) );
  NAND4X1 U13722 ( .A(n13115), .B(n13116), .C(n13117), .D(n13118), .Y(n12682)
         );
  NOR4X1 U13723 ( .A(n13119), .B(n13120), .C(n13121), .D(n13122), .Y(n13118)
         );
  NOR2X1 U13724 ( .A(n10940), .B(n11539), .Y(n13122) );
  NOR2X1 U13725 ( .A(n10939), .B(n11549), .Y(n13121) );
  NOR2X1 U13726 ( .A(n10927), .B(n11548), .Y(n13120) );
  NOR2X1 U13727 ( .A(n10916), .B(n11547), .Y(n13119) );
  NOR4X1 U13728 ( .A(n13123), .B(n13124), .C(n13125), .D(n13126), .Y(n13117)
         );
  NOR2X1 U13729 ( .A(n10929), .B(n11532), .Y(n13126) );
  NOR2X1 U13730 ( .A(n10922), .B(n11531), .Y(n13125) );
  NOR2X1 U13731 ( .A(n10942), .B(n11541), .Y(n13124) );
  NOR2X1 U13732 ( .A(n10941), .B(n11540), .Y(n13123) );
  NOR4X1 U13733 ( .A(n13127), .B(n13128), .C(n13129), .D(n13130), .Y(n13116)
         );
  NOR2X1 U13734 ( .A(n10918), .B(n11525), .Y(n13130) );
  NOR2X1 U13735 ( .A(n10911), .B(n11524), .Y(n13129) );
  NOR2X1 U13736 ( .A(n10909), .B(n11523), .Y(n13128) );
  NOR2X1 U13737 ( .A(n10931), .B(n11533), .Y(n13127) );
  NOR4X1 U13738 ( .A(n13131), .B(n13132), .C(n13133), .D(n13134), .Y(n13115)
         );
  NOR2X1 U13739 ( .A(n10904), .B(n11546), .Y(n13134) );
  NOR2X1 U13740 ( .A(n10907), .B(n11522), .Y(n13133) );
  NOR2X1 U13741 ( .A(n10919), .B(n11530), .Y(n13132) );
  NOR2X1 U13742 ( .A(n10932), .B(n11538), .Y(n13131) );
  NAND4X1 U13743 ( .A(n13135), .B(n13136), .C(n13137), .D(n13138), .Y(n12965)
         );
  NAND2X1 U13744 ( .A(G21607), .B(n7564), .Y(n13138) );
  NAND2X1 U13745 ( .A(G21702), .B(n10236), .Y(n13137) );
  NAND2X1 U13746 ( .A(G21734), .B(n10333), .Y(n13136) );
  NAND2X1 U13747 ( .A(G21575), .B(n10503), .Y(n13135) );
  NAND2X1 U13748 ( .A(n13139), .B(n13140), .Y(n12897) );
  NAND2X1 U13749 ( .A(n9755), .B(n12690), .Y(n13140) );
  ADDHXL U13750 ( .A(n10227), .B(n13141), .S(n13139) );
  NAND3X1 U13751 ( .A(n13141), .B(n12690), .C(n9755), .Y(n12896) );
  NAND4X1 U13752 ( .A(n13142), .B(n13143), .C(n13144), .D(n13145), .Y(n12690)
         );
  NOR4X1 U13753 ( .A(n13146), .B(n13147), .C(n13148), .D(n13149), .Y(n13145)
         );
  NOR2X1 U13754 ( .A(n10842), .B(n11539), .Y(n13149) );
  NOR2X1 U13755 ( .A(n10841), .B(n11549), .Y(n13148) );
  NOR2X1 U13756 ( .A(n10833), .B(n11548), .Y(n13147) );
  NOR2X1 U13757 ( .A(n10825), .B(n11547), .Y(n13146) );
  NOR4X1 U13758 ( .A(n13150), .B(n13151), .C(n13152), .D(n13153), .Y(n13144)
         );
  NOR2X1 U13759 ( .A(n10834), .B(n11532), .Y(n13153) );
  NOR2X1 U13760 ( .A(n10828), .B(n11531), .Y(n13152) );
  NOR2X1 U13761 ( .A(n10844), .B(n11541), .Y(n13151) );
  NOR2X1 U13762 ( .A(n10843), .B(n11540), .Y(n13150) );
  NOR4X1 U13763 ( .A(n13154), .B(n13155), .C(n13156), .D(n13157), .Y(n13143)
         );
  NOR2X1 U13764 ( .A(n10826), .B(n11525), .Y(n13157) );
  NOR2X1 U13765 ( .A(n10820), .B(n11524), .Y(n13156) );
  NOR2X1 U13766 ( .A(n10819), .B(n11523), .Y(n13155) );
  NOR2X1 U13767 ( .A(n10835), .B(n11533), .Y(n13154) );
  NOR4X1 U13768 ( .A(n13158), .B(n13159), .C(n13160), .D(n13161), .Y(n13142)
         );
  NOR2X1 U13769 ( .A(n10817), .B(n11546), .Y(n13161) );
  NOR2X1 U13770 ( .A(n10818), .B(n11522), .Y(n13160) );
  NOR2X1 U13771 ( .A(n10827), .B(n11530), .Y(n13159) );
  NOR2X1 U13772 ( .A(n10836), .B(n11538), .Y(n13158) );
  NAND4X1 U13773 ( .A(n13162), .B(n13163), .C(n13164), .D(n13165), .Y(n13141)
         );
  NAND2X1 U13774 ( .A(G21608), .B(n7564), .Y(n13165) );
  NAND2X1 U13775 ( .A(G21703), .B(n10236), .Y(n13164) );
  NAND2X1 U13776 ( .A(G21735), .B(n10333), .Y(n13163) );
  NAND2X1 U13777 ( .A(G21576), .B(n10503), .Y(n13162) );
  NAND3X1 U13778 ( .A(n12960), .B(n12698), .C(n9755), .Y(n12738) );
  INVX1 U13779 ( .A(n9138), .Y(n7428) );
  NOR4X1 U13780 ( .A(n12809), .B(n13166), .C(n12060), .D(n7455), .Y(n9138) );
  INVX1 U13781 ( .A(n11808), .Y(n12060) );
  NOR2X1 U13782 ( .A(n7446), .B(n9076), .Y(n11808) );
  NAND4X1 U13783 ( .A(n13167), .B(n13168), .C(n13169), .D(n13170), .Y(n12698)
         );
  NOR4X1 U13784 ( .A(n13171), .B(n13172), .C(n13173), .D(n13174), .Y(n13170)
         );
  NOR2X1 U13785 ( .A(n10752), .B(n11539), .Y(n13174) );
  NAND2X1 U13786 ( .A(n13175), .B(n10952), .Y(n11539) );
  NOR2X1 U13787 ( .A(n10751), .B(n11549), .Y(n13173) );
  NAND2X1 U13788 ( .A(n13175), .B(n10944), .Y(n11549) );
  NOR2X1 U13789 ( .A(n10743), .B(n11548), .Y(n13172) );
  NAND2X1 U13790 ( .A(n13176), .B(n10944), .Y(n11548) );
  NOR2X1 U13791 ( .A(n10735), .B(n11547), .Y(n13171) );
  NAND2X1 U13792 ( .A(n13177), .B(n9135), .Y(n11547) );
  NOR4X1 U13793 ( .A(n13178), .B(n13179), .C(n13180), .D(n13181), .Y(n13169)
         );
  NOR2X1 U13794 ( .A(n10744), .B(n11532), .Y(n13181) );
  NAND2X1 U13795 ( .A(n13176), .B(n10952), .Y(n11532) );
  NOR2X1 U13796 ( .A(n10738), .B(n11531), .Y(n13180) );
  NAND2X1 U13797 ( .A(n13177), .B(n10944), .Y(n11531) );
  NOR2X1 U13798 ( .A(n10754), .B(n11541), .Y(n13179) );
  NAND2X1 U13799 ( .A(n13175), .B(n9135), .Y(n11541) );
  NOR2X1 U13800 ( .A(n10753), .B(n11540), .Y(n13178) );
  NAND2X1 U13801 ( .A(n13175), .B(n8889), .Y(n11540) );
  AND2X1 U13802 ( .A(n13182), .B(n13183), .Y(n13175) );
  NOR4X1 U13803 ( .A(n13184), .B(n13185), .C(n13186), .D(n13187), .Y(n13168)
         );
  NOR2X1 U13804 ( .A(n10736), .B(n11525), .Y(n13187) );
  NAND2X1 U13805 ( .A(n13177), .B(n8889), .Y(n11525) );
  NOR2X1 U13806 ( .A(n10730), .B(n11524), .Y(n13186) );
  NAND2X1 U13807 ( .A(n13188), .B(n10944), .Y(n11524) );
  NOR2X1 U13808 ( .A(n10729), .B(n11523), .Y(n13185) );
  NAND2X1 U13809 ( .A(n13188), .B(n10952), .Y(n11523) );
  NOR2X1 U13810 ( .A(n10745), .B(n11533), .Y(n13184) );
  NAND2X1 U13811 ( .A(n13176), .B(n8889), .Y(n11533) );
  NOR4X1 U13812 ( .A(n13189), .B(n13190), .C(n13191), .D(n13192), .Y(n13167)
         );
  NOR2X1 U13813 ( .A(n10727), .B(n11546), .Y(n13192) );
  NAND2X1 U13814 ( .A(n13188), .B(n9135), .Y(n11546) );
  NOR2X1 U13815 ( .A(n10728), .B(n11522), .Y(n13191) );
  NAND2X1 U13816 ( .A(n13188), .B(n8889), .Y(n11522) );
  AND2X1 U13817 ( .A(n13183), .B(n13193), .Y(n13188) );
  NOR2X1 U13818 ( .A(n10737), .B(n11530), .Y(n13190) );
  NAND2X1 U13819 ( .A(n13177), .B(n10952), .Y(n11530) );
  NOR2X1 U13820 ( .A(n13183), .B(n13182), .Y(n13177) );
  INVX1 U13821 ( .A(n13193), .Y(n13182) );
  NOR2X1 U13822 ( .A(n10746), .B(n11538), .Y(n13189) );
  NAND2X1 U13823 ( .A(n13176), .B(n9135), .Y(n11538) );
  NOR2X1 U13824 ( .A(n13193), .B(n13183), .Y(n13176) );
  ADDHXL U13825 ( .A(n10945), .B(n8893), .S(n13183) );
  NAND3X1 U13826 ( .A(n13194), .B(n13195), .C(n13196), .Y(n13193) );
  INVX1 U13827 ( .A(n13197), .Y(n13196) );
  NAND2X1 U13828 ( .A(G21558), .B(n10945), .Y(n13195) );
  NAND2X1 U13829 ( .A(n13198), .B(G21560), .Y(n13194) );
  NAND4X1 U13830 ( .A(n13199), .B(n13200), .C(n13201), .D(n13202), .Y(n12960)
         );
  NAND2X1 U13831 ( .A(G21609), .B(n7564), .Y(n13202) );
  NAND2X1 U13832 ( .A(G21704), .B(n10236), .Y(n13201) );
  NOR2X1 U13833 ( .A(n7426), .B(n8817), .Y(n10236) );
  NAND4X1 U13834 ( .A(n13203), .B(n9194), .C(n9076), .D(n7451), .Y(n7426) );
  NOR2X1 U13835 ( .A(n7442), .B(n8762), .Y(n9194) );
  NAND2X1 U13836 ( .A(G21736), .B(n10333), .Y(n13200) );
  NAND2X1 U13837 ( .A(n10227), .B(n9753), .Y(n10333) );
  NAND2X1 U13838 ( .A(n9174), .B(G21428), .Y(n9753) );
  INVX1 U13839 ( .A(n12907), .Y(n9174) );
  NAND4X1 U13840 ( .A(n13203), .B(n9195), .C(n8772), .D(n8711), .Y(n12907) );
  NOR3X1 U13841 ( .A(n8782), .B(n7458), .C(n9193), .Y(n13203) );
  INVX1 U13842 ( .A(n9212), .Y(n7429) );
  NOR4X1 U13843 ( .A(n9223), .B(n12809), .C(n12708), .D(n9076), .Y(n9212) );
  NAND3X1 U13844 ( .A(n8743), .B(n8782), .C(n7439), .Y(n12809) );
  INVX1 U13845 ( .A(n9281), .Y(n9223) );
  NOR2X1 U13846 ( .A(n8772), .B(n7458), .Y(n9281) );
  NAND2X1 U13847 ( .A(G21577), .B(n10503), .Y(n13199) );
  NAND3X1 U13848 ( .A(n13021), .B(n12843), .C(n13204), .Y(n10503) );
  NAND2X1 U13849 ( .A(G21428), .B(n13205), .Y(n13204) );
  NAND3X1 U13850 ( .A(n13206), .B(n12911), .C(n12846), .Y(n13205) );
  AND2X1 U13851 ( .A(n13207), .B(n13208), .Y(n12846) );
  NAND3X1 U13852 ( .A(n13209), .B(n7458), .C(n9202), .Y(n13208) );
  NAND2X1 U13853 ( .A(n13210), .B(n9632), .Y(n13209) );
  INVX1 U13854 ( .A(n9203), .Y(n9632) );
  NAND2X1 U13855 ( .A(n7442), .B(n9059), .Y(n13210) );
  OR2X1 U13856 ( .A(n9218), .B(n9200), .Y(n13207) );
  NAND3X1 U13857 ( .A(n7451), .B(n7455), .C(n9202), .Y(n9200) );
  NOR3X1 U13858 ( .A(n8711), .B(n12784), .C(n9193), .Y(n9202) );
  NAND2X1 U13859 ( .A(n9751), .B(n7439), .Y(n9193) );
  NAND2X1 U13860 ( .A(n7458), .B(n8772), .Y(n9218) );
  NAND4X1 U13861 ( .A(n12784), .B(n9751), .C(n9203), .D(n13211), .Y(n12911) );
  NOR3X1 U13862 ( .A(n7458), .B(n7439), .C(n8762), .Y(n13211) );
  NOR2X1 U13863 ( .A(n8772), .B(n7444), .Y(n9203) );
  NAND2X1 U13864 ( .A(n9092), .B(n8861), .Y(n13206) );
  NOR2X1 U13865 ( .A(n9179), .B(n13082), .Y(n8861) );
  NAND2X1 U13866 ( .A(n8711), .B(n8743), .Y(n13082) );
  NAND2X1 U13867 ( .A(n13212), .B(n7439), .Y(n9179) );
  INVX1 U13868 ( .A(n7457), .Y(n9092) );
  NAND2X1 U13869 ( .A(n13213), .B(n13214), .Y(n7457) );
  NAND3X1 U13870 ( .A(n13215), .B(n12673), .C(n13216), .Y(n13214) );
  INVX1 U13871 ( .A(n13217), .Y(n13215) );
  NAND2X1 U13872 ( .A(n13218), .B(n13219), .Y(n13213) );
  NAND3X1 U13873 ( .A(n13220), .B(n13221), .C(n13222), .Y(n13219) );
  OR2X1 U13874 ( .A(n13217), .B(n13223), .Y(n13222) );
  NAND2X1 U13875 ( .A(n13224), .B(n13217), .Y(n13221) );
  NAND2X1 U13876 ( .A(n13225), .B(n13226), .Y(n13224) );
  NAND3X1 U13877 ( .A(n12927), .B(n12928), .C(n13227), .Y(n13226) );
  NAND2X1 U13878 ( .A(n13228), .B(n13229), .Y(n12928) );
  ADDHXL U13879 ( .A(n7474), .B(n8848), .S(n13228) );
  NAND2X1 U13880 ( .A(n13230), .B(n13231), .Y(n12927) );
  ADDHXL U13881 ( .A(G21562), .B(n8848), .S(n13230) );
  NAND2X1 U13882 ( .A(n13232), .B(n13233), .Y(n13225) );
  NAND4X1 U13883 ( .A(n13234), .B(n13235), .C(n13236), .D(n13237), .Y(n13233)
         );
  NAND2X1 U13884 ( .A(n13238), .B(n13239), .Y(n13237) );
  NAND2X1 U13885 ( .A(n8827), .B(n13240), .Y(n13238) );
  NAND3X1 U13886 ( .A(n13241), .B(n13242), .C(n13243), .Y(n13236) );
  NAND2X1 U13887 ( .A(n13244), .B(n13245), .Y(n13243) );
  NAND3X1 U13888 ( .A(n7442), .B(n13246), .C(n8827), .Y(n13245) );
  INVX1 U13889 ( .A(n13247), .Y(n13244) );
  NAND3X1 U13890 ( .A(n8827), .B(n13240), .C(n13248), .Y(n13242) );
  INVX1 U13891 ( .A(n13239), .Y(n13248) );
  NAND4X1 U13892 ( .A(n13249), .B(n13250), .C(n13217), .D(n9070), .Y(n13239)
         );
  INVX1 U13893 ( .A(G21425), .Y(n9070) );
  NAND2X1 U13894 ( .A(G21427), .B(n13251), .Y(n13250) );
  NAND2X1 U13895 ( .A(G21559), .B(n13252), .Y(n13251) );
  NAND2X1 U13896 ( .A(n13227), .B(n12922), .Y(n13249) );
  ADDFXL U13897 ( .A(G21564), .B(n8893), .CI(n13253), .S(n12922) );
  NAND2X1 U13898 ( .A(n13166), .B(n13254), .Y(n13240) );
  NAND4X1 U13899 ( .A(n13255), .B(n13256), .C(n13257), .D(n13258), .Y(n13241)
         );
  NAND2X1 U13900 ( .A(G21427), .B(n8890), .Y(n13258) );
  NAND3X1 U13901 ( .A(n13254), .B(n13166), .C(n9093), .Y(n13257) );
  NAND2X1 U13902 ( .A(n7442), .B(n8762), .Y(n13254) );
  NAND3X1 U13903 ( .A(n13246), .B(n13247), .C(n8827), .Y(n13256) );
  NAND2X1 U13904 ( .A(n13259), .B(n13260), .Y(n13247) );
  NAND3X1 U13905 ( .A(n13261), .B(n13262), .C(G21427), .Y(n13260) );
  NAND2X1 U13906 ( .A(G21560), .B(n13252), .Y(n13262) );
  NAND3X1 U13907 ( .A(G21567), .B(n9124), .C(G21795), .Y(n13261) );
  NAND2X1 U13908 ( .A(n13227), .B(n12926), .Y(n13259) );
  NAND3X1 U13909 ( .A(n13263), .B(n13264), .C(n13265), .Y(n12926) );
  OR2X1 U13910 ( .A(n8887), .B(n13266), .Y(n13265) );
  NAND3X1 U13911 ( .A(n13266), .B(G21560), .C(G21565), .Y(n13264) );
  INVX1 U13912 ( .A(n13267), .Y(n13266) );
  NAND2X1 U13913 ( .A(n13268), .B(n8880), .Y(n13263) );
  ADDHXL U13914 ( .A(n10945), .B(n13267), .S(n13268) );
  NAND2X1 U13915 ( .A(n12906), .B(n13269), .Y(n13246) );
  NAND2X1 U13916 ( .A(n8743), .B(n8762), .Y(n13269) );
  INVX1 U13917 ( .A(n9059), .Y(n12906) );
  NOR2X1 U13918 ( .A(n7444), .B(n7455), .Y(n9059) );
  NAND2X1 U13919 ( .A(n13227), .B(n12925), .Y(n13255) );
  NAND2X1 U13920 ( .A(n13267), .B(n13270), .Y(n12925) );
  NAND2X1 U13921 ( .A(G21566), .B(n8890), .Y(n13270) );
  NAND2X1 U13922 ( .A(G21427), .B(n8870), .Y(n13235) );
  NAND2X1 U13923 ( .A(n13271), .B(n13227), .Y(n13234) );
  INVX1 U13924 ( .A(n12915), .Y(n13271) );
  ADDFXL U13925 ( .A(G21563), .B(n8870), .CI(n13272), .S(n12915) );
  NAND2X1 U13926 ( .A(G21425), .B(G21557), .Y(n13232) );
  OR2X1 U13927 ( .A(n12673), .B(n13217), .Y(n13220) );
  NAND3X1 U13928 ( .A(n8743), .B(n8772), .C(n8827), .Y(n13217) );
  NAND4X1 U13929 ( .A(n13273), .B(n13274), .C(n13275), .D(n13276), .Y(n12673)
         );
  NOR4X1 U13930 ( .A(n13277), .B(n13278), .C(n13279), .D(n13280), .Y(n13276)
         );
  NOR2X1 U13931 ( .A(n10312), .B(n8688), .Y(n13280) );
  NAND2X1 U13932 ( .A(n13281), .B(n13282), .Y(n8688) );
  NOR2X1 U13933 ( .A(n10314), .B(n8610), .Y(n13279) );
  NAND2X1 U13934 ( .A(n13283), .B(n13281), .Y(n8610) );
  NOR2X1 U13935 ( .A(n10316), .B(n8528), .Y(n13278) );
  NAND2X1 U13936 ( .A(n13281), .B(n13284), .Y(n8528) );
  NOR2X1 U13937 ( .A(n10324), .B(n8371), .Y(n13277) );
  NAND2X1 U13938 ( .A(n13285), .B(n13282), .Y(n8371) );
  NOR4X1 U13939 ( .A(n13286), .B(n13287), .C(n13288), .D(n13289), .Y(n13275)
         );
  NOR2X1 U13940 ( .A(n10326), .B(n8293), .Y(n13289) );
  NAND2X1 U13941 ( .A(n13283), .B(n13285), .Y(n8293) );
  NOR2X1 U13942 ( .A(n10328), .B(n8213), .Y(n13288) );
  NAND2X1 U13943 ( .A(n13284), .B(n13285), .Y(n8213) );
  NOR2X1 U13944 ( .A(n10972), .B(n8056), .Y(n13287) );
  NAND2X1 U13945 ( .A(n13290), .B(n13282), .Y(n8056) );
  NOR2X1 U13946 ( .A(n10967), .B(n7978), .Y(n13286) );
  NAND2X1 U13947 ( .A(n13290), .B(n13283), .Y(n7978) );
  NOR4X1 U13948 ( .A(n13291), .B(n13292), .C(n13293), .D(n13294), .Y(n13274)
         );
  NOR2X1 U13949 ( .A(n10983), .B(n7898), .Y(n13294) );
  NAND2X1 U13950 ( .A(n13290), .B(n13284), .Y(n7898) );
  NOR2X1 U13951 ( .A(n10965), .B(n7736), .Y(n13293) );
  NAND2X1 U13952 ( .A(n13295), .B(n13282), .Y(n7736) );
  NOR2X1 U13953 ( .A(n9137), .B(n9084), .Y(n13282) );
  NOR2X1 U13954 ( .A(n10964), .B(n7656), .Y(n13292) );
  NAND2X1 U13955 ( .A(n13295), .B(n13283), .Y(n7656) );
  NOR2X1 U13956 ( .A(n9112), .B(n9124), .Y(n13283) );
  NOR2X1 U13957 ( .A(n10982), .B(n7570), .Y(n13291) );
  NAND2X1 U13958 ( .A(n13295), .B(n13284), .Y(n7570) );
  NOR2X1 U13959 ( .A(n9124), .B(n9084), .Y(n13284) );
  INVX1 U13960 ( .A(n9112), .Y(n9084) );
  NOR4X1 U13961 ( .A(n13296), .B(n13297), .C(n13298), .D(n13299), .Y(n13273)
         );
  NOR2X1 U13962 ( .A(n10310), .B(n8803), .Y(n13299) );
  NAND2X1 U13963 ( .A(n13300), .B(n13281), .Y(n8803) );
  NOR2X1 U13964 ( .A(n9154), .B(n9171), .Y(n13281) );
  NOR2X1 U13965 ( .A(n10322), .B(n8449), .Y(n13298) );
  NAND2X1 U13966 ( .A(n13300), .B(n13285), .Y(n8449) );
  NOR2X1 U13967 ( .A(n9171), .B(n9146), .Y(n13285) );
  NOR2X1 U13968 ( .A(n10973), .B(n8134), .Y(n13297) );
  NAND2X1 U13969 ( .A(n13300), .B(n13290), .Y(n8134) );
  NOR2X1 U13970 ( .A(n9154), .B(n7473), .Y(n13290) );
  NOR2X1 U13971 ( .A(n10966), .B(n7816), .Y(n13296) );
  NAND2X1 U13972 ( .A(n13300), .B(n13295), .Y(n7816) );
  NOR2X1 U13973 ( .A(n7473), .B(n9146), .Y(n13295) );
  INVX1 U13974 ( .A(n9154), .Y(n9146) );
  NAND2X1 U13975 ( .A(n13301), .B(n13302), .Y(n9154) );
  NAND2X1 U13976 ( .A(n13303), .B(n13304), .Y(n13302) );
  INVX1 U13977 ( .A(n9171), .Y(n7473) );
  ADDHXL U13978 ( .A(n13305), .B(n13301), .S(n9171) );
  OR2X1 U13979 ( .A(n13304), .B(n13303), .Y(n13301) );
  AND3X1 U13980 ( .A(n13306), .B(n13307), .C(n13308), .Y(n13303) );
  NAND2X1 U13981 ( .A(n9646), .B(G21559), .Y(n13308) );
  NAND2X1 U13982 ( .A(n7828), .B(n7430), .Y(n13307) );
  ADDHXL U13983 ( .A(n7824), .B(G21564), .S(n7828) );
  NAND2X1 U13984 ( .A(n9071), .B(G21564), .Y(n13306) );
  NAND2X1 U13985 ( .A(n13309), .B(n13310), .Y(n13304) );
  NAND2X1 U13986 ( .A(n13311), .B(n13312), .Y(n13310) );
  NAND2X1 U13987 ( .A(n13313), .B(n13314), .Y(n13312) );
  OR2X1 U13988 ( .A(n13314), .B(n13313), .Y(n13309) );
  INVX1 U13989 ( .A(n13315), .Y(n13313) );
  NAND3X1 U13990 ( .A(n13316), .B(n13317), .C(n13318), .Y(n13305) );
  NAND2X1 U13991 ( .A(n9646), .B(G21558), .Y(n13318) );
  NAND2X1 U13992 ( .A(n7827), .B(n7430), .Y(n13317) );
  INVX1 U13993 ( .A(n8458), .Y(n7827) );
  NOR3X1 U13994 ( .A(n8221), .B(n8137), .C(n13319), .Y(n8458) );
  NOR2X1 U13995 ( .A(n8799), .B(n7824), .Y(n13319) );
  INVX1 U13996 ( .A(n8073), .Y(n8137) );
  NAND2X1 U13997 ( .A(n7906), .B(n7824), .Y(n8073) );
  NOR2X1 U13998 ( .A(n8540), .B(n8880), .Y(n7824) );
  NOR2X1 U13999 ( .A(n8800), .B(G21563), .Y(n7906) );
  NOR2X1 U14000 ( .A(n8799), .B(G21564), .Y(n8221) );
  NAND2X1 U14001 ( .A(n9071), .B(G21563), .Y(n13316) );
  NOR2X1 U14002 ( .A(n9112), .B(n9137), .Y(n13300) );
  INVX1 U14003 ( .A(n9124), .Y(n9137) );
  ADDFXL U14004 ( .A(n13315), .B(n13311), .CI(n13314), .S(n9124) );
  NAND2X1 U14005 ( .A(n13320), .B(n13321), .Y(n13314) );
  NAND2X1 U14006 ( .A(n8815), .B(n13322), .Y(n13321) );
  ADDHXL U14007 ( .A(G21568), .B(n13323), .S(n13322) );
  NOR2X1 U14008 ( .A(n11440), .B(n9629), .Y(n13323) );
  NAND2X1 U14009 ( .A(n13324), .B(n13325), .Y(n9629) );
  NAND2X1 U14010 ( .A(G21427), .B(n7014), .Y(n13325) );
  INVX1 U14011 ( .A(G21598), .Y(n7014) );
  NAND2X1 U14012 ( .A(n9093), .B(n9320), .Y(n13324) );
  INVX1 U14013 ( .A(G21757), .Y(n9320) );
  NAND2X1 U14014 ( .A(n9195), .B(n9646), .Y(n13320) );
  AND3X1 U14015 ( .A(n13326), .B(n13327), .C(n13328), .Y(n13311) );
  NAND2X1 U14016 ( .A(n9646), .B(G21560), .Y(n13328) );
  NAND2X1 U14017 ( .A(n8539), .B(n7430), .Y(n13327) );
  INVX1 U14018 ( .A(n8697), .Y(n8539) );
  NOR2X1 U14019 ( .A(n7664), .B(n7744), .Y(n8697) );
  NOR2X1 U14020 ( .A(n8880), .B(G21566), .Y(n7744) );
  NOR2X1 U14021 ( .A(n8540), .B(G21565), .Y(n7664) );
  NAND2X1 U14022 ( .A(n9071), .B(G21565), .Y(n13326) );
  NAND2X1 U14023 ( .A(n13329), .B(n13315), .Y(n9112) );
  NAND2X1 U14024 ( .A(n13330), .B(n13331), .Y(n13315) );
  OR2X1 U14025 ( .A(n13331), .B(n13330), .Y(n13329) );
  NAND4X1 U14026 ( .A(n13332), .B(n8897), .C(n13333), .D(n13334), .Y(n13330)
         );
  NAND2X1 U14027 ( .A(n7430), .B(n8540), .Y(n13334) );
  NAND2X1 U14028 ( .A(n9071), .B(G21566), .Y(n13333) );
  NOR2X1 U14029 ( .A(n7430), .B(G21428), .Y(n9071) );
  NAND2X1 U14030 ( .A(n9646), .B(G21561), .Y(n13332) );
  NOR2X1 U14031 ( .A(n8817), .B(G21427), .Y(n9646) );
  OR3X1 U14032 ( .A(n13335), .B(n9123), .C(n8817), .Y(n13331) );
  NOR2X1 U14033 ( .A(n11440), .B(n9093), .Y(n9123) );
  INVX1 U14034 ( .A(G21567), .Y(n11440) );
  AND2X1 U14035 ( .A(n8897), .B(n13336), .Y(n13335) );
  NAND2X1 U14036 ( .A(n9060), .B(G21426), .Y(n13336) );
  NOR3X1 U14037 ( .A(n7456), .B(n9076), .C(n12708), .Y(n9060) );
  INVX1 U14038 ( .A(n9195), .Y(n12708) );
  NOR2X1 U14039 ( .A(n8762), .B(n7451), .Y(n9195) );
  INVX1 U14040 ( .A(n8815), .Y(n8897) );
  NOR2X1 U14041 ( .A(n9093), .B(n7430), .Y(n8815) );
  INVX1 U14042 ( .A(G21426), .Y(n7430) );
  INVX1 U14043 ( .A(G21427), .Y(n9093) );
  INVX1 U14044 ( .A(n13216), .Y(n13218) );
  NAND2X1 U14045 ( .A(n13337), .B(n13338), .Y(n13216) );
  NAND3X1 U14046 ( .A(G21427), .B(n13252), .C(G21557), .Y(n13338) );
  INVX1 U14047 ( .A(G21795), .Y(n13252) );
  NAND2X1 U14048 ( .A(n13227), .B(n12913), .Y(n13337) );
  NAND2X1 U14049 ( .A(n13339), .B(n13340), .Y(n12913) );
  NAND2X1 U14050 ( .A(n13341), .B(n7474), .Y(n13340) );
  INVX1 U14051 ( .A(G21562), .Y(n7474) );
  NAND2X1 U14052 ( .A(n13231), .B(n8848), .Y(n13341) );
  INVX1 U14053 ( .A(G21557), .Y(n8848) );
  INVX1 U14054 ( .A(n13229), .Y(n13231) );
  NAND2X1 U14055 ( .A(G21557), .B(n13229), .Y(n13339) );
  NAND2X1 U14056 ( .A(n13342), .B(n13343), .Y(n13229) );
  NAND2X1 U14057 ( .A(n13344), .B(n8799), .Y(n13343) );
  INVX1 U14058 ( .A(G21563), .Y(n8799) );
  OR2X1 U14059 ( .A(n13272), .B(G21558), .Y(n13344) );
  NAND2X1 U14060 ( .A(G21558), .B(n13272), .Y(n13342) );
  NAND2X1 U14061 ( .A(n13345), .B(n13346), .Y(n13272) );
  NAND2X1 U14062 ( .A(n13347), .B(n8800), .Y(n13346) );
  INVX1 U14063 ( .A(G21564), .Y(n8800) );
  NAND2X1 U14064 ( .A(n8893), .B(n13253), .Y(n13347) );
  OR2X1 U14065 ( .A(n8893), .B(n13253), .Y(n13345) );
  NAND2X1 U14066 ( .A(n8887), .B(n13348), .Y(n13253) );
  NAND2X1 U14067 ( .A(n13349), .B(n13267), .Y(n13348) );
  NAND2X1 U14068 ( .A(G21561), .B(n8540), .Y(n13267) );
  INVX1 U14069 ( .A(G21566), .Y(n8540) );
  NAND2X1 U14070 ( .A(G21560), .B(n8880), .Y(n13349) );
  INVX1 U14071 ( .A(G21565), .Y(n8880) );
  NAND2X1 U14072 ( .A(G21565), .B(n10945), .Y(n8887) );
  AND2X1 U14073 ( .A(n8827), .B(n13350), .Y(n13227) );
  NAND2X1 U14074 ( .A(n13223), .B(n13166), .Y(n13350) );
  INVX1 U14075 ( .A(n9631), .Y(n13166) );
  NOR2X1 U14076 ( .A(n8772), .B(n7451), .Y(n9631) );
  NOR3X1 U14077 ( .A(n7455), .B(n7451), .C(n9751), .Y(n13223) );
  INVX1 U14078 ( .A(n8762), .Y(n7455) );
  NOR2X1 U14079 ( .A(G21425), .B(G21427), .Y(n8827) );
  INVX1 U14080 ( .A(n10013), .Y(n12843) );
  NOR2X1 U14081 ( .A(n7424), .B(n8817), .Y(n10013) );
  INVX1 U14082 ( .A(n9207), .Y(n7424) );
  NOR3X1 U14083 ( .A(n8711), .B(n7444), .C(n8858), .Y(n9207) );
  NAND2X1 U14084 ( .A(n9285), .B(n7456), .Y(n8858) );
  AND2X1 U14085 ( .A(n9751), .B(n13212), .Y(n9285) );
  NOR3X1 U14086 ( .A(n12784), .B(n7442), .C(n12707), .Y(n13212) );
  INVX1 U14087 ( .A(n8782), .Y(n12784) );
  NAND4X1 U14088 ( .A(n13351), .B(n13352), .C(n13353), .D(n13354), .Y(n8782)
         );
  NOR4X1 U14089 ( .A(n13355), .B(n13356), .C(n13357), .D(n13358), .Y(n13354)
         );
  NOR2X1 U14090 ( .A(n13359), .B(n10312), .Y(n13358) );
  INVX1 U14091 ( .A(G21437), .Y(n10312) );
  NOR2X1 U14092 ( .A(n13360), .B(n10314), .Y(n13357) );
  INVX1 U14093 ( .A(G21445), .Y(n10314) );
  NOR2X1 U14094 ( .A(n13361), .B(n10316), .Y(n13356) );
  INVX1 U14095 ( .A(G21453), .Y(n10316) );
  NOR2X1 U14096 ( .A(n13362), .B(n10324), .Y(n13355) );
  INVX1 U14097 ( .A(G21469), .Y(n10324) );
  NOR4X1 U14098 ( .A(n13363), .B(n13364), .C(n13365), .D(n13366), .Y(n13353)
         );
  NOR2X1 U14099 ( .A(n13367), .B(n10326), .Y(n13366) );
  INVX1 U14100 ( .A(G21477), .Y(n10326) );
  NOR2X1 U14101 ( .A(n13368), .B(n10328), .Y(n13365) );
  INVX1 U14102 ( .A(G21485), .Y(n10328) );
  NOR2X1 U14103 ( .A(n13369), .B(n10972), .Y(n13364) );
  INVX1 U14104 ( .A(G21501), .Y(n10972) );
  NOR2X1 U14105 ( .A(n13370), .B(n10967), .Y(n13363) );
  INVX1 U14106 ( .A(G21509), .Y(n10967) );
  NOR4X1 U14107 ( .A(n13371), .B(n13372), .C(n13373), .D(n13374), .Y(n13352)
         );
  NOR2X1 U14108 ( .A(n13375), .B(n10983), .Y(n13374) );
  INVX1 U14109 ( .A(G21517), .Y(n10983) );
  NOR2X1 U14110 ( .A(n13376), .B(n10965), .Y(n13373) );
  INVX1 U14111 ( .A(G21533), .Y(n10965) );
  NOR2X1 U14112 ( .A(n13377), .B(n10964), .Y(n13372) );
  INVX1 U14113 ( .A(G21541), .Y(n10964) );
  NOR2X1 U14114 ( .A(n13378), .B(n10982), .Y(n13371) );
  INVX1 U14115 ( .A(G21549), .Y(n10982) );
  NOR4X1 U14116 ( .A(n13379), .B(n13380), .C(n13381), .D(n13382), .Y(n13351)
         );
  NOR2X1 U14117 ( .A(n13383), .B(n10310), .Y(n13382) );
  INVX1 U14118 ( .A(G21429), .Y(n10310) );
  NOR2X1 U14119 ( .A(n13384), .B(n10322), .Y(n13381) );
  INVX1 U14120 ( .A(G21461), .Y(n10322) );
  NOR2X1 U14121 ( .A(n13385), .B(n10973), .Y(n13380) );
  INVX1 U14122 ( .A(G21493), .Y(n10973) );
  NOR2X1 U14123 ( .A(n13386), .B(n10966), .Y(n13379) );
  INVX1 U14124 ( .A(G21525), .Y(n10966) );
  NAND2X1 U14125 ( .A(n12910), .B(n13026), .Y(n13021) );
  NOR2X1 U14126 ( .A(n8817), .B(n10116), .Y(n13026) );
  NOR2X1 U14127 ( .A(n8929), .B(n13387), .Y(n10116) );
  NOR2X1 U14128 ( .A(n8955), .B(G21391), .Y(n13387) );
  INVX1 U14129 ( .A(G21390), .Y(n8955) );
  NOR2X1 U14130 ( .A(n8938), .B(G21390), .Y(n8929) );
  INVX1 U14131 ( .A(G21391), .Y(n8938) );
  INVX1 U14132 ( .A(G21428), .Y(n8817) );
  AND3X1 U14133 ( .A(n9185), .B(n9751), .C(n13388), .Y(n12910) );
  NOR3X1 U14134 ( .A(n12707), .B(n7442), .C(n7439), .Y(n13388) );
  INVX1 U14135 ( .A(n7456), .Y(n7439) );
  NAND4X1 U14136 ( .A(n13389), .B(n13390), .C(n13391), .D(n13392), .Y(n7456)
         );
  NOR4X1 U14137 ( .A(n13393), .B(n13394), .C(n13395), .D(n13396), .Y(n13392)
         );
  NOR2X1 U14138 ( .A(n13359), .B(n10728), .Y(n13396) );
  INVX1 U14139 ( .A(G21442), .Y(n10728) );
  NOR2X1 U14140 ( .A(n13360), .B(n10729), .Y(n13395) );
  INVX1 U14141 ( .A(G21450), .Y(n10729) );
  NOR2X1 U14142 ( .A(n13361), .B(n10730), .Y(n13394) );
  INVX1 U14143 ( .A(G21458), .Y(n10730) );
  NOR2X1 U14144 ( .A(n13362), .B(n10736), .Y(n13393) );
  INVX1 U14145 ( .A(G21474), .Y(n10736) );
  NOR4X1 U14146 ( .A(n13397), .B(n13398), .C(n13399), .D(n13400), .Y(n13391)
         );
  NOR2X1 U14147 ( .A(n13367), .B(n10737), .Y(n13400) );
  INVX1 U14148 ( .A(G21482), .Y(n10737) );
  NOR2X1 U14149 ( .A(n13368), .B(n10738), .Y(n13399) );
  INVX1 U14150 ( .A(G21490), .Y(n10738) );
  NOR2X1 U14151 ( .A(n13369), .B(n10753), .Y(n13398) );
  INVX1 U14152 ( .A(G21506), .Y(n10753) );
  NOR2X1 U14153 ( .A(n13370), .B(n10752), .Y(n13397) );
  INVX1 U14154 ( .A(G21514), .Y(n10752) );
  NOR4X1 U14155 ( .A(n13401), .B(n13402), .C(n13403), .D(n13404), .Y(n13390)
         );
  NOR2X1 U14156 ( .A(n13375), .B(n10751), .Y(n13404) );
  INVX1 U14157 ( .A(G21522), .Y(n10751) );
  NOR2X1 U14158 ( .A(n13376), .B(n10745), .Y(n13403) );
  INVX1 U14159 ( .A(G21538), .Y(n10745) );
  NOR2X1 U14160 ( .A(n13377), .B(n10744), .Y(n13402) );
  INVX1 U14161 ( .A(G21546), .Y(n10744) );
  NOR2X1 U14162 ( .A(n13378), .B(n10743), .Y(n13401) );
  INVX1 U14163 ( .A(G21554), .Y(n10743) );
  NOR4X1 U14164 ( .A(n13405), .B(n13406), .C(n13407), .D(n13408), .Y(n13389)
         );
  NOR2X1 U14165 ( .A(n13383), .B(n10727), .Y(n13408) );
  INVX1 U14166 ( .A(G21434), .Y(n10727) );
  NOR2X1 U14167 ( .A(n13384), .B(n10735), .Y(n13407) );
  INVX1 U14168 ( .A(G21466), .Y(n10735) );
  NOR2X1 U14169 ( .A(n13385), .B(n10754), .Y(n13406) );
  INVX1 U14170 ( .A(G21498), .Y(n10754) );
  NOR2X1 U14171 ( .A(n13386), .B(n10746), .Y(n13405) );
  INVX1 U14172 ( .A(G21530), .Y(n10746) );
  INVX1 U14173 ( .A(n8772), .Y(n7442) );
  NAND4X1 U14174 ( .A(n13409), .B(n13410), .C(n13411), .D(n13412), .Y(n8772)
         );
  NOR4X1 U14175 ( .A(n13413), .B(n13414), .C(n13415), .D(n13416), .Y(n13412)
         );
  NOR2X1 U14176 ( .A(n13359), .B(n10390), .Y(n13416) );
  INVX1 U14177 ( .A(G21438), .Y(n10390) );
  NOR2X1 U14178 ( .A(n13360), .B(n10391), .Y(n13415) );
  INVX1 U14179 ( .A(G21446), .Y(n10391) );
  NOR2X1 U14180 ( .A(n13361), .B(n10392), .Y(n13414) );
  INVX1 U14181 ( .A(G21454), .Y(n10392) );
  NOR2X1 U14182 ( .A(n13362), .B(n10398), .Y(n13413) );
  INVX1 U14183 ( .A(G21470), .Y(n10398) );
  NOR4X1 U14184 ( .A(n13417), .B(n13418), .C(n13419), .D(n13420), .Y(n13411)
         );
  NOR2X1 U14185 ( .A(n13367), .B(n10399), .Y(n13420) );
  INVX1 U14186 ( .A(G21478), .Y(n10399) );
  NOR2X1 U14187 ( .A(n13368), .B(n10400), .Y(n13419) );
  INVX1 U14188 ( .A(G21486), .Y(n10400) );
  NOR2X1 U14189 ( .A(n13369), .B(n10421), .Y(n13418) );
  INVX1 U14190 ( .A(G21502), .Y(n10421) );
  NOR2X1 U14191 ( .A(n13370), .B(n10419), .Y(n13417) );
  INVX1 U14192 ( .A(G21510), .Y(n10419) );
  NOR4X1 U14193 ( .A(n13421), .B(n13422), .C(n13423), .D(n13424), .Y(n13410)
         );
  NOR2X1 U14194 ( .A(n13375), .B(n10417), .Y(n13424) );
  INVX1 U14195 ( .A(G21518), .Y(n10417) );
  NOR2X1 U14196 ( .A(n13376), .B(n10409), .Y(n13423) );
  INVX1 U14197 ( .A(G21534), .Y(n10409) );
  NOR2X1 U14198 ( .A(n13377), .B(n10407), .Y(n13422) );
  INVX1 U14199 ( .A(G21542), .Y(n10407) );
  NOR2X1 U14200 ( .A(n13378), .B(n10405), .Y(n13421) );
  INVX1 U14201 ( .A(G21550), .Y(n10405) );
  NOR4X1 U14202 ( .A(n13425), .B(n13426), .C(n13427), .D(n13428), .Y(n13409)
         );
  NOR2X1 U14203 ( .A(n13383), .B(n10389), .Y(n13428) );
  INVX1 U14204 ( .A(G21430), .Y(n10389) );
  NOR2X1 U14205 ( .A(n13384), .B(n10397), .Y(n13427) );
  INVX1 U14206 ( .A(G21462), .Y(n10397) );
  NOR2X1 U14207 ( .A(n13385), .B(n10423), .Y(n13426) );
  INVX1 U14208 ( .A(G21494), .Y(n10423) );
  NOR2X1 U14209 ( .A(n13386), .B(n10411), .Y(n13425) );
  INVX1 U14210 ( .A(G21526), .Y(n10411) );
  NAND2X1 U14211 ( .A(n7446), .B(n8762), .Y(n12707) );
  NAND4X1 U14212 ( .A(n13429), .B(n13430), .C(n13431), .D(n13432), .Y(n8762)
         );
  NOR4X1 U14213 ( .A(n13433), .B(n13434), .C(n13435), .D(n13436), .Y(n13432)
         );
  NOR2X1 U14214 ( .A(n13359), .B(n10492), .Y(n13436) );
  INVX1 U14215 ( .A(G21439), .Y(n10492) );
  NOR2X1 U14216 ( .A(n13360), .B(n10493), .Y(n13435) );
  INVX1 U14217 ( .A(G21447), .Y(n10493) );
  NOR2X1 U14218 ( .A(n13361), .B(n10494), .Y(n13434) );
  INVX1 U14219 ( .A(G21455), .Y(n10494) );
  NOR2X1 U14220 ( .A(n13362), .B(n10500), .Y(n13433) );
  INVX1 U14221 ( .A(G21471), .Y(n10500) );
  NOR4X1 U14222 ( .A(n13437), .B(n13438), .C(n13439), .D(n13440), .Y(n13431)
         );
  NOR2X1 U14223 ( .A(n13367), .B(n10501), .Y(n13440) );
  INVX1 U14224 ( .A(G21479), .Y(n10501) );
  NOR2X1 U14225 ( .A(n13368), .B(n10502), .Y(n13439) );
  INVX1 U14226 ( .A(G21487), .Y(n10502) );
  NOR2X1 U14227 ( .A(n13369), .B(n11105), .Y(n13438) );
  INVX1 U14228 ( .A(G21503), .Y(n11105) );
  NOR2X1 U14229 ( .A(n13370), .B(n11100), .Y(n13437) );
  INVX1 U14230 ( .A(G21511), .Y(n11100) );
  NOR4X1 U14231 ( .A(n13441), .B(n13442), .C(n13443), .D(n13444), .Y(n13430)
         );
  NOR2X1 U14232 ( .A(n13375), .B(n11116), .Y(n13444) );
  INVX1 U14233 ( .A(G21519), .Y(n11116) );
  NOR2X1 U14234 ( .A(n13376), .B(n11098), .Y(n13443) );
  INVX1 U14235 ( .A(G21535), .Y(n11098) );
  NOR2X1 U14236 ( .A(n13377), .B(n11097), .Y(n13442) );
  INVX1 U14237 ( .A(G21543), .Y(n11097) );
  NOR2X1 U14238 ( .A(n13378), .B(n11115), .Y(n13441) );
  INVX1 U14239 ( .A(G21551), .Y(n11115) );
  NOR4X1 U14240 ( .A(n13445), .B(n13446), .C(n13447), .D(n13448), .Y(n13429)
         );
  NOR2X1 U14241 ( .A(n13383), .B(n10491), .Y(n13448) );
  INVX1 U14242 ( .A(G21431), .Y(n10491) );
  NOR2X1 U14243 ( .A(n13384), .B(n10499), .Y(n13447) );
  INVX1 U14244 ( .A(G21463), .Y(n10499) );
  NOR2X1 U14245 ( .A(n13385), .B(n11106), .Y(n13446) );
  INVX1 U14246 ( .A(G21495), .Y(n11106) );
  NOR2X1 U14247 ( .A(n13386), .B(n11099), .Y(n13445) );
  INVX1 U14248 ( .A(G21527), .Y(n11099) );
  INVX1 U14249 ( .A(n7458), .Y(n7446) );
  NAND4X1 U14250 ( .A(n13449), .B(n13450), .C(n13451), .D(n13452), .Y(n7458)
         );
  NOR4X1 U14251 ( .A(n13453), .B(n13454), .C(n13455), .D(n13456), .Y(n13452)
         );
  NOR2X1 U14252 ( .A(n13359), .B(n10557), .Y(n13456) );
  INVX1 U14253 ( .A(G21440), .Y(n10557) );
  NOR2X1 U14254 ( .A(n13360), .B(n10558), .Y(n13455) );
  INVX1 U14255 ( .A(G21448), .Y(n10558) );
  NOR2X1 U14256 ( .A(n13361), .B(n10559), .Y(n13454) );
  INVX1 U14257 ( .A(G21456), .Y(n10559) );
  NOR2X1 U14258 ( .A(n13362), .B(n10565), .Y(n13453) );
  INVX1 U14259 ( .A(G21472), .Y(n10565) );
  NOR4X1 U14260 ( .A(n13457), .B(n13458), .C(n13459), .D(n13460), .Y(n13451)
         );
  NOR2X1 U14261 ( .A(n13367), .B(n10566), .Y(n13460) );
  INVX1 U14262 ( .A(G21480), .Y(n10566) );
  NOR2X1 U14263 ( .A(n13368), .B(n10567), .Y(n13459) );
  INVX1 U14264 ( .A(G21488), .Y(n10567) );
  NOR2X1 U14265 ( .A(n13369), .B(n10582), .Y(n13458) );
  INVX1 U14266 ( .A(G21504), .Y(n10582) );
  NOR2X1 U14267 ( .A(n13370), .B(n10581), .Y(n13457) );
  INVX1 U14268 ( .A(G21512), .Y(n10581) );
  NOR4X1 U14269 ( .A(n13461), .B(n13462), .C(n13463), .D(n13464), .Y(n13450)
         );
  NOR2X1 U14270 ( .A(n13375), .B(n10580), .Y(n13464) );
  INVX1 U14271 ( .A(G21520), .Y(n10580) );
  NOR2X1 U14272 ( .A(n13376), .B(n10574), .Y(n13463) );
  INVX1 U14273 ( .A(G21536), .Y(n10574) );
  NOR2X1 U14274 ( .A(n13377), .B(n10573), .Y(n13462) );
  INVX1 U14275 ( .A(G21544), .Y(n10573) );
  NOR2X1 U14276 ( .A(n13378), .B(n10572), .Y(n13461) );
  INVX1 U14277 ( .A(G21552), .Y(n10572) );
  NOR4X1 U14278 ( .A(n13465), .B(n13466), .C(n13467), .D(n13468), .Y(n13449)
         );
  NOR2X1 U14279 ( .A(n13383), .B(n10556), .Y(n13468) );
  INVX1 U14280 ( .A(G21432), .Y(n10556) );
  NOR2X1 U14281 ( .A(n13384), .B(n10564), .Y(n13467) );
  INVX1 U14282 ( .A(G21464), .Y(n10564) );
  NOR2X1 U14283 ( .A(n13385), .B(n10583), .Y(n13466) );
  INVX1 U14284 ( .A(G21496), .Y(n10583) );
  NOR2X1 U14285 ( .A(n13386), .B(n10575), .Y(n13465) );
  INVX1 U14286 ( .A(G21528), .Y(n10575) );
  INVX1 U14287 ( .A(n8743), .Y(n9751) );
  NAND4X1 U14288 ( .A(n13469), .B(n13470), .C(n13471), .D(n13472), .Y(n8743)
         );
  NOR4X1 U14289 ( .A(n13473), .B(n13474), .C(n13475), .D(n13476), .Y(n13472)
         );
  NOR2X1 U14290 ( .A(n13359), .B(n10639), .Y(n13476) );
  INVX1 U14291 ( .A(G21441), .Y(n10639) );
  NOR2X1 U14292 ( .A(n13360), .B(n10640), .Y(n13475) );
  INVX1 U14293 ( .A(G21449), .Y(n10640) );
  NOR2X1 U14294 ( .A(n13361), .B(n10641), .Y(n13474) );
  INVX1 U14295 ( .A(G21457), .Y(n10641) );
  NOR2X1 U14296 ( .A(n13362), .B(n10647), .Y(n13473) );
  INVX1 U14297 ( .A(G21473), .Y(n10647) );
  NOR4X1 U14298 ( .A(n13477), .B(n13478), .C(n13479), .D(n13480), .Y(n13471)
         );
  NOR2X1 U14299 ( .A(n13367), .B(n10648), .Y(n13480) );
  INVX1 U14300 ( .A(G21481), .Y(n10648) );
  NOR2X1 U14301 ( .A(n13368), .B(n10649), .Y(n13479) );
  INVX1 U14302 ( .A(G21489), .Y(n10649) );
  NOR2X1 U14303 ( .A(n13369), .B(n10664), .Y(n13478) );
  INVX1 U14304 ( .A(G21505), .Y(n10664) );
  NOR2X1 U14305 ( .A(n13370), .B(n10663), .Y(n13477) );
  INVX1 U14306 ( .A(G21513), .Y(n10663) );
  NOR4X1 U14307 ( .A(n13481), .B(n13482), .C(n13483), .D(n13484), .Y(n13470)
         );
  NOR2X1 U14308 ( .A(n13375), .B(n10662), .Y(n13484) );
  INVX1 U14309 ( .A(G21521), .Y(n10662) );
  NOR2X1 U14310 ( .A(n13376), .B(n10656), .Y(n13483) );
  INVX1 U14311 ( .A(G21537), .Y(n10656) );
  NOR2X1 U14312 ( .A(n13377), .B(n10655), .Y(n13482) );
  INVX1 U14313 ( .A(G21545), .Y(n10655) );
  NOR2X1 U14314 ( .A(n13378), .B(n10654), .Y(n13481) );
  INVX1 U14315 ( .A(G21553), .Y(n10654) );
  NOR4X1 U14316 ( .A(n13485), .B(n13486), .C(n13487), .D(n13488), .Y(n13469)
         );
  NOR2X1 U14317 ( .A(n13383), .B(n10638), .Y(n13488) );
  INVX1 U14318 ( .A(G21433), .Y(n10638) );
  NOR2X1 U14319 ( .A(n13384), .B(n10646), .Y(n13487) );
  INVX1 U14320 ( .A(G21465), .Y(n10646) );
  NOR2X1 U14321 ( .A(n13385), .B(n10665), .Y(n13486) );
  INVX1 U14322 ( .A(G21497), .Y(n10665) );
  NOR2X1 U14323 ( .A(n13386), .B(n10657), .Y(n13485) );
  INVX1 U14324 ( .A(G21529), .Y(n10657) );
  NOR2X1 U14325 ( .A(n8711), .B(n7451), .Y(n9185) );
  INVX1 U14326 ( .A(n7444), .Y(n7451) );
  NAND4X1 U14327 ( .A(n13489), .B(n13490), .C(n13491), .D(n13492), .Y(n7444)
         );
  NOR4X1 U14328 ( .A(n13493), .B(n13494), .C(n13495), .D(n13496), .Y(n13492)
         );
  NOR2X1 U14329 ( .A(n13359), .B(n10818), .Y(n13496) );
  INVX1 U14330 ( .A(G21443), .Y(n10818) );
  NOR2X1 U14331 ( .A(n13360), .B(n10819), .Y(n13495) );
  INVX1 U14332 ( .A(G21451), .Y(n10819) );
  NOR2X1 U14333 ( .A(n13361), .B(n10820), .Y(n13494) );
  INVX1 U14334 ( .A(G21459), .Y(n10820) );
  NOR2X1 U14335 ( .A(n13362), .B(n10826), .Y(n13493) );
  INVX1 U14336 ( .A(G21475), .Y(n10826) );
  NOR4X1 U14337 ( .A(n13497), .B(n13498), .C(n13499), .D(n13500), .Y(n13491)
         );
  NOR2X1 U14338 ( .A(n13367), .B(n10827), .Y(n13500) );
  INVX1 U14339 ( .A(G21483), .Y(n10827) );
  NOR2X1 U14340 ( .A(n13368), .B(n10828), .Y(n13499) );
  INVX1 U14341 ( .A(G21491), .Y(n10828) );
  NOR2X1 U14342 ( .A(n13369), .B(n10843), .Y(n13498) );
  INVX1 U14343 ( .A(G21507), .Y(n10843) );
  NOR2X1 U14344 ( .A(n13370), .B(n10842), .Y(n13497) );
  INVX1 U14345 ( .A(G21515), .Y(n10842) );
  NOR4X1 U14346 ( .A(n13501), .B(n13502), .C(n13503), .D(n13504), .Y(n13490)
         );
  NOR2X1 U14347 ( .A(n13375), .B(n10841), .Y(n13504) );
  INVX1 U14348 ( .A(G21523), .Y(n10841) );
  NOR2X1 U14349 ( .A(n13376), .B(n10835), .Y(n13503) );
  INVX1 U14350 ( .A(G21539), .Y(n10835) );
  NOR2X1 U14351 ( .A(n13377), .B(n10834), .Y(n13502) );
  INVX1 U14352 ( .A(G21547), .Y(n10834) );
  NOR2X1 U14353 ( .A(n13378), .B(n10833), .Y(n13501) );
  INVX1 U14354 ( .A(G21555), .Y(n10833) );
  NOR4X1 U14355 ( .A(n13505), .B(n13506), .C(n13507), .D(n13508), .Y(n13489)
         );
  NOR2X1 U14356 ( .A(n13383), .B(n10817), .Y(n13508) );
  INVX1 U14357 ( .A(G21435), .Y(n10817) );
  NOR2X1 U14358 ( .A(n13384), .B(n10825), .Y(n13507) );
  INVX1 U14359 ( .A(G21467), .Y(n10825) );
  NOR2X1 U14360 ( .A(n13385), .B(n10844), .Y(n13506) );
  INVX1 U14361 ( .A(G21499), .Y(n10844) );
  NOR2X1 U14362 ( .A(n13386), .B(n10836), .Y(n13505) );
  INVX1 U14363 ( .A(G21531), .Y(n10836) );
  NOR4X1 U14364 ( .A(n13513), .B(n13514), .C(n13515), .D(n13516), .Y(n13512)
         );
  NOR2X1 U14365 ( .A(n13359), .B(n10907), .Y(n13516) );
  INVX1 U14366 ( .A(G21444), .Y(n10907) );
  NAND2X1 U14367 ( .A(n13517), .B(n10944), .Y(n13359) );
  NOR2X1 U14368 ( .A(n13360), .B(n10909), .Y(n13515) );
  INVX1 U14369 ( .A(G21452), .Y(n10909) );
  NAND2X1 U14370 ( .A(n9135), .B(n13517), .Y(n13360) );
  NOR2X1 U14371 ( .A(n13361), .B(n10911), .Y(n13514) );
  INVX1 U14372 ( .A(G21460), .Y(n10911) );
  NAND2X1 U14373 ( .A(n8889), .B(n13517), .Y(n13361) );
  NOR2X1 U14374 ( .A(n13362), .B(n10918), .Y(n13513) );
  INVX1 U14375 ( .A(G21476), .Y(n10918) );
  NAND2X1 U14376 ( .A(n13197), .B(n10944), .Y(n13362) );
  NOR4X1 U14377 ( .A(n13518), .B(n13519), .C(n13520), .D(n13521), .Y(n13511)
         );
  NOR2X1 U14378 ( .A(n13367), .B(n10919), .Y(n13521) );
  INVX1 U14379 ( .A(G21484), .Y(n10919) );
  NAND2X1 U14380 ( .A(n9135), .B(n13197), .Y(n13367) );
  NOR2X1 U14381 ( .A(n13368), .B(n10922), .Y(n13520) );
  INVX1 U14382 ( .A(G21492), .Y(n10922) );
  NAND2X1 U14383 ( .A(n8889), .B(n13197), .Y(n13368) );
  NOR2X1 U14384 ( .A(n13369), .B(n10941), .Y(n13519) );
  INVX1 U14385 ( .A(G21508), .Y(n10941) );
  NAND2X1 U14386 ( .A(n13198), .B(n10944), .Y(n13369) );
  NOR2X1 U14387 ( .A(n13370), .B(n10940), .Y(n13518) );
  INVX1 U14388 ( .A(G21516), .Y(n10940) );
  NAND2X1 U14389 ( .A(n13198), .B(n9135), .Y(n13370) );
  NOR4X1 U14390 ( .A(n13522), .B(n13523), .C(n13524), .D(n13525), .Y(n13510)
         );
  NOR2X1 U14391 ( .A(n13375), .B(n10939), .Y(n13525) );
  INVX1 U14392 ( .A(G21524), .Y(n10939) );
  NAND2X1 U14393 ( .A(n13198), .B(n8889), .Y(n13375) );
  NOR2X1 U14394 ( .A(n13376), .B(n10931), .Y(n13524) );
  INVX1 U14395 ( .A(G21540), .Y(n10931) );
  NAND2X1 U14396 ( .A(n10949), .B(n10944), .Y(n13376) );
  NOR2X1 U14397 ( .A(n10945), .B(G21561), .Y(n10944) );
  NOR2X1 U14398 ( .A(n13377), .B(n10929), .Y(n13523) );
  INVX1 U14399 ( .A(G21548), .Y(n10929) );
  NAND2X1 U14400 ( .A(n10949), .B(n9135), .Y(n13377) );
  NOR2X1 U14401 ( .A(n8890), .B(G21560), .Y(n9135) );
  NOR2X1 U14402 ( .A(n13378), .B(n10927), .Y(n13522) );
  INVX1 U14403 ( .A(G21556), .Y(n10927) );
  NAND2X1 U14404 ( .A(n10949), .B(n8889), .Y(n13378) );
  NOR2X1 U14405 ( .A(G21560), .B(G21561), .Y(n8889) );
  NOR4X1 U14406 ( .A(n13526), .B(n13527), .C(n13528), .D(n13529), .Y(n13509)
         );
  NOR2X1 U14407 ( .A(n13383), .B(n10904), .Y(n13529) );
  INVX1 U14408 ( .A(G21436), .Y(n10904) );
  NAND2X1 U14409 ( .A(n10952), .B(n13517), .Y(n13383) );
  NOR2X1 U14410 ( .A(n8870), .B(n8893), .Y(n13517) );
  NOR2X1 U14411 ( .A(n13384), .B(n10916), .Y(n13528) );
  INVX1 U14412 ( .A(G21468), .Y(n10916) );
  NAND2X1 U14413 ( .A(n10952), .B(n13197), .Y(n13384) );
  NOR2X1 U14414 ( .A(n8870), .B(G21559), .Y(n13197) );
  INVX1 U14415 ( .A(G21558), .Y(n8870) );
  NOR2X1 U14416 ( .A(n13385), .B(n10942), .Y(n13527) );
  INVX1 U14417 ( .A(G21500), .Y(n10942) );
  NAND2X1 U14418 ( .A(n10952), .B(n13198), .Y(n13385) );
  NOR2X1 U14419 ( .A(n8893), .B(G21558), .Y(n13198) );
  INVX1 U14420 ( .A(G21559), .Y(n8893) );
  NOR2X1 U14421 ( .A(n13386), .B(n10932), .Y(n13526) );
  INVX1 U14422 ( .A(G21532), .Y(n10932) );
  NAND2X1 U14423 ( .A(n10952), .B(n10949), .Y(n13386) );
  NOR2X1 U14424 ( .A(G21558), .B(G21559), .Y(n10949) );
  NOR2X1 U14425 ( .A(n10945), .B(n8890), .Y(n10952) );
  INVX1 U14426 ( .A(G21561), .Y(n8890) );
  INVX1 U14427 ( .A(G21560), .Y(n10945) );
endmodule

